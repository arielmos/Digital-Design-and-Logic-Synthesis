
module Block_To_Pixel ( clk, rst, M2, block_in, block_done, Pixel_Data, Ready, 
        new_pixel, last_Block, Image_Done );
  input [19:0] M2;
  input [31:0] block_in;
  output [7:0] Pixel_Data;
  input clk, rst, block_done, last_Block;
  output Ready, new_pixel, Image_Done;
  wire   block_done_down, Image_DoneHelp, N36, n5, n15, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n51,
         n52, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n1,
         n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17, n18,
         n48, n53, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92;
  wire   [1:0] state;
  wire   [3:0] i;

  NOR3X4 U36 ( .A(i[0]), .B(i[2]), .C(n88), .Y(n24) );
  NOR3X4 U37 ( .A(i[1]), .B(i[2]), .C(n87), .Y(n23) );
  NOR3X4 U39 ( .A(i[0]), .B(i[1]), .C(n89), .Y(n26) );
  DFFHQX1 \Pixel_Data_reg[7]  ( .D(n73), .CK(clk), .Q(Pixel_Data[7]) );
  DFFHQX1 \Pixel_Data_reg[6]  ( .D(n72), .CK(clk), .Q(Pixel_Data[6]) );
  DFFHQX1 \Pixel_Data_reg[5]  ( .D(n71), .CK(clk), .Q(Pixel_Data[5]) );
  DFFHQX1 \Pixel_Data_reg[4]  ( .D(n70), .CK(clk), .Q(Pixel_Data[4]) );
  DFFHQX1 \Pixel_Data_reg[3]  ( .D(n69), .CK(clk), .Q(Pixel_Data[3]) );
  DFFHQX1 \Pixel_Data_reg[2]  ( .D(n68), .CK(clk), .Q(Pixel_Data[2]) );
  DFFHQX1 \Pixel_Data_reg[1]  ( .D(n67), .CK(clk), .Q(Pixel_Data[1]) );
  DFFHQX1 \Pixel_Data_reg[0]  ( .D(n66), .CK(clk), .Q(Pixel_Data[0]) );
  DFFHQX1 Image_DoneHelp_reg ( .D(n74), .CK(clk), .Q(Image_DoneHelp) );
  DFFHQX1 block_done_down_reg ( .D(n78), .CK(clk), .Q(block_done_down) );
  DFFTRX1 \state_reg[1]  ( .D(n92), .RN(n82), .CK(clk), .Q(state[1]), .QN(n15)
         );
  DFFHQX1 Ready_reg ( .D(n85), .CK(clk), .Q(Ready) );
  DFFHQX1 \state_reg[0]  ( .D(n79), .CK(clk), .Q(state[0]) );
  DFFX1 \i_reg[3]  ( .D(n77), .CK(clk), .Q(i[3]), .QN(n5) );
  EDFFTRX1 new_pixel_reg ( .RN(n92), .D(n63), .E(n82), .CK(clk), .Q(new_pixel)
         );
  DFFTRX1 Image_Done_reg ( .D(n92), .RN(n2), .CK(clk), .Q(Image_Done) );
  DFFHQX2 \i_reg[2]  ( .D(n83), .CK(clk), .Q(i[2]) );
  DFFHQX2 \i_reg[0]  ( .D(n76), .CK(clk), .Q(i[0]) );
  DFFHQX2 \i_reg[1]  ( .D(n75), .CK(clk), .Q(i[1]) );
  AOI22XL U3 ( .A0(i[1]), .A1(n53), .B0(n6), .B1(i[0]), .Y(n10) );
  NAND4XL U4 ( .A(i[0]), .B(n1), .C(n84), .D(n88), .Y(n58) );
  CLKINVX3 U5 ( .A(n59), .Y(n84) );
  CLKINVX3 U6 ( .A(n3), .Y(n81) );
  AOI21X1 U7 ( .A0(n63), .A1(N36), .B0(n86), .Y(n59) );
  OAI2BB1X1 U8 ( .A0N(n56), .A1N(n1), .B0(n84), .Y(n55) );
  BUFX3 U9 ( .A(n19), .Y(n3) );
  NAND2X1 U10 ( .A(N36), .B(n1), .Y(n19) );
  OAI21XL U11 ( .A0(n87), .A1(n84), .B0(n60), .Y(n76) );
  OAI21XL U12 ( .A0(n87), .A1(n86), .B0(n84), .Y(n60) );
  AND2X2 U13 ( .A(n63), .B(n92), .Y(n1) );
  INVX1 U14 ( .A(n50), .Y(n86) );
  INVX1 U15 ( .A(rst), .Y(n92) );
  OAI32X1 U16 ( .A0(n61), .A1(n56), .A2(n89), .B0(n62), .B1(n5), .Y(n77) );
  NAND3X1 U17 ( .A(n84), .B(n5), .C(n1), .Y(n61) );
  AOI21X1 U18 ( .A0(n1), .A1(n89), .B0(n55), .Y(n62) );
  INVX1 U19 ( .A(n54), .Y(n83) );
  AOI32X1 U20 ( .A0(n4), .A1(n84), .A2(n1), .B0(n55), .B1(i[2]), .Y(n54) );
  OAI21XL U21 ( .A0(n57), .A1(n88), .B0(n58), .Y(n75) );
  AOI21X1 U22 ( .A0(n1), .A1(n87), .B0(n59), .Y(n57) );
  AOI21X1 U23 ( .A0(n3), .A1(n64), .B0(n65), .Y(n79) );
  NAND2X1 U24 ( .A(n51), .B(n92), .Y(n64) );
  AOI21X1 U25 ( .A0(block_done), .A1(block_done_down), .B0(n63), .Y(n65) );
  OAI2BB1X1 U26 ( .A0N(Pixel_Data[0]), .A1N(n3), .B0(n20), .Y(n66) );
  OAI2BB1X1 U27 ( .A0N(n21), .A1N(n22), .B0(n81), .Y(n20) );
  AOI22X1 U28 ( .A0(block_in[0]), .A1(n23), .B0(block_in[8]), .B1(n24), .Y(n22) );
  AOI22X1 U29 ( .A0(block_in[16]), .A1(n4), .B0(block_in[24]), .B1(n26), .Y(
        n21) );
  OAI2BB1X1 U30 ( .A0N(Pixel_Data[1]), .A1N(n3), .B0(n27), .Y(n67) );
  OAI2BB1X1 U31 ( .A0N(n28), .A1N(n29), .B0(n81), .Y(n27) );
  AOI22X1 U32 ( .A0(block_in[1]), .A1(n23), .B0(block_in[9]), .B1(n24), .Y(n29) );
  AOI22X1 U33 ( .A0(block_in[17]), .A1(n4), .B0(block_in[25]), .B1(n26), .Y(
        n28) );
  OAI2BB1X1 U34 ( .A0N(Pixel_Data[2]), .A1N(n3), .B0(n30), .Y(n68) );
  OAI2BB1X1 U35 ( .A0N(n31), .A1N(n32), .B0(n81), .Y(n30) );
  AOI22X1 U38 ( .A0(block_in[2]), .A1(n23), .B0(block_in[10]), .B1(n24), .Y(
        n32) );
  AOI22X1 U40 ( .A0(block_in[18]), .A1(n4), .B0(block_in[26]), .B1(n26), .Y(
        n31) );
  OAI2BB1X1 U41 ( .A0N(Pixel_Data[3]), .A1N(n3), .B0(n33), .Y(n69) );
  OAI2BB1X1 U42 ( .A0N(n34), .A1N(n35), .B0(n81), .Y(n33) );
  AOI22X1 U43 ( .A0(block_in[3]), .A1(n23), .B0(block_in[11]), .B1(n24), .Y(
        n35) );
  AOI22X1 U44 ( .A0(block_in[19]), .A1(n4), .B0(block_in[27]), .B1(n26), .Y(
        n34) );
  OAI2BB1X1 U45 ( .A0N(Pixel_Data[4]), .A1N(n3), .B0(n36), .Y(n70) );
  OAI2BB1X1 U46 ( .A0N(n37), .A1N(n38), .B0(n81), .Y(n36) );
  AOI22X1 U47 ( .A0(block_in[4]), .A1(n23), .B0(block_in[12]), .B1(n24), .Y(
        n38) );
  AOI22X1 U48 ( .A0(block_in[20]), .A1(n4), .B0(block_in[28]), .B1(n26), .Y(
        n37) );
  OAI2BB1X1 U49 ( .A0N(Pixel_Data[5]), .A1N(n3), .B0(n39), .Y(n71) );
  OAI2BB1X1 U50 ( .A0N(n40), .A1N(n41), .B0(n81), .Y(n39) );
  AOI22X1 U51 ( .A0(block_in[5]), .A1(n23), .B0(block_in[13]), .B1(n24), .Y(
        n41) );
  AOI22X1 U52 ( .A0(block_in[21]), .A1(n4), .B0(block_in[29]), .B1(n26), .Y(
        n40) );
  OAI2BB1X1 U53 ( .A0N(Pixel_Data[6]), .A1N(n3), .B0(n42), .Y(n72) );
  OAI2BB1X1 U54 ( .A0N(n43), .A1N(n44), .B0(n81), .Y(n42) );
  AOI22X1 U55 ( .A0(block_in[6]), .A1(n23), .B0(block_in[14]), .B1(n24), .Y(
        n44) );
  AOI22X1 U56 ( .A0(block_in[22]), .A1(n4), .B0(block_in[30]), .B1(n26), .Y(
        n43) );
  OAI2BB1X1 U57 ( .A0N(Pixel_Data[7]), .A1N(n3), .B0(n45), .Y(n73) );
  OAI2BB1X1 U58 ( .A0N(n46), .A1N(n47), .B0(n81), .Y(n45) );
  AOI22X1 U59 ( .A0(block_in[7]), .A1(n23), .B0(block_in[15]), .B1(n24), .Y(
        n47) );
  AOI22X1 U60 ( .A0(block_in[23]), .A1(n4), .B0(block_in[31]), .B1(n26), .Y(
        n46) );
  INVX1 U61 ( .A(M2[2]), .Y(n80) );
  INVX1 U62 ( .A(M2[1]), .Y(n53) );
  INVX1 U63 ( .A(n52), .Y(n82) );
  AOI21X1 U64 ( .A0(n63), .A1(N36), .B0(state[0]), .Y(n52) );
  NOR2X2 U65 ( .A(n15), .B(state[0]), .Y(n63) );
  INVX1 U66 ( .A(i[0]), .Y(n87) );
  INVX1 U67 ( .A(i[2]), .Y(n89) );
  INVX1 U68 ( .A(i[1]), .Y(n88) );
  AOI21X1 U69 ( .A0(n15), .A1(state[0]), .B0(rst), .Y(n50) );
  NOR2X1 U70 ( .A(state[0]), .B(state[1]), .Y(n51) );
  NAND2X1 U71 ( .A(i[1]), .B(i[0]), .Y(n56) );
  BUFX3 U72 ( .A(n25), .Y(n4) );
  NOR2X1 U73 ( .A(n56), .B(i[2]), .Y(n25) );
  INVX1 U74 ( .A(n49), .Y(n85) );
  AOI211X1 U75 ( .A0(Ready), .A1(n50), .B0(n51), .C0(rst), .Y(n49) );
  AND3X2 U76 ( .A(Ready), .B(Image_DoneHelp), .C(last_Block), .Y(n2) );
  OAI32X1 U77 ( .A0(n90), .A1(rst), .A2(n51), .B0(rst), .B1(block_done), .Y(
        n78) );
  INVX1 U78 ( .A(block_done_down), .Y(n90) );
  AOI211X1 U79 ( .A0(Ready), .A1(n91), .B0(rst), .C0(n2), .Y(n74) );
  INVX1 U80 ( .A(Image_DoneHelp), .Y(n91) );
  INVX1 U81 ( .A(M2[3]), .Y(n48) );
  AOI2BB1X1 U82 ( .A0N(n53), .A1N(i[1]), .B0(M2[0]), .Y(n6) );
  NAND2BX1 U83 ( .AN(i[3]), .B(M2[3]), .Y(n7) );
  AOI32X1 U84 ( .A0(i[2]), .A1(n80), .A2(n7), .B0(n48), .B1(i[3]), .Y(n9) );
  OAI21XL U85 ( .A0(i[2]), .A1(n80), .B0(n7), .Y(n8) );
  AOI22X1 U86 ( .A0(n10), .A1(n9), .B0(n9), .B1(n8), .Y(n18) );
  NOR2X1 U87 ( .A(M2[11]), .B(M2[10]), .Y(n17) );
  NOR2X1 U88 ( .A(M2[16]), .B(M2[15]), .Y(n11) );
  NOR4BX1 U89 ( .AN(n11), .B(M2[13]), .C(M2[12]), .D(M2[14]), .Y(n16) );
  NOR3X1 U90 ( .A(M2[7]), .B(M2[9]), .C(M2[8]), .Y(n13) );
  OR4X1 U91 ( .A(M2[18]), .B(M2[17]), .C(M2[4]), .D(M2[19]), .Y(n12) );
  NOR4BX1 U92 ( .AN(n13), .B(n12), .C(M2[6]), .D(M2[5]), .Y(n14) );
  NAND4X1 U93 ( .A(n18), .B(n17), .C(n16), .D(n14), .Y(N36) );
endmodule


module Power2 ( Mu, pow );
  input [9:0] Mu;
  output [9:0] pow;
  wire   pow_7, pow_6, pow_5, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33;
  assign pow[8] = 1'b1;
  assign pow[9] = 1'b1;
  assign pow[4] = 1'b0;
  assign pow[2] = pow_7;
  assign pow[7] = pow_7;
  assign pow[0] = pow_6;
  assign pow[6] = pow_6;
  assign pow[5] = pow_5;

  NAND2X2 U3 ( .A(n6), .B(n7), .Y(pow_5) );
  OAI31X4 U4 ( .A0(n19), .A1(Mu[8]), .A2(Mu[7]), .B0(Mu[9]), .Y(n3) );
  AOI21XL U5 ( .A0(n2), .A1(n8), .B0(n3), .Y(n10) );
  AND2X2 U6 ( .A(n1), .B(n2), .Y(pow_7) );
  OAI2BB1X1 U7 ( .A0N(n3), .A1N(n4), .B0(n5), .Y(pow_6) );
  OAI21XL U8 ( .A0(n3), .A1(n8), .B0(n4), .Y(n6) );
  NAND3X1 U9 ( .A(n7), .B(n5), .C(n3), .Y(pow[1]) );
  INVX1 U10 ( .A(pow[3]), .Y(n5) );
  NAND2X1 U11 ( .A(n1), .B(n9), .Y(pow[3]) );
  OAI21XL U12 ( .A0(n10), .A1(n11), .B0(n7), .Y(n9) );
  INVX1 U13 ( .A(n4), .Y(n11) );
  NOR2BX1 U14 ( .AN(n12), .B(n13), .Y(n4) );
  OAI211X1 U15 ( .A0(n14), .A1(n15), .B0(n16), .C0(n17), .Y(n12) );
  AOI21X1 U16 ( .A0(n18), .A1(Mu[2]), .B0(Mu[3]), .Y(n14) );
  AOI31X1 U17 ( .A0(n20), .A1(n21), .A2(n22), .B0(n15), .Y(n19) );
  NOR2X1 U18 ( .A(Mu[3]), .B(Mu[2]), .Y(n22) );
  OAI31X1 U19 ( .A0(n16), .A1(n23), .A2(n24), .B0(n25), .Y(n8) );
  AOI21X1 U20 ( .A0(Mu[1]), .A1(Mu[2]), .B0(Mu[4]), .Y(n23) );
  INVX1 U21 ( .A(n26), .Y(n2) );
  AOI211X1 U22 ( .A0(n16), .A1(n27), .B0(n25), .C0(n17), .Y(n26) );
  INVX1 U23 ( .A(Mu[9]), .Y(n17) );
  INVX1 U24 ( .A(Mu[8]), .Y(n25) );
  OAI31X1 U25 ( .A0(Mu[2]), .A1(Mu[4]), .A2(n18), .B0(n28), .Y(n27) );
  INVX1 U26 ( .A(n24), .Y(n28) );
  OAI211X1 U27 ( .A0(Mu[4]), .A1(Mu[3]), .B0(Mu[5]), .C0(Mu[6]), .Y(n24) );
  NOR2X1 U28 ( .A(n21), .B(n20), .Y(n18) );
  INVX1 U29 ( .A(Mu[0]), .Y(n20) );
  INVX1 U30 ( .A(Mu[1]), .Y(n21) );
  OAI211X1 U31 ( .A0(n29), .A1(n30), .B0(n16), .C0(n13), .Y(n1) );
  NAND2X1 U32 ( .A(Mu[3]), .B(Mu[2]), .Y(n30) );
  OAI21XL U33 ( .A0(Mu[1]), .A1(Mu[0]), .B0(n31), .Y(n29) );
  OAI31X1 U34 ( .A0(n32), .A1(n33), .A2(n16), .B0(n13), .Y(n7) );
  NOR2X1 U35 ( .A(Mu[8]), .B(Mu[9]), .Y(n13) );
  INVX1 U36 ( .A(Mu[7]), .Y(n16) );
  INVX1 U37 ( .A(Mu[3]), .Y(n33) );
  OAI21XL U38 ( .A0(Mu[2]), .A1(Mu[1]), .B0(n31), .Y(n32) );
  INVX1 U39 ( .A(n15), .Y(n31) );
  NAND3X1 U40 ( .A(Mu[5]), .B(Mu[4]), .C(Mu[6]), .Y(n15) );
endmodule


module Equation_Implementation_DW_div_uns_5 ( a, b, quotient, remainder, 
        divide_by_0 );
  input [11:0] a;
  input [2:0] b;
  output [11:0] quotient;
  output [2:0] remainder;
  output divide_by_0;
  wire   n79, n80, \u_div/SumTmp[1][0] , \u_div/SumTmp[1][1] ,
         \u_div/SumTmp[1][2] , \u_div/SumTmp[2][0] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[3][0] , \u_div/SumTmp[3][1] ,
         \u_div/SumTmp[3][2] , \u_div/SumTmp[4][0] , \u_div/SumTmp[4][1] ,
         \u_div/SumTmp[4][2] , \u_div/SumTmp[5][0] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[6][0] , \u_div/SumTmp[6][1] ,
         \u_div/SumTmp[6][2] , \u_div/SumTmp[7][0] , \u_div/SumTmp[7][1] ,
         \u_div/SumTmp[7][2] , \u_div/SumTmp[8][0] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[9][0] , \u_div/SumTmp[9][1] ,
         \u_div/SumTmp[9][2] , \u_div/SumTmp[10][0] , \u_div/SumTmp[10][1] ,
         \u_div/SumTmp[11][0] , \u_div/CryTmp[0][1] , \u_div/CryTmp[1][1] ,
         \u_div/CryTmp[2][1] , \u_div/CryTmp[3][1] , \u_div/CryTmp[4][1] ,
         \u_div/CryTmp[5][1] , \u_div/CryTmp[6][1] , \u_div/CryTmp[7][1] ,
         \u_div/CryTmp[8][1] , \u_div/CryTmp[9][1] , \u_div/CryTmp[10][1] ,
         \u_div/PartRem[1][1] , \u_div/PartRem[1][3] , \u_div/PartRem[2][1] ,
         \u_div/PartRem[2][2] , \u_div/PartRem[2][3] , \u_div/PartRem[3][1] ,
         \u_div/PartRem[3][2] , \u_div/PartRem[3][3] , \u_div/PartRem[4][1] ,
         \u_div/PartRem[4][2] , \u_div/PartRem[4][3] , \u_div/PartRem[5][1] ,
         \u_div/PartRem[5][2] , \u_div/PartRem[5][3] , \u_div/PartRem[6][1] ,
         \u_div/PartRem[6][2] , \u_div/PartRem[6][3] , \u_div/PartRem[7][1] ,
         \u_div/PartRem[7][2] , \u_div/PartRem[7][3] , \u_div/PartRem[8][1] ,
         \u_div/PartRem[8][2] , \u_div/PartRem[8][3] , \u_div/PartRem[9][1] ,
         \u_div/PartRem[9][2] , \u_div/PartRem[9][3] , \u_div/PartRem[10][1] ,
         \u_div/PartRem[10][2] , \u_div/PartRem[11][1] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78;

  MX2X1 \u_div/u_mx_PartRem_0_1_0  ( .A(a[1]), .B(\u_div/SumTmp[1][0] ), .S0(
        quotient[1]), .Y(\u_div/PartRem[1][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_10_0  ( .A(a[10]), .B(\u_div/SumTmp[10][0] ), 
        .S0(n79), .Y(\u_div/PartRem[10][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_9_0  ( .A(a[9]), .B(\u_div/SumTmp[9][0] ), .S0(
        n80), .Y(\u_div/PartRem[9][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_0  ( .A(a[2]), .B(\u_div/SumTmp[2][0] ), .S0(
        quotient[2]), .Y(\u_div/PartRem[2][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_0  ( .A(a[4]), .B(\u_div/SumTmp[4][0] ), .S0(
        quotient[4]), .Y(\u_div/PartRem[4][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_5_0  ( .A(a[5]), .B(\u_div/SumTmp[5][0] ), .S0(
        quotient[5]), .Y(\u_div/PartRem[5][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_6_0  ( .A(a[6]), .B(\u_div/SumTmp[6][0] ), .S0(
        quotient[6]), .Y(\u_div/PartRem[6][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_7_0  ( .A(a[7]), .B(\u_div/SumTmp[7][0] ), .S0(
        quotient[7]), .Y(\u_div/PartRem[7][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_8_0  ( .A(a[8]), .B(\u_div/SumTmp[8][0] ), .S0(
        quotient[8]), .Y(\u_div/PartRem[8][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_0  ( .A(a[3]), .B(\u_div/SumTmp[3][0] ), .S0(
        quotient[3]), .Y(\u_div/PartRem[3][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_9_1  ( .A(\u_div/PartRem[10][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(n80), .Y(\u_div/PartRem[9][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/PartRem[5][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_5_1  ( .A(\u_div/PartRem[6][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_6_1  ( .A(\u_div/PartRem[7][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_7_1  ( .A(\u_div/PartRem[8][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_8_1  ( .A(\u_div/PartRem[9][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_10_1  ( .A(\u_div/PartRem[11][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(n79), .Y(\u_div/PartRem[10][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/PartRem[5][2] ), .B(
        \u_div/SumTmp[4][2] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_5_2  ( .A(\u_div/PartRem[6][2] ), .B(
        \u_div/SumTmp[5][2] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_6_2  ( .A(\u_div/PartRem[7][2] ), .B(
        \u_div/SumTmp[6][2] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_7_2  ( .A(\u_div/PartRem[8][2] ), .B(
        \u_div/SumTmp[7][2] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_8_2  ( .A(\u_div/PartRem[9][2] ), .B(
        \u_div/SumTmp[8][2] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_9_2  ( .A(\u_div/PartRem[10][2] ), .B(
        \u_div/SumTmp[9][2] ), .S0(n80), .Y(\u_div/PartRem[9][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][3] ) );
  INVX8 U1 ( .A(b[1]), .Y(n5) );
  MXI2X1 U2 ( .A(\u_div/PartRem[2][1] ), .B(\u_div/SumTmp[1][1] ), .S0(
        quotient[1]), .Y(n1) );
  OAI221X1 U3 ( .A0(n42), .A1(n10), .B0(n4), .B1(n10), .C0(n41), .Y(
        quotient[1]) );
  OAI221X1 U4 ( .A0(n46), .A1(n12), .B0(n4), .B1(n12), .C0(n45), .Y(
        quotient[2]) );
  OAI221X1 U5 ( .A0(n50), .A1(n14), .B0(n4), .B1(n14), .C0(n49), .Y(
        quotient[3]) );
  OAI221X1 U6 ( .A0(n54), .A1(n16), .B0(n4), .B1(n16), .C0(n53), .Y(
        quotient[4]) );
  OAI221X1 U7 ( .A0(n58), .A1(n18), .B0(n4), .B1(n18), .C0(n57), .Y(
        quotient[5]) );
  OAI221X1 U8 ( .A0(n62), .A1(n20), .B0(n4), .B1(n20), .C0(n61), .Y(
        quotient[6]) );
  OAI221X1 U9 ( .A0(n66), .A1(n22), .B0(n4), .B1(n22), .C0(n65), .Y(
        quotient[7]) );
  OAI221X1 U10 ( .A0(n75), .A1(n24), .B0(n4), .B1(n24), .C0(n74), .Y(
        quotient[8]) );
  OAI222X1 U11 ( .A0(n72), .A1(n25), .B0(n72), .B1(n4), .C0(n4), .C1(n25), .Y(
        n80) );
  INVXL U12 ( .A(a[11]), .Y(n38) );
  INVXL U13 ( .A(a[7]), .Y(n34) );
  INVXL U14 ( .A(a[6]), .Y(n33) );
  INVXL U15 ( .A(a[5]), .Y(n32) );
  INVXL U16 ( .A(a[4]), .Y(n31) );
  INVXL U17 ( .A(a[3]), .Y(n30) );
  INVXL U18 ( .A(a[2]), .Y(n29) );
  INVXL U19 ( .A(a[1]), .Y(n28) );
  CLKINVX3 U20 ( .A(n8), .Y(n6) );
  CLKINVX3 U21 ( .A(n8), .Y(n7) );
  INVX1 U22 ( .A(b[0]), .Y(n8) );
  INVX1 U23 ( .A(n75), .Y(n23) );
  INVX1 U24 ( .A(n66), .Y(n21) );
  INVX1 U25 ( .A(n62), .Y(n19) );
  INVX1 U26 ( .A(n58), .Y(n17) );
  INVX1 U27 ( .A(n54), .Y(n15) );
  INVX1 U28 ( .A(n50), .Y(n13) );
  INVX1 U29 ( .A(n46), .Y(n11) );
  INVX1 U30 ( .A(n42), .Y(n9) );
  INVX1 U31 ( .A(\u_div/PartRem[8][2] ), .Y(n22) );
  INVX1 U32 ( .A(\u_div/PartRem[7][2] ), .Y(n20) );
  INVX1 U33 ( .A(\u_div/PartRem[6][2] ), .Y(n18) );
  INVX1 U34 ( .A(\u_div/PartRem[5][2] ), .Y(n16) );
  INVX1 U35 ( .A(\u_div/PartRem[4][2] ), .Y(n14) );
  INVX1 U36 ( .A(\u_div/PartRem[3][2] ), .Y(n12) );
  INVX1 U37 ( .A(\u_div/PartRem[2][2] ), .Y(n10) );
  INVX1 U38 ( .A(\u_div/PartRem[9][2] ), .Y(n24) );
  INVX1 U39 ( .A(\u_div/PartRem[10][2] ), .Y(n25) );
  INVX1 U40 ( .A(n69), .Y(n26) );
  BUFX4 U41 ( .A(n27), .Y(n3) );
  INVX1 U42 ( .A(n4), .Y(n27) );
  MX2X1 U43 ( .A(\u_div/SumTmp[11][0] ), .B(a[11]), .S0(n2), .Y(
        \u_div/PartRem[11][1] ) );
  NAND3X1 U44 ( .A(n78), .B(n3), .C(n5), .Y(n2) );
  INVX1 U45 ( .A(a[10]), .Y(n37) );
  BUFX3 U46 ( .A(b[2]), .Y(n4) );
  INVX1 U47 ( .A(a[9]), .Y(n36) );
  INVX1 U48 ( .A(a[8]), .Y(n35) );
  AOI222X1 U49 ( .A0(\u_div/CryTmp[0][1] ), .A1(\u_div/PartRem[1][1] ), .B0(n5), .B1(\u_div/CryTmp[0][1] ), .C0(n5), .C1(\u_div/PartRem[1][1] ), .Y(n40) );
  AOI2BB1X1 U50 ( .A0N(n4), .A1N(n40), .B0(\u_div/PartRem[1][3] ), .Y(n39) );
  OAI221XL U51 ( .A0(n40), .A1(n1), .B0(n4), .B1(n1), .C0(n39), .Y(quotient[0]) );
  AOI222X1 U52 ( .A0(\u_div/CryTmp[1][1] ), .A1(\u_div/PartRem[2][1] ), .B0(n5), .B1(\u_div/CryTmp[1][1] ), .C0(n5), .C1(\u_div/PartRem[2][1] ), .Y(n42) );
  AOI21X1 U53 ( .A0(n3), .A1(n9), .B0(\u_div/PartRem[2][3] ), .Y(n41) );
  XOR2X1 U54 ( .A(\u_div/CryTmp[1][1] ), .B(n5), .Y(n43) );
  XOR2X1 U55 ( .A(\u_div/PartRem[2][1] ), .B(n43), .Y(\u_div/SumTmp[1][1] ) );
  XOR2X1 U56 ( .A(n10), .B(n3), .Y(n44) );
  XNOR2X1 U57 ( .A(n44), .B(n9), .Y(\u_div/SumTmp[1][2] ) );
  AOI222X1 U58 ( .A0(\u_div/CryTmp[2][1] ), .A1(\u_div/PartRem[3][1] ), .B0(n5), .B1(\u_div/CryTmp[2][1] ), .C0(n5), .C1(\u_div/PartRem[3][1] ), .Y(n46) );
  AOI21X1 U59 ( .A0(n3), .A1(n11), .B0(\u_div/PartRem[3][3] ), .Y(n45) );
  XOR2X1 U60 ( .A(\u_div/CryTmp[2][1] ), .B(n5), .Y(n47) );
  XOR2X1 U61 ( .A(\u_div/PartRem[3][1] ), .B(n47), .Y(\u_div/SumTmp[2][1] ) );
  XOR2X1 U62 ( .A(n12), .B(n3), .Y(n48) );
  XNOR2X1 U63 ( .A(n48), .B(n11), .Y(\u_div/SumTmp[2][2] ) );
  AOI222X1 U64 ( .A0(\u_div/CryTmp[3][1] ), .A1(\u_div/PartRem[4][1] ), .B0(n5), .B1(\u_div/CryTmp[3][1] ), .C0(n5), .C1(\u_div/PartRem[4][1] ), .Y(n50) );
  AOI21X1 U65 ( .A0(n3), .A1(n13), .B0(\u_div/PartRem[4][3] ), .Y(n49) );
  XOR2X1 U66 ( .A(\u_div/CryTmp[3][1] ), .B(n5), .Y(n51) );
  XOR2X1 U67 ( .A(\u_div/PartRem[4][1] ), .B(n51), .Y(\u_div/SumTmp[3][1] ) );
  XOR2X1 U68 ( .A(n14), .B(n3), .Y(n52) );
  XNOR2X1 U69 ( .A(n52), .B(n13), .Y(\u_div/SumTmp[3][2] ) );
  AOI222X1 U70 ( .A0(\u_div/CryTmp[4][1] ), .A1(\u_div/PartRem[5][1] ), .B0(n5), .B1(\u_div/CryTmp[4][1] ), .C0(n5), .C1(\u_div/PartRem[5][1] ), .Y(n54) );
  AOI21X1 U71 ( .A0(n3), .A1(n15), .B0(\u_div/PartRem[5][3] ), .Y(n53) );
  XOR2X1 U72 ( .A(\u_div/CryTmp[4][1] ), .B(n5), .Y(n55) );
  XOR2X1 U73 ( .A(\u_div/PartRem[5][1] ), .B(n55), .Y(\u_div/SumTmp[4][1] ) );
  XOR2X1 U74 ( .A(n16), .B(n3), .Y(n56) );
  XNOR2X1 U75 ( .A(n56), .B(n15), .Y(\u_div/SumTmp[4][2] ) );
  AOI222X1 U76 ( .A0(\u_div/CryTmp[5][1] ), .A1(\u_div/PartRem[6][1] ), .B0(n5), .B1(\u_div/CryTmp[5][1] ), .C0(n5), .C1(\u_div/PartRem[6][1] ), .Y(n58) );
  AOI21X1 U77 ( .A0(n3), .A1(n17), .B0(\u_div/PartRem[6][3] ), .Y(n57) );
  XOR2X1 U78 ( .A(\u_div/CryTmp[5][1] ), .B(n5), .Y(n59) );
  XOR2X1 U79 ( .A(\u_div/PartRem[6][1] ), .B(n59), .Y(\u_div/SumTmp[5][1] ) );
  XOR2X1 U80 ( .A(n18), .B(n3), .Y(n60) );
  XNOR2X1 U81 ( .A(n60), .B(n17), .Y(\u_div/SumTmp[5][2] ) );
  AOI222X1 U82 ( .A0(\u_div/CryTmp[6][1] ), .A1(\u_div/PartRem[7][1] ), .B0(n5), .B1(\u_div/CryTmp[6][1] ), .C0(n5), .C1(\u_div/PartRem[7][1] ), .Y(n62) );
  AOI21X1 U83 ( .A0(n3), .A1(n19), .B0(\u_div/PartRem[7][3] ), .Y(n61) );
  XOR2X1 U84 ( .A(\u_div/CryTmp[6][1] ), .B(n5), .Y(n63) );
  XOR2X1 U85 ( .A(\u_div/PartRem[7][1] ), .B(n63), .Y(\u_div/SumTmp[6][1] ) );
  XOR2X1 U86 ( .A(n20), .B(n3), .Y(n64) );
  XNOR2X1 U87 ( .A(n64), .B(n19), .Y(\u_div/SumTmp[6][2] ) );
  AOI222X1 U88 ( .A0(\u_div/CryTmp[7][1] ), .A1(\u_div/PartRem[8][1] ), .B0(n5), .B1(\u_div/CryTmp[7][1] ), .C0(n5), .C1(\u_div/PartRem[8][1] ), .Y(n66) );
  AOI21X1 U89 ( .A0(n3), .A1(n21), .B0(\u_div/PartRem[8][3] ), .Y(n65) );
  XOR2X1 U90 ( .A(\u_div/CryTmp[7][1] ), .B(n5), .Y(n67) );
  XOR2X1 U91 ( .A(\u_div/PartRem[8][1] ), .B(n67), .Y(\u_div/SumTmp[7][1] ) );
  XOR2X1 U92 ( .A(n22), .B(n3), .Y(n68) );
  XNOR2X1 U93 ( .A(n68), .B(n21), .Y(\u_div/SumTmp[7][2] ) );
  AOI222X1 U94 ( .A0(\u_div/CryTmp[10][1] ), .A1(\u_div/PartRem[11][1] ), .B0(
        \u_div/CryTmp[10][1] ), .B1(n5), .C0(n5), .C1(\u_div/PartRem[11][1] ), 
        .Y(n69) );
  XOR2X1 U95 ( .A(\u_div/CryTmp[10][1] ), .B(n5), .Y(n70) );
  XOR2X1 U96 ( .A(\u_div/PartRem[11][1] ), .B(n70), .Y(\u_div/SumTmp[10][1] )
         );
  AOI222X1 U97 ( .A0(\u_div/CryTmp[9][1] ), .A1(\u_div/PartRem[10][1] ), .B0(
        n5), .B1(\u_div/CryTmp[9][1] ), .C0(n5), .C1(\u_div/PartRem[10][1] ), 
        .Y(n72) );
  XOR2X1 U98 ( .A(\u_div/CryTmp[9][1] ), .B(n5), .Y(n71) );
  XOR2X1 U99 ( .A(\u_div/PartRem[10][1] ), .B(n71), .Y(\u_div/SumTmp[9][1] )
         );
  XNOR2X1 U100 ( .A(\u_div/PartRem[10][2] ), .B(n3), .Y(n73) );
  XOR2X1 U101 ( .A(n73), .B(n72), .Y(\u_div/SumTmp[9][2] ) );
  AOI222X1 U102 ( .A0(\u_div/CryTmp[8][1] ), .A1(\u_div/PartRem[9][1] ), .B0(
        n5), .B1(\u_div/CryTmp[8][1] ), .C0(n5), .C1(\u_div/PartRem[9][1] ), 
        .Y(n75) );
  AOI21X1 U103 ( .A0(n3), .A1(n23), .B0(\u_div/PartRem[9][3] ), .Y(n74) );
  XOR2X1 U104 ( .A(\u_div/CryTmp[8][1] ), .B(n5), .Y(n76) );
  XOR2X1 U105 ( .A(\u_div/PartRem[9][1] ), .B(n76), .Y(\u_div/SumTmp[8][1] )
         );
  XOR2X1 U106 ( .A(n24), .B(n3), .Y(n77) );
  XNOR2X1 U107 ( .A(n77), .B(n23), .Y(\u_div/SumTmp[8][2] ) );
  OAI21XL U108 ( .A0(n7), .A1(n36), .B0(\u_div/CryTmp[9][1] ), .Y(
        \u_div/SumTmp[9][0] ) );
  OAI21XL U109 ( .A0(n7), .A1(n35), .B0(\u_div/CryTmp[8][1] ), .Y(
        \u_div/SumTmp[8][0] ) );
  OAI21XL U110 ( .A0(n7), .A1(n34), .B0(\u_div/CryTmp[7][1] ), .Y(
        \u_div/SumTmp[7][0] ) );
  OAI21XL U111 ( .A0(n7), .A1(n33), .B0(\u_div/CryTmp[6][1] ), .Y(
        \u_div/SumTmp[6][0] ) );
  OAI21XL U112 ( .A0(n7), .A1(n32), .B0(\u_div/CryTmp[5][1] ), .Y(
        \u_div/SumTmp[5][0] ) );
  OAI21XL U113 ( .A0(n7), .A1(n31), .B0(\u_div/CryTmp[4][1] ), .Y(
        \u_div/SumTmp[4][0] ) );
  OAI21XL U114 ( .A0(n7), .A1(n30), .B0(\u_div/CryTmp[3][1] ), .Y(
        \u_div/SumTmp[3][0] ) );
  OAI21XL U115 ( .A0(n7), .A1(n29), .B0(\u_div/CryTmp[2][1] ), .Y(
        \u_div/SumTmp[2][0] ) );
  OAI21XL U116 ( .A0(n7), .A1(n28), .B0(\u_div/CryTmp[1][1] ), .Y(
        \u_div/SumTmp[1][0] ) );
  OAI21XL U117 ( .A0(n7), .A1(n38), .B0(n78), .Y(\u_div/SumTmp[11][0] ) );
  OAI21XL U118 ( .A0(n6), .A1(n37), .B0(\u_div/CryTmp[10][1] ), .Y(
        \u_div/SumTmp[10][0] ) );
  NAND2X1 U119 ( .A(n6), .B(n36), .Y(\u_div/CryTmp[9][1] ) );
  NAND2X1 U120 ( .A(n6), .B(n35), .Y(\u_div/CryTmp[8][1] ) );
  NAND2X1 U121 ( .A(n6), .B(n34), .Y(\u_div/CryTmp[7][1] ) );
  NAND2X1 U122 ( .A(n6), .B(n33), .Y(\u_div/CryTmp[6][1] ) );
  NAND2X1 U123 ( .A(n6), .B(n32), .Y(\u_div/CryTmp[5][1] ) );
  NAND2X1 U124 ( .A(n6), .B(n31), .Y(\u_div/CryTmp[4][1] ) );
  NAND2X1 U125 ( .A(n6), .B(n30), .Y(\u_div/CryTmp[3][1] ) );
  NAND2X1 U126 ( .A(n6), .B(n29), .Y(\u_div/CryTmp[2][1] ) );
  NAND2X1 U127 ( .A(n6), .B(n28), .Y(\u_div/CryTmp[1][1] ) );
  NAND2X1 U128 ( .A(n6), .B(n37), .Y(\u_div/CryTmp[10][1] ) );
  NAND2BX1 U129 ( .AN(a[0]), .B(n6), .Y(\u_div/CryTmp[0][1] ) );
  NAND2X1 U130 ( .A(n6), .B(n38), .Y(n78) );
  AND2X1 U131 ( .A(n26), .B(n3), .Y(n79) );
endmodule


module Equation_Implementation_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [12:0] carry;

  ADDFX2 U2_5 ( .A(A[5]), .B(n7), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n6), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFX2 U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFX2 U2_2 ( .A(A[2]), .B(n4), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFX2 U2_1 ( .A(A[1]), .B(n3), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(n8), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFX2 U2_7 ( .A(A[7]), .B(n9), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  INVX1 U1 ( .A(B[0]), .Y(n2) );
  INVX1 U2 ( .A(B[7]), .Y(n9) );
  OR2X2 U3 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  OR2X2 U4 ( .A(carry[8]), .B(A[8]), .Y(carry[9]) );
  XOR2X1 U5 ( .A(A[11]), .B(n1), .Y(DIFF[11]) );
  NOR2X1 U6 ( .A(carry[10]), .B(A[10]), .Y(n1) );
  INVX1 U7 ( .A(B[6]), .Y(n8) );
  INVX1 U8 ( .A(B[1]), .Y(n3) );
  OR2X2 U9 ( .A(A[0]), .B(n2), .Y(carry[1]) );
  INVX1 U10 ( .A(B[2]), .Y(n4) );
  INVX1 U11 ( .A(B[3]), .Y(n5) );
  INVX1 U12 ( .A(B[4]), .Y(n6) );
  INVX1 U13 ( .A(B[5]), .Y(n7) );
  XNOR2X1 U14 ( .A(n2), .B(A[0]), .Y(DIFF[0]) );
  XNOR2X1 U15 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  XNOR2X1 U16 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2X1 U17 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
endmodule


module Equation_Implementation_DW01_add_141 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [11:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
  AND2X2 U2 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  XOR2X1 U3 ( .A(A[9]), .B(carry[9]), .Y(SUM[9]) );
  XNOR2X1 U4 ( .A(A[11]), .B(n1), .Y(SUM[11]) );
  NAND2X1 U5 ( .A(A[10]), .B(carry[10]), .Y(n1) );
  XOR2X1 U6 ( .A(A[10]), .B(carry[10]), .Y(SUM[10]) );
  AND2X2 U7 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XOR2X1 U8 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U9 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Equation_Implementation_DW01_add_142 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [11:1] carry;

  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(A[10]), .B(carry[10]), .Y(SUM[10]) );
  XOR2X1 U3 ( .A(A[9]), .B(carry[9]), .Y(SUM[9]) );
  XOR2X1 U4 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X2 U5 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
  AND2X2 U6 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  AND2X2 U7 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XNOR2X1 U8 ( .A(A[11]), .B(n1), .Y(SUM[11]) );
  NAND2X1 U9 ( .A(A[10]), .B(carry[10]), .Y(n1) );
endmodule


module Equation_Implementation_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  CMPR22X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CMPR22X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  CMPR22X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module Equation_Implementation_DW01_sub_6 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [12:0] carry;

  ADDFX2 U2_5 ( .A(A[5]), .B(n6), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFX2 U2_3 ( .A(A[3]), .B(n4), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFX2 U2_2 ( .A(A[2]), .B(n3), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFX2 U2_1 ( .A(A[1]), .B(n2), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFX2 U2_7 ( .A(A[7]), .B(n8), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  INVX1 U1 ( .A(B[0]), .Y(n1) );
  INVX1 U2 ( .A(B[7]), .Y(n8) );
  OR2X2 U3 ( .A(carry[8]), .B(A[8]), .Y(carry[9]) );
  OR2X2 U4 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  XNOR2X1 U5 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  XNOR2X1 U6 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  XNOR2X1 U7 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  INVX1 U8 ( .A(B[6]), .Y(n7) );
  INVX1 U9 ( .A(B[1]), .Y(n2) );
  OR2X2 U10 ( .A(A[0]), .B(n1), .Y(carry[1]) );
  INVX1 U11 ( .A(B[2]), .Y(n3) );
  INVX1 U12 ( .A(B[3]), .Y(n4) );
  INVX1 U13 ( .A(B[4]), .Y(n5) );
  INVX1 U14 ( .A(B[5]), .Y(n6) );
  XNOR2X1 U15 ( .A(A[11]), .B(carry[11]), .Y(DIFF[11]) );
  OR2X2 U16 ( .A(carry[10]), .B(A[10]), .Y(carry[11]) );
  XNOR2X1 U17 ( .A(n1), .B(A[0]), .Y(DIFF[0]) );
endmodule


module Equation_Implementation_DW01_add_148 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  XOR3X2 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Y(SUM[11]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Equation_Implementation_DW01_add_147 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U3 ( .A(A[9]), .B(carry[9]), .Y(SUM[9]) );
  XOR2X1 U4 ( .A(A[10]), .B(carry[10]), .Y(SUM[10]) );
  AND2X2 U5 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
  AND2X2 U6 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  AND2X2 U7 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XOR2X1 U8 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  AND2X2 U9 ( .A(A[10]), .B(carry[10]), .Y(carry[11]) );
endmodule


module Equation_Implementation_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [12:0] carry;

  ADDFX2 U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFX2 U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFX2 U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFX2 U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFX2 U2_7 ( .A(A[7]), .B(n1), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  INVX1 U1 ( .A(B[7]), .Y(n1) );
  OR2X2 U2 ( .A(carry[8]), .B(A[8]), .Y(carry[9]) );
  OR2X2 U3 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  INVX1 U4 ( .A(B[6]), .Y(n2) );
  INVX1 U5 ( .A(B[1]), .Y(n7) );
  OR2X2 U6 ( .A(A[0]), .B(n8), .Y(carry[1]) );
  INVX1 U7 ( .A(B[4]), .Y(n4) );
  INVX1 U8 ( .A(B[5]), .Y(n3) );
  INVX1 U9 ( .A(B[2]), .Y(n6) );
  INVX1 U10 ( .A(B[3]), .Y(n5) );
  XNOR2X1 U11 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  XNOR2X1 U12 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2X1 U13 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  INVX1 U14 ( .A(B[0]), .Y(n8) );
  XNOR2X1 U15 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
  XNOR2X1 U16 ( .A(A[11]), .B(carry[11]), .Y(DIFF[11]) );
  OR2X2 U17 ( .A(carry[10]), .B(A[10]), .Y(carry[11]) );
endmodule


module Equation_Implementation_DW01_sub_9 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [12:0] carry;

  ADDFX2 U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFX2 U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFX2 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFX2 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFX2 U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFX2 U2_7 ( .A(A[7]), .B(n2), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  XNOR2X1 U1 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  XNOR2X1 U2 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2X1 U3 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  INVX1 U4 ( .A(B[7]), .Y(n2) );
  XNOR2X1 U5 ( .A(n9), .B(A[0]), .Y(DIFF[0]) );
  OR2X2 U6 ( .A(carry[8]), .B(A[8]), .Y(carry[9]) );
  OR2X2 U7 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  XOR2X1 U8 ( .A(A[11]), .B(n1), .Y(DIFF[11]) );
  NOR2X1 U9 ( .A(carry[10]), .B(A[10]), .Y(n1) );
  INVX1 U10 ( .A(B[1]), .Y(n8) );
  OR2X2 U11 ( .A(A[0]), .B(n9), .Y(carry[1]) );
  INVX1 U12 ( .A(B[2]), .Y(n7) );
  INVX1 U13 ( .A(B[3]), .Y(n6) );
  INVX1 U14 ( .A(B[4]), .Y(n5) );
  INVX1 U15 ( .A(B[5]), .Y(n4) );
  INVX1 U16 ( .A(B[6]), .Y(n3) );
  INVX1 U17 ( .A(B[0]), .Y(n9) );
endmodule


module Equation_Implementation_DW01_add_150 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  XOR3X2 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Y(SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Equation_Implementation_DW01_add_152 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;
  assign SUM[0] = B[0];

  XOR3X2 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .Y(SUM[9]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(carry[2]) );
  XOR2X1 U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module Equation_Implementation_DW_mult_uns_5 ( a, b, product );
  input [9:0] a;
  input [7:0] b;
  output [17:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259;

  ADDFX2 U2 ( .A(n17), .B(n105), .CI(n2), .CO(product[17]), .S(product[16]) );
  ADDFX2 U3 ( .A(n20), .B(n18), .CI(n3), .CO(n2), .S(product[15]) );
  ADDFX2 U4 ( .A(n23), .B(n21), .CI(n4), .CO(n3), .S(product[14]) );
  ADDFX2 U5 ( .A(n24), .B(n28), .CI(n5), .CO(n4), .S(product[13]) );
  ADDFX2 U6 ( .A(n29), .B(n34), .CI(n6), .CO(n5), .S(product[12]) );
  ADDFX2 U7 ( .A(n35), .B(n42), .CI(n7), .CO(n6), .S(product[11]) );
  ADDFX2 U8 ( .A(n43), .B(n52), .CI(n8), .CO(n7), .S(product[10]) );
  ADDFX2 U9 ( .A(n53), .B(n61), .CI(n9), .CO(n8), .S(product[9]) );
  ADDFX2 U10 ( .A(n62), .B(n70), .CI(n10), .CO(n9), .S(product[8]) );
  ADDFX2 U11 ( .A(n71), .B(n80), .CI(n11), .CO(n10), .S(product[7]) );
  ADDFX2 U12 ( .A(n81), .B(n88), .CI(n12), .CO(n11), .S(product[6]) );
  ADDFX2 U13 ( .A(n89), .B(n95), .CI(n13), .CO(n12), .S(product[5]) );
  ADDFX2 U14 ( .A(n96), .B(n99), .CI(n14), .CO(n13), .S(product[4]) );
  ADDFX2 U15 ( .A(n100), .B(n102), .CI(n15), .CO(n14), .S(product[3]) );
  ADDFX2 U16 ( .A(n16), .B(n164), .CI(n104), .CO(n15), .S(product[2]) );
  ADDHXL U17 ( .A(n174), .B(n183), .CO(n16), .S(product[1]) );
  ADDFX2 U18 ( .A(n106), .B(n115), .CI(n19), .CO(n17), .S(n18) );
  CMPR42X1 U19 ( .A(n107), .B(n125), .C(n25), .D(n116), .ICI(n22), .S(n21), 
        .ICO(n19), .CO(n20) );
  CMPR42X1 U20 ( .A(n30), .B(n117), .C(n31), .D(n26), .ICI(n27), .S(n24), 
        .ICO(n22), .CO(n23) );
  ADDFX2 U21 ( .A(n126), .B(n135), .CI(n108), .CO(n25), .S(n26) );
  CMPR42X1 U22 ( .A(n32), .B(n39), .C(n37), .D(n36), .ICI(n33), .S(n29), .ICO(
        n27), .CO(n28) );
  CMPR42X1 U23 ( .A(n109), .B(n145), .C(n136), .D(n118), .ICI(n127), .S(n32), 
        .ICO(n30), .CO(n31) );
  CMPR42X1 U24 ( .A(n44), .B(n40), .C(n45), .D(n38), .ICI(n41), .S(n35), .ICO(
        n33), .CO(n34) );
  CMPR42X1 U25 ( .A(n146), .B(n128), .C(n49), .D(n137), .ICI(n47), .S(n38), 
        .ICO(n36), .CO(n37) );
  ADDFX2 U26 ( .A(n110), .B(n155), .CI(n119), .CO(n39), .S(n40) );
  CMPR42X1 U27 ( .A(n54), .B(n58), .C(n46), .D(n55), .ICI(n51), .S(n43), .ICO(
        n41), .CO(n42) );
  CMPR42X1 U28 ( .A(n156), .B(n147), .C(n48), .D(n57), .ICI(n50), .S(n46), 
        .ICO(n44), .CO(n45) );
  ADDFX2 U29 ( .A(n129), .B(n138), .CI(n165), .CO(n47), .S(n48) );
  ADDHXL U30 ( .A(n120), .B(n111), .CO(n49), .S(n50) );
  CMPR42X1 U31 ( .A(n63), .B(n59), .C(n56), .D(n64), .ICI(n60), .S(n53), .ICO(
        n51), .CO(n52) );
  CMPR42X1 U32 ( .A(n175), .B(n157), .C(n66), .D(n166), .ICI(n67), .S(n56), 
        .ICO(n54), .CO(n55) );
  CMPR42X1 U33 ( .A(n112), .B(n121), .C(n139), .D(n130), .ICI(n148), .S(n59), 
        .ICO(n57), .CO(n58) );
  CMPR42X1 U34 ( .A(n72), .B(n68), .C(n65), .D(n73), .ICI(n69), .S(n62), .ICO(
        n60), .CO(n61) );
  CMPR42X1 U35 ( .A(n176), .B(n158), .C(n77), .D(n167), .ICI(n75), .S(n65), 
        .ICO(n63), .CO(n64) );
  CMPR42X1 U36 ( .A(n113), .B(n122), .C(n140), .D(n131), .ICI(n149), .S(n68), 
        .ICO(n66), .CO(n67) );
  CMPR42X1 U37 ( .A(n78), .B(n76), .C(n74), .D(n83), .ICI(n79), .S(n71), .ICO(
        n69), .CO(n70) );
  CMPR42X1 U38 ( .A(n168), .B(n141), .C(n82), .D(n159), .ICI(n85), .S(n74), 
        .ICO(n72), .CO(n73) );
  ADDFX2 U39 ( .A(n177), .B(n150), .CI(n132), .CO(n75), .S(n76) );
  ADDHXL U40 ( .A(n123), .B(n114), .CO(n77), .S(n78) );
  CMPR42X1 U41 ( .A(n90), .B(n92), .C(n84), .D(n86), .ICI(n87), .S(n81), .ICO(
        n79), .CO(n80) );
  CMPR42X1 U42 ( .A(n142), .B(n178), .C(n160), .D(n151), .ICI(n169), .S(n84), 
        .ICO(n82), .CO(n83) );
  ADDHXL U43 ( .A(n133), .B(n124), .CO(n85), .S(n86) );
  CMPR42X1 U44 ( .A(n97), .B(n170), .C(n93), .D(n91), .ICI(n94), .S(n89), 
        .ICO(n87), .CO(n88) );
  ADDFX2 U45 ( .A(n152), .B(n179), .CI(n161), .CO(n90), .S(n91) );
  ADDHXL U46 ( .A(n143), .B(n134), .CO(n92), .S(n93) );
  CMPR42X1 U47 ( .A(n162), .B(n180), .C(n101), .D(n171), .ICI(n98), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDHXL U48 ( .A(n153), .B(n144), .CO(n97), .S(n98) );
  ADDFX2 U49 ( .A(n172), .B(n181), .CI(n103), .CO(n99), .S(n100) );
  ADDHXL U50 ( .A(n163), .B(n154), .CO(n101), .S(n102) );
  ADDHXL U51 ( .A(n182), .B(n173), .CO(n103), .S(n104) );
  CLKINVX3 U152 ( .A(b[0]), .Y(n249) );
  CLKINVX3 U153 ( .A(b[1]), .Y(n248) );
  CLKINVX3 U154 ( .A(b[3]), .Y(n246) );
  CLKINVX3 U155 ( .A(b[2]), .Y(n247) );
  CLKINVX3 U156 ( .A(b[4]), .Y(n245) );
  CLKINVX3 U157 ( .A(b[7]), .Y(n242) );
  CLKINVX3 U158 ( .A(b[5]), .Y(n244) );
  CLKINVX3 U159 ( .A(b[6]), .Y(n243) );
  CLKINVX3 U160 ( .A(a[0]), .Y(n259) );
  CLKINVX3 U161 ( .A(a[1]), .Y(n258) );
  CLKINVX3 U162 ( .A(a[2]), .Y(n257) );
  CLKINVX3 U163 ( .A(a[3]), .Y(n256) );
  CLKINVX3 U164 ( .A(a[4]), .Y(n255) );
  CLKINVX3 U165 ( .A(a[5]), .Y(n254) );
  CLKINVX3 U166 ( .A(a[6]), .Y(n253) );
  CLKINVX3 U167 ( .A(a[7]), .Y(n252) );
  CLKINVX3 U168 ( .A(a[9]), .Y(n250) );
  CLKINVX3 U169 ( .A(a[8]), .Y(n251) );
  NOR2X1 U170 ( .A(n259), .B(n249), .Y(product[0]) );
  NOR2X1 U171 ( .A(n249), .B(n258), .Y(n183) );
  NOR2X1 U172 ( .A(n249), .B(n257), .Y(n182) );
  NOR2X1 U173 ( .A(n249), .B(n256), .Y(n181) );
  NOR2X1 U174 ( .A(n249), .B(n255), .Y(n180) );
  NOR2X1 U175 ( .A(n249), .B(n254), .Y(n179) );
  NOR2X1 U176 ( .A(n249), .B(n253), .Y(n178) );
  NOR2X1 U177 ( .A(n249), .B(n252), .Y(n177) );
  NOR2X1 U178 ( .A(n249), .B(n251), .Y(n176) );
  NOR2X1 U179 ( .A(n249), .B(n250), .Y(n175) );
  NOR2X1 U180 ( .A(n259), .B(n248), .Y(n174) );
  NOR2X1 U181 ( .A(n258), .B(n248), .Y(n173) );
  NOR2X1 U182 ( .A(n257), .B(n248), .Y(n172) );
  NOR2X1 U183 ( .A(n256), .B(n248), .Y(n171) );
  NOR2X1 U184 ( .A(n255), .B(n248), .Y(n170) );
  NOR2X1 U185 ( .A(n254), .B(n248), .Y(n169) );
  NOR2X1 U186 ( .A(n253), .B(n248), .Y(n168) );
  NOR2X1 U187 ( .A(n252), .B(n248), .Y(n167) );
  NOR2X1 U188 ( .A(n251), .B(n248), .Y(n166) );
  NOR2X1 U189 ( .A(n250), .B(n248), .Y(n165) );
  NOR2X1 U190 ( .A(n259), .B(n247), .Y(n164) );
  NOR2X1 U191 ( .A(n258), .B(n247), .Y(n163) );
  NOR2X1 U192 ( .A(n257), .B(n247), .Y(n162) );
  NOR2X1 U193 ( .A(n256), .B(n247), .Y(n161) );
  NOR2X1 U194 ( .A(n255), .B(n247), .Y(n160) );
  NOR2X1 U195 ( .A(n254), .B(n247), .Y(n159) );
  NOR2X1 U196 ( .A(n253), .B(n247), .Y(n158) );
  NOR2X1 U197 ( .A(n252), .B(n247), .Y(n157) );
  NOR2X1 U198 ( .A(n251), .B(n247), .Y(n156) );
  NOR2X1 U199 ( .A(n250), .B(n247), .Y(n155) );
  NOR2X1 U200 ( .A(n259), .B(n246), .Y(n154) );
  NOR2X1 U201 ( .A(n258), .B(n246), .Y(n153) );
  NOR2X1 U202 ( .A(n257), .B(n246), .Y(n152) );
  NOR2X1 U203 ( .A(n256), .B(n246), .Y(n151) );
  NOR2X1 U204 ( .A(n255), .B(n246), .Y(n150) );
  NOR2X1 U205 ( .A(n254), .B(n246), .Y(n149) );
  NOR2X1 U206 ( .A(n253), .B(n246), .Y(n148) );
  NOR2X1 U207 ( .A(n252), .B(n246), .Y(n147) );
  NOR2X1 U208 ( .A(n251), .B(n246), .Y(n146) );
  NOR2X1 U209 ( .A(n250), .B(n246), .Y(n145) );
  NOR2X1 U210 ( .A(n259), .B(n245), .Y(n144) );
  NOR2X1 U211 ( .A(n258), .B(n245), .Y(n143) );
  NOR2X1 U212 ( .A(n257), .B(n245), .Y(n142) );
  NOR2X1 U213 ( .A(n256), .B(n245), .Y(n141) );
  NOR2X1 U214 ( .A(n255), .B(n245), .Y(n140) );
  NOR2X1 U215 ( .A(n254), .B(n245), .Y(n139) );
  NOR2X1 U216 ( .A(n253), .B(n245), .Y(n138) );
  NOR2X1 U217 ( .A(n252), .B(n245), .Y(n137) );
  NOR2X1 U218 ( .A(n251), .B(n245), .Y(n136) );
  NOR2X1 U219 ( .A(n250), .B(n245), .Y(n135) );
  NOR2X1 U220 ( .A(n259), .B(n244), .Y(n134) );
  NOR2X1 U221 ( .A(n258), .B(n244), .Y(n133) );
  NOR2X1 U222 ( .A(n257), .B(n244), .Y(n132) );
  NOR2X1 U223 ( .A(n256), .B(n244), .Y(n131) );
  NOR2X1 U224 ( .A(n255), .B(n244), .Y(n130) );
  NOR2X1 U225 ( .A(n254), .B(n244), .Y(n129) );
  NOR2X1 U226 ( .A(n253), .B(n244), .Y(n128) );
  NOR2X1 U227 ( .A(n252), .B(n244), .Y(n127) );
  NOR2X1 U228 ( .A(n251), .B(n244), .Y(n126) );
  NOR2X1 U229 ( .A(n250), .B(n244), .Y(n125) );
  NOR2X1 U230 ( .A(n259), .B(n243), .Y(n124) );
  NOR2X1 U231 ( .A(n258), .B(n243), .Y(n123) );
  NOR2X1 U232 ( .A(n257), .B(n243), .Y(n122) );
  NOR2X1 U233 ( .A(n256), .B(n243), .Y(n121) );
  NOR2X1 U234 ( .A(n255), .B(n243), .Y(n120) );
  NOR2X1 U235 ( .A(n254), .B(n243), .Y(n119) );
  NOR2X1 U236 ( .A(n253), .B(n243), .Y(n118) );
  NOR2X1 U237 ( .A(n252), .B(n243), .Y(n117) );
  NOR2X1 U238 ( .A(n251), .B(n243), .Y(n116) );
  NOR2X1 U239 ( .A(n250), .B(n243), .Y(n115) );
  NOR2X1 U240 ( .A(n259), .B(n242), .Y(n114) );
  NOR2X1 U241 ( .A(n258), .B(n242), .Y(n113) );
  NOR2X1 U242 ( .A(n257), .B(n242), .Y(n112) );
  NOR2X1 U243 ( .A(n256), .B(n242), .Y(n111) );
  NOR2X1 U244 ( .A(n255), .B(n242), .Y(n110) );
  NOR2X1 U245 ( .A(n254), .B(n242), .Y(n109) );
  NOR2X1 U246 ( .A(n253), .B(n242), .Y(n108) );
  NOR2X1 U247 ( .A(n252), .B(n242), .Y(n107) );
  NOR2X1 U248 ( .A(n251), .B(n242), .Y(n106) );
  NOR2X1 U249 ( .A(n250), .B(n242), .Y(n105) );
endmodule


module Equation_Implementation_DW_mult_uns_4 ( a, b, product );
  input [9:0] a;
  input [7:0] b;
  output [17:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259;

  ADDFX2 U2 ( .A(n17), .B(n105), .CI(n2), .CO(product[17]), .S(product[16]) );
  ADDFX2 U3 ( .A(n20), .B(n18), .CI(n3), .CO(n2), .S(product[15]) );
  ADDFX2 U4 ( .A(n23), .B(n21), .CI(n4), .CO(n3), .S(product[14]) );
  ADDFX2 U5 ( .A(n24), .B(n28), .CI(n5), .CO(n4), .S(product[13]) );
  ADDFX2 U6 ( .A(n29), .B(n34), .CI(n6), .CO(n5), .S(product[12]) );
  ADDFX2 U7 ( .A(n35), .B(n42), .CI(n7), .CO(n6), .S(product[11]) );
  ADDFX2 U8 ( .A(n43), .B(n52), .CI(n8), .CO(n7), .S(product[10]) );
  ADDFX2 U9 ( .A(n53), .B(n61), .CI(n9), .CO(n8), .S(product[9]) );
  ADDFX2 U10 ( .A(n62), .B(n70), .CI(n10), .CO(n9), .S(product[8]) );
  ADDFX2 U11 ( .A(n71), .B(n80), .CI(n11), .CO(n10), .S(product[7]) );
  ADDFX2 U12 ( .A(n81), .B(n88), .CI(n12), .CO(n11), .S(product[6]) );
  ADDFX2 U13 ( .A(n89), .B(n95), .CI(n13), .CO(n12), .S(product[5]) );
  ADDFX2 U14 ( .A(n96), .B(n99), .CI(n14), .CO(n13), .S(product[4]) );
  ADDFX2 U15 ( .A(n100), .B(n102), .CI(n15), .CO(n14), .S(product[3]) );
  ADDFX2 U16 ( .A(n16), .B(n164), .CI(n104), .CO(n15), .S(product[2]) );
  ADDHXL U17 ( .A(n174), .B(n183), .CO(n16), .S(product[1]) );
  ADDFX2 U18 ( .A(n106), .B(n115), .CI(n19), .CO(n17), .S(n18) );
  CMPR42X1 U19 ( .A(n107), .B(n125), .C(n25), .D(n116), .ICI(n22), .S(n21), 
        .ICO(n19), .CO(n20) );
  CMPR42X1 U20 ( .A(n30), .B(n117), .C(n31), .D(n26), .ICI(n27), .S(n24), 
        .ICO(n22), .CO(n23) );
  ADDFX2 U21 ( .A(n126), .B(n135), .CI(n108), .CO(n25), .S(n26) );
  CMPR42X1 U22 ( .A(n32), .B(n39), .C(n37), .D(n36), .ICI(n33), .S(n29), .ICO(
        n27), .CO(n28) );
  CMPR42X1 U23 ( .A(n109), .B(n145), .C(n136), .D(n118), .ICI(n127), .S(n32), 
        .ICO(n30), .CO(n31) );
  CMPR42X1 U24 ( .A(n44), .B(n40), .C(n45), .D(n38), .ICI(n41), .S(n35), .ICO(
        n33), .CO(n34) );
  CMPR42X1 U25 ( .A(n146), .B(n128), .C(n49), .D(n137), .ICI(n47), .S(n38), 
        .ICO(n36), .CO(n37) );
  ADDFX2 U26 ( .A(n110), .B(n155), .CI(n119), .CO(n39), .S(n40) );
  CMPR42X1 U27 ( .A(n54), .B(n58), .C(n46), .D(n55), .ICI(n51), .S(n43), .ICO(
        n41), .CO(n42) );
  CMPR42X1 U28 ( .A(n156), .B(n147), .C(n48), .D(n57), .ICI(n50), .S(n46), 
        .ICO(n44), .CO(n45) );
  ADDFX2 U29 ( .A(n129), .B(n138), .CI(n165), .CO(n47), .S(n48) );
  ADDHXL U30 ( .A(n120), .B(n111), .CO(n49), .S(n50) );
  CMPR42X1 U31 ( .A(n63), .B(n59), .C(n56), .D(n64), .ICI(n60), .S(n53), .ICO(
        n51), .CO(n52) );
  CMPR42X1 U32 ( .A(n175), .B(n157), .C(n66), .D(n166), .ICI(n67), .S(n56), 
        .ICO(n54), .CO(n55) );
  CMPR42X1 U33 ( .A(n112), .B(n121), .C(n139), .D(n130), .ICI(n148), .S(n59), 
        .ICO(n57), .CO(n58) );
  CMPR42X1 U34 ( .A(n72), .B(n68), .C(n65), .D(n73), .ICI(n69), .S(n62), .ICO(
        n60), .CO(n61) );
  CMPR42X1 U35 ( .A(n176), .B(n158), .C(n77), .D(n167), .ICI(n75), .S(n65), 
        .ICO(n63), .CO(n64) );
  CMPR42X1 U36 ( .A(n113), .B(n122), .C(n140), .D(n131), .ICI(n149), .S(n68), 
        .ICO(n66), .CO(n67) );
  CMPR42X1 U37 ( .A(n78), .B(n76), .C(n74), .D(n83), .ICI(n79), .S(n71), .ICO(
        n69), .CO(n70) );
  CMPR42X1 U38 ( .A(n168), .B(n141), .C(n82), .D(n159), .ICI(n85), .S(n74), 
        .ICO(n72), .CO(n73) );
  ADDFX2 U39 ( .A(n177), .B(n150), .CI(n132), .CO(n75), .S(n76) );
  ADDHXL U40 ( .A(n123), .B(n114), .CO(n77), .S(n78) );
  CMPR42X1 U41 ( .A(n90), .B(n92), .C(n84), .D(n86), .ICI(n87), .S(n81), .ICO(
        n79), .CO(n80) );
  CMPR42X1 U42 ( .A(n142), .B(n178), .C(n160), .D(n151), .ICI(n169), .S(n84), 
        .ICO(n82), .CO(n83) );
  ADDHXL U43 ( .A(n133), .B(n124), .CO(n85), .S(n86) );
  CMPR42X1 U44 ( .A(n97), .B(n170), .C(n93), .D(n91), .ICI(n94), .S(n89), 
        .ICO(n87), .CO(n88) );
  ADDFX2 U45 ( .A(n152), .B(n179), .CI(n161), .CO(n90), .S(n91) );
  ADDHXL U46 ( .A(n143), .B(n134), .CO(n92), .S(n93) );
  CMPR42X1 U47 ( .A(n162), .B(n180), .C(n101), .D(n171), .ICI(n98), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDHXL U48 ( .A(n153), .B(n144), .CO(n97), .S(n98) );
  ADDFX2 U49 ( .A(n172), .B(n181), .CI(n103), .CO(n99), .S(n100) );
  ADDHXL U50 ( .A(n163), .B(n154), .CO(n101), .S(n102) );
  ADDHXL U51 ( .A(n182), .B(n173), .CO(n103), .S(n104) );
  CLKINVX3 U152 ( .A(b[0]), .Y(n249) );
  CLKINVX3 U153 ( .A(b[1]), .Y(n248) );
  CLKINVX3 U154 ( .A(b[3]), .Y(n246) );
  CLKINVX3 U155 ( .A(b[2]), .Y(n247) );
  CLKINVX3 U156 ( .A(b[4]), .Y(n245) );
  CLKINVX3 U157 ( .A(b[5]), .Y(n244) );
  CLKINVX3 U158 ( .A(b[6]), .Y(n243) );
  CLKINVX3 U159 ( .A(b[7]), .Y(n242) );
  CLKINVX3 U160 ( .A(a[0]), .Y(n259) );
  CLKINVX3 U161 ( .A(a[1]), .Y(n258) );
  CLKINVX3 U162 ( .A(a[2]), .Y(n257) );
  CLKINVX3 U163 ( .A(a[3]), .Y(n256) );
  CLKINVX3 U164 ( .A(a[4]), .Y(n255) );
  CLKINVX3 U165 ( .A(a[5]), .Y(n254) );
  CLKINVX3 U166 ( .A(a[6]), .Y(n253) );
  CLKINVX3 U167 ( .A(a[7]), .Y(n252) );
  CLKINVX3 U168 ( .A(a[9]), .Y(n250) );
  CLKINVX3 U169 ( .A(a[8]), .Y(n251) );
  NOR2X1 U170 ( .A(n259), .B(n249), .Y(product[0]) );
  NOR2X1 U171 ( .A(n249), .B(n258), .Y(n183) );
  NOR2X1 U172 ( .A(n249), .B(n257), .Y(n182) );
  NOR2X1 U173 ( .A(n249), .B(n256), .Y(n181) );
  NOR2X1 U174 ( .A(n249), .B(n255), .Y(n180) );
  NOR2X1 U175 ( .A(n249), .B(n254), .Y(n179) );
  NOR2X1 U176 ( .A(n249), .B(n253), .Y(n178) );
  NOR2X1 U177 ( .A(n249), .B(n252), .Y(n177) );
  NOR2X1 U178 ( .A(n249), .B(n251), .Y(n176) );
  NOR2X1 U179 ( .A(n249), .B(n250), .Y(n175) );
  NOR2X1 U180 ( .A(n259), .B(n248), .Y(n174) );
  NOR2X1 U181 ( .A(n258), .B(n248), .Y(n173) );
  NOR2X1 U182 ( .A(n257), .B(n248), .Y(n172) );
  NOR2X1 U183 ( .A(n256), .B(n248), .Y(n171) );
  NOR2X1 U184 ( .A(n255), .B(n248), .Y(n170) );
  NOR2X1 U185 ( .A(n254), .B(n248), .Y(n169) );
  NOR2X1 U186 ( .A(n253), .B(n248), .Y(n168) );
  NOR2X1 U187 ( .A(n252), .B(n248), .Y(n167) );
  NOR2X1 U188 ( .A(n251), .B(n248), .Y(n166) );
  NOR2X1 U189 ( .A(n250), .B(n248), .Y(n165) );
  NOR2X1 U190 ( .A(n259), .B(n247), .Y(n164) );
  NOR2X1 U191 ( .A(n258), .B(n247), .Y(n163) );
  NOR2X1 U192 ( .A(n257), .B(n247), .Y(n162) );
  NOR2X1 U193 ( .A(n256), .B(n247), .Y(n161) );
  NOR2X1 U194 ( .A(n255), .B(n247), .Y(n160) );
  NOR2X1 U195 ( .A(n254), .B(n247), .Y(n159) );
  NOR2X1 U196 ( .A(n253), .B(n247), .Y(n158) );
  NOR2X1 U197 ( .A(n252), .B(n247), .Y(n157) );
  NOR2X1 U198 ( .A(n251), .B(n247), .Y(n156) );
  NOR2X1 U199 ( .A(n250), .B(n247), .Y(n155) );
  NOR2X1 U200 ( .A(n259), .B(n246), .Y(n154) );
  NOR2X1 U201 ( .A(n258), .B(n246), .Y(n153) );
  NOR2X1 U202 ( .A(n257), .B(n246), .Y(n152) );
  NOR2X1 U203 ( .A(n256), .B(n246), .Y(n151) );
  NOR2X1 U204 ( .A(n255), .B(n246), .Y(n150) );
  NOR2X1 U205 ( .A(n254), .B(n246), .Y(n149) );
  NOR2X1 U206 ( .A(n253), .B(n246), .Y(n148) );
  NOR2X1 U207 ( .A(n252), .B(n246), .Y(n147) );
  NOR2X1 U208 ( .A(n251), .B(n246), .Y(n146) );
  NOR2X1 U209 ( .A(n250), .B(n246), .Y(n145) );
  NOR2X1 U210 ( .A(n259), .B(n245), .Y(n144) );
  NOR2X1 U211 ( .A(n258), .B(n245), .Y(n143) );
  NOR2X1 U212 ( .A(n257), .B(n245), .Y(n142) );
  NOR2X1 U213 ( .A(n256), .B(n245), .Y(n141) );
  NOR2X1 U214 ( .A(n255), .B(n245), .Y(n140) );
  NOR2X1 U215 ( .A(n254), .B(n245), .Y(n139) );
  NOR2X1 U216 ( .A(n253), .B(n245), .Y(n138) );
  NOR2X1 U217 ( .A(n252), .B(n245), .Y(n137) );
  NOR2X1 U218 ( .A(n251), .B(n245), .Y(n136) );
  NOR2X1 U219 ( .A(n250), .B(n245), .Y(n135) );
  NOR2X1 U220 ( .A(n259), .B(n244), .Y(n134) );
  NOR2X1 U221 ( .A(n258), .B(n244), .Y(n133) );
  NOR2X1 U222 ( .A(n257), .B(n244), .Y(n132) );
  NOR2X1 U223 ( .A(n256), .B(n244), .Y(n131) );
  NOR2X1 U224 ( .A(n255), .B(n244), .Y(n130) );
  NOR2X1 U225 ( .A(n254), .B(n244), .Y(n129) );
  NOR2X1 U226 ( .A(n253), .B(n244), .Y(n128) );
  NOR2X1 U227 ( .A(n252), .B(n244), .Y(n127) );
  NOR2X1 U228 ( .A(n251), .B(n244), .Y(n126) );
  NOR2X1 U229 ( .A(n250), .B(n244), .Y(n125) );
  NOR2X1 U230 ( .A(n259), .B(n243), .Y(n124) );
  NOR2X1 U231 ( .A(n258), .B(n243), .Y(n123) );
  NOR2X1 U232 ( .A(n257), .B(n243), .Y(n122) );
  NOR2X1 U233 ( .A(n256), .B(n243), .Y(n121) );
  NOR2X1 U234 ( .A(n255), .B(n243), .Y(n120) );
  NOR2X1 U235 ( .A(n254), .B(n243), .Y(n119) );
  NOR2X1 U236 ( .A(n253), .B(n243), .Y(n118) );
  NOR2X1 U237 ( .A(n252), .B(n243), .Y(n117) );
  NOR2X1 U238 ( .A(n251), .B(n243), .Y(n116) );
  NOR2X1 U239 ( .A(n250), .B(n243), .Y(n115) );
  NOR2X1 U240 ( .A(n259), .B(n242), .Y(n114) );
  NOR2X1 U241 ( .A(n258), .B(n242), .Y(n113) );
  NOR2X1 U242 ( .A(n257), .B(n242), .Y(n112) );
  NOR2X1 U243 ( .A(n256), .B(n242), .Y(n111) );
  NOR2X1 U244 ( .A(n255), .B(n242), .Y(n110) );
  NOR2X1 U245 ( .A(n254), .B(n242), .Y(n109) );
  NOR2X1 U246 ( .A(n253), .B(n242), .Y(n108) );
  NOR2X1 U247 ( .A(n252), .B(n242), .Y(n107) );
  NOR2X1 U248 ( .A(n251), .B(n242), .Y(n106) );
  NOR2X1 U249 ( .A(n250), .B(n242), .Y(n105) );
endmodule


module Equation_Implementation_DW01_add_143 ( A, B, CI, SUM, CO );
  input [18:0] A;
  input [18:0] B;
  output [18:0] SUM;
  input CI;
  output CO;

  wire   [18:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(SUM[18]), .S(
        SUM[17]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module Equation_Implementation_DW01_inc_1 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
endmodule


module Equation_Implementation_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [9:0] carry;

  ADDFX2 U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFX2 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFX2 U2_7 ( .A(A[7]), .B(n2), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADDFX2 U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFX2 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  INVX1 U1 ( .A(carry[8]), .Y(DIFF[8]) );
  INVX1 U2 ( .A(B[2]), .Y(n7) );
  INVX1 U3 ( .A(B[5]), .Y(n4) );
  INVX1 U4 ( .A(B[7]), .Y(n2) );
  INVX1 U5 ( .A(B[0]), .Y(n9) );
  INVX1 U6 ( .A(B[3]), .Y(n6) );
  INVX1 U7 ( .A(B[4]), .Y(n5) );
  INVX1 U8 ( .A(B[6]), .Y(n3) );
  INVX1 U9 ( .A(B[1]), .Y(n8) );
  OR2X2 U10 ( .A(A[0]), .B(n9), .Y(carry[1]) );
  XNOR2X1 U11 ( .A(n9), .B(A[0]), .Y(DIFF[0]) );
endmodule


module Equation_Implementation_DW01_add_146 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  XOR3X2 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Y(SUM[11]) );
  XOR2XL U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module Equation_Implementation_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [9:0] carry;

  ADDFX2 U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFX2 U2_7 ( .A(A[7]), .B(n2), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFX2 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFX2 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFX2 U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  INVX1 U1 ( .A(carry[8]), .Y(DIFF[8]) );
  XNOR2X1 U2 ( .A(n9), .B(A[0]), .Y(DIFF[0]) );
  INVX1 U3 ( .A(B[6]), .Y(n3) );
  INVX1 U4 ( .A(B[5]), .Y(n4) );
  INVX1 U5 ( .A(B[2]), .Y(n7) );
  INVX1 U6 ( .A(B[3]), .Y(n6) );
  INVX1 U7 ( .A(B[4]), .Y(n5) );
  INVX1 U8 ( .A(B[7]), .Y(n2) );
  INVX1 U9 ( .A(B[1]), .Y(n8) );
  OR2X2 U10 ( .A(A[0]), .B(n9), .Y(carry[1]) );
  INVX1 U11 ( .A(B[0]), .Y(n9) );
endmodule


module Equation_Implementation_DW01_add_145 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  XOR3X2 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Y(SUM[11]) );
  XOR2XL U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module Equation_Implementation_DW_mult_uns_7 ( a, b, product );
  input [6:0] a;
  input [7:0] b;
  output [14:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190;

  ADDFX2 U2 ( .A(n14), .B(n72), .CI(n2), .CO(product[14]), .S(product[13]) );
  ADDFX2 U3 ( .A(n17), .B(n15), .CI(n3), .CO(n2), .S(product[12]) );
  ADDFX2 U4 ( .A(n18), .B(n20), .CI(n4), .CO(n3), .S(product[11]) );
  ADDFX2 U5 ( .A(n21), .B(n25), .CI(n5), .CO(n4), .S(product[10]) );
  ADDFX2 U6 ( .A(n26), .B(n31), .CI(n6), .CO(n5), .S(product[9]) );
  ADDFX2 U7 ( .A(n32), .B(n39), .CI(n7), .CO(n6), .S(product[8]) );
  ADDFX2 U8 ( .A(n40), .B(n47), .CI(n8), .CO(n7), .S(product[7]) );
  ADDFX2 U9 ( .A(n48), .B(n55), .CI(n9), .CO(n8), .S(product[6]) );
  ADDFX2 U10 ( .A(n56), .B(n62), .CI(n10), .CO(n9), .S(product[5]) );
  ADDFX2 U11 ( .A(n63), .B(n66), .CI(n11), .CO(n10), .S(product[4]) );
  ADDFX2 U12 ( .A(n67), .B(n69), .CI(n12), .CO(n11), .S(product[3]) );
  ADDFX2 U13 ( .A(n13), .B(n111), .CI(n71), .CO(n12), .S(product[2]) );
  ADDHXL U14 ( .A(n119), .B(n126), .CO(n13), .S(product[1]) );
  ADDFX2 U15 ( .A(n73), .B(n80), .CI(n16), .CO(n14), .S(n15) );
  CMPR42X1 U16 ( .A(n74), .B(n88), .C(n22), .D(n81), .ICI(n19), .S(n18), .ICO(
        n16), .CO(n17) );
  CMPR42X1 U17 ( .A(n27), .B(n82), .C(n28), .D(n23), .ICI(n24), .S(n21), .ICO(
        n19), .CO(n20) );
  ADDFX2 U18 ( .A(n89), .B(n96), .CI(n75), .CO(n22), .S(n23) );
  CMPR42X1 U19 ( .A(n36), .B(n33), .C(n34), .D(n29), .ICI(n30), .S(n26), .ICO(
        n24), .CO(n25) );
  CMPR42X1 U20 ( .A(n76), .B(n90), .C(n97), .D(n104), .ICI(n83), .S(n29), 
        .ICO(n27), .CO(n28) );
  CMPR42X1 U21 ( .A(n37), .B(n44), .C(n35), .D(n42), .ICI(n38), .S(n32), .ICO(
        n30), .CO(n31) );
  CMPR42X1 U22 ( .A(n105), .B(n91), .C(n77), .D(n98), .ICI(n41), .S(n35), 
        .ICO(n33), .CO(n34) );
  ADDHXL U23 ( .A(n84), .B(n112), .CO(n36), .S(n37) );
  CMPR42X1 U24 ( .A(n45), .B(n52), .C(n43), .D(n50), .ICI(n46), .S(n40), .ICO(
        n38), .CO(n39) );
  CMPR42X1 U25 ( .A(n113), .B(n99), .C(n92), .D(n106), .ICI(n49), .S(n43), 
        .ICO(n41), .CO(n42) );
  ADDFX2 U26 ( .A(n78), .B(n85), .CI(n120), .CO(n44), .S(n45) );
  CMPR42X1 U27 ( .A(n57), .B(n59), .C(n51), .D(n53), .ICI(n54), .S(n48), .ICO(
        n46), .CO(n47) );
  CMPR42X1 U28 ( .A(n93), .B(n121), .C(n107), .D(n100), .ICI(n114), .S(n51), 
        .ICO(n49), .CO(n50) );
  ADDHXL U29 ( .A(n86), .B(n79), .CO(n52), .S(n53) );
  CMPR42X1 U30 ( .A(n64), .B(n115), .C(n60), .D(n58), .ICI(n61), .S(n56), 
        .ICO(n54), .CO(n55) );
  ADDFX2 U31 ( .A(n101), .B(n122), .CI(n108), .CO(n57), .S(n58) );
  ADDHXL U32 ( .A(n94), .B(n87), .CO(n59), .S(n60) );
  CMPR42X1 U33 ( .A(n109), .B(n123), .C(n68), .D(n116), .ICI(n65), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDHXL U34 ( .A(n102), .B(n95), .CO(n64), .S(n65) );
  ADDFX2 U35 ( .A(n117), .B(n124), .CI(n70), .CO(n66), .S(n67) );
  ADDHXL U36 ( .A(n110), .B(n103), .CO(n68), .S(n69) );
  ADDHXL U37 ( .A(n125), .B(n118), .CO(n70), .S(n71) );
  CLKINVX3 U111 ( .A(b[0]), .Y(n190) );
  CLKINVX3 U112 ( .A(b[1]), .Y(n189) );
  CLKINVX3 U113 ( .A(b[2]), .Y(n188) );
  CLKINVX3 U114 ( .A(b[4]), .Y(n186) );
  CLKINVX3 U115 ( .A(b[5]), .Y(n185) );
  CLKINVX3 U116 ( .A(b[6]), .Y(n184) );
  CLKINVX3 U117 ( .A(b[3]), .Y(n187) );
  CLKINVX3 U118 ( .A(b[7]), .Y(n183) );
  CLKINVX3 U119 ( .A(a[0]), .Y(n182) );
  CLKINVX3 U120 ( .A(a[3]), .Y(n179) );
  CLKINVX3 U121 ( .A(a[4]), .Y(n178) );
  CLKINVX3 U122 ( .A(a[1]), .Y(n181) );
  CLKINVX3 U123 ( .A(a[2]), .Y(n180) );
  CLKINVX3 U124 ( .A(a[5]), .Y(n177) );
  CLKINVX3 U125 ( .A(a[6]), .Y(n176) );
  NOR2X1 U126 ( .A(n182), .B(n190), .Y(product[0]) );
  NOR2X1 U127 ( .A(n179), .B(n186), .Y(n99) );
  NOR2X1 U128 ( .A(n179), .B(n185), .Y(n98) );
  NOR2X1 U129 ( .A(n179), .B(n184), .Y(n97) );
  NOR2X1 U130 ( .A(n179), .B(n183), .Y(n96) );
  NOR2X1 U131 ( .A(n190), .B(n178), .Y(n95) );
  NOR2X1 U132 ( .A(n178), .B(n189), .Y(n94) );
  NOR2X1 U133 ( .A(n178), .B(n188), .Y(n93) );
  NOR2X1 U134 ( .A(n178), .B(n187), .Y(n92) );
  NOR2X1 U135 ( .A(n186), .B(n178), .Y(n91) );
  NOR2X1 U136 ( .A(n185), .B(n178), .Y(n90) );
  NOR2X1 U137 ( .A(n184), .B(n178), .Y(n89) );
  NOR2X1 U138 ( .A(n183), .B(n178), .Y(n88) );
  NOR2X1 U139 ( .A(n190), .B(n177), .Y(n87) );
  NOR2X1 U140 ( .A(n189), .B(n177), .Y(n86) );
  NOR2X1 U141 ( .A(n188), .B(n177), .Y(n85) );
  NOR2X1 U142 ( .A(n187), .B(n177), .Y(n84) );
  NOR2X1 U143 ( .A(n186), .B(n177), .Y(n83) );
  NOR2X1 U144 ( .A(n185), .B(n177), .Y(n82) );
  NOR2X1 U145 ( .A(n184), .B(n177), .Y(n81) );
  NOR2X1 U146 ( .A(n183), .B(n177), .Y(n80) );
  NOR2X1 U147 ( .A(n190), .B(n176), .Y(n79) );
  NOR2X1 U148 ( .A(n189), .B(n176), .Y(n78) );
  NOR2X1 U149 ( .A(n188), .B(n176), .Y(n77) );
  NOR2X1 U150 ( .A(n187), .B(n176), .Y(n76) );
  NOR2X1 U151 ( .A(n186), .B(n176), .Y(n75) );
  NOR2X1 U152 ( .A(n185), .B(n176), .Y(n74) );
  NOR2X1 U153 ( .A(n184), .B(n176), .Y(n73) );
  NOR2X1 U154 ( .A(n183), .B(n176), .Y(n72) );
  NOR2X1 U155 ( .A(n182), .B(n189), .Y(n126) );
  NOR2X1 U156 ( .A(n182), .B(n188), .Y(n125) );
  NOR2X1 U157 ( .A(n182), .B(n187), .Y(n124) );
  NOR2X1 U158 ( .A(n182), .B(n186), .Y(n123) );
  NOR2X1 U159 ( .A(n182), .B(n185), .Y(n122) );
  NOR2X1 U160 ( .A(n182), .B(n184), .Y(n121) );
  NOR2X1 U161 ( .A(n182), .B(n183), .Y(n120) );
  NOR2X1 U162 ( .A(n190), .B(n181), .Y(n119) );
  NOR2X1 U163 ( .A(n189), .B(n181), .Y(n118) );
  NOR2X1 U164 ( .A(n188), .B(n181), .Y(n117) );
  NOR2X1 U165 ( .A(n187), .B(n181), .Y(n116) );
  NOR2X1 U166 ( .A(n186), .B(n181), .Y(n115) );
  NOR2X1 U167 ( .A(n185), .B(n181), .Y(n114) );
  NOR2X1 U168 ( .A(n184), .B(n181), .Y(n113) );
  NOR2X1 U169 ( .A(n183), .B(n181), .Y(n112) );
  NOR2X1 U170 ( .A(n190), .B(n180), .Y(n111) );
  NOR2X1 U171 ( .A(n189), .B(n180), .Y(n110) );
  NOR2X1 U172 ( .A(n188), .B(n180), .Y(n109) );
  NOR2X1 U173 ( .A(n187), .B(n180), .Y(n108) );
  NOR2X1 U174 ( .A(n186), .B(n180), .Y(n107) );
  NOR2X1 U175 ( .A(n185), .B(n180), .Y(n106) );
  NOR2X1 U176 ( .A(n184), .B(n180), .Y(n105) );
  NOR2X1 U177 ( .A(n183), .B(n180), .Y(n104) );
  NOR2X1 U178 ( .A(n190), .B(n179), .Y(n103) );
  NOR2X1 U179 ( .A(n179), .B(n189), .Y(n102) );
  NOR2X1 U180 ( .A(n179), .B(n188), .Y(n101) );
  NOR2X1 U181 ( .A(n179), .B(n187), .Y(n100) );
endmodule


module Equation_Implementation_DW_mult_uns_6 ( a, b, product );
  input [5:0] a;
  input [7:0] b;
  output [13:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166;

  ADDFX2 U2 ( .A(n13), .B(n60), .CI(n2), .CO(product[13]), .S(product[12]) );
  ADDFX2 U3 ( .A(n16), .B(n14), .CI(n3), .CO(n2), .S(product[11]) );
  ADDFX2 U4 ( .A(n19), .B(n17), .CI(n4), .CO(n3), .S(product[10]) );
  ADDFX2 U5 ( .A(n20), .B(n24), .CI(n5), .CO(n4), .S(product[9]) );
  ADDFX2 U6 ( .A(n25), .B(n31), .CI(n6), .CO(n5), .S(product[8]) );
  ADDFX2 U7 ( .A(n32), .B(n37), .CI(n7), .CO(n6), .S(product[7]) );
  ADDFX2 U8 ( .A(n38), .B(n43), .CI(n8), .CO(n7), .S(product[6]) );
  ADDFX2 U9 ( .A(n44), .B(n50), .CI(n9), .CO(n8), .S(product[5]) );
  ADDFX2 U10 ( .A(n51), .B(n54), .CI(n10), .CO(n9), .S(product[4]) );
  ADDFX2 U11 ( .A(n55), .B(n57), .CI(n11), .CO(n10), .S(product[3]) );
  ADDFX2 U12 ( .A(n12), .B(n91), .CI(n59), .CO(n11), .S(product[2]) );
  ADDHXL U13 ( .A(n99), .B(n106), .CO(n12), .S(product[1]) );
  ADDFX2 U14 ( .A(n61), .B(n68), .CI(n15), .CO(n13), .S(n14) );
  CMPR42X1 U15 ( .A(n62), .B(n76), .C(n21), .D(n69), .ICI(n18), .S(n17), .ICO(
        n15), .CO(n16) );
  CMPR42X1 U16 ( .A(n28), .B(n77), .C(n22), .D(n26), .ICI(n23), .S(n20), .ICO(
        n18), .CO(n19) );
  ADDFX2 U17 ( .A(n63), .B(n84), .CI(n70), .CO(n21), .S(n22) );
  CMPR42X1 U18 ( .A(n27), .B(n33), .C(n34), .D(n29), .ICI(n30), .S(n25), .ICO(
        n23), .CO(n24) );
  ADDFX2 U19 ( .A(n85), .B(n78), .CI(n92), .CO(n26), .S(n27) );
  ADDHXL U20 ( .A(n71), .B(n64), .CO(n28), .S(n29) );
  CMPR42X1 U21 ( .A(n39), .B(n93), .C(n35), .D(n40), .ICI(n36), .S(n32), .ICO(
        n30), .CO(n31) );
  CMPR42X1 U22 ( .A(n65), .B(n72), .C(n100), .D(n79), .ICI(n86), .S(n35), 
        .ICO(n33), .CO(n34) );
  CMPR42X1 U23 ( .A(n47), .B(n101), .C(n41), .D(n45), .ICI(n42), .S(n38), 
        .ICO(n36), .CO(n37) );
  CMPR42X1 U24 ( .A(n66), .B(n73), .C(n87), .D(n80), .ICI(n94), .S(n41), .ICO(
        n39), .CO(n40) );
  CMPR42X1 U25 ( .A(n52), .B(n95), .C(n48), .D(n46), .ICI(n49), .S(n44), .ICO(
        n42), .CO(n43) );
  ADDFX2 U26 ( .A(n81), .B(n102), .CI(n88), .CO(n45), .S(n46) );
  ADDHXL U27 ( .A(n74), .B(n67), .CO(n47), .S(n48) );
  CMPR42X1 U28 ( .A(n89), .B(n103), .C(n56), .D(n96), .ICI(n53), .S(n51), 
        .ICO(n49), .CO(n50) );
  ADDHXL U29 ( .A(n82), .B(n75), .CO(n52), .S(n53) );
  ADDFX2 U30 ( .A(n97), .B(n104), .CI(n58), .CO(n54), .S(n55) );
  ADDHXL U31 ( .A(n90), .B(n83), .CO(n56), .S(n57) );
  ADDHXL U32 ( .A(n105), .B(n98), .CO(n58), .S(n59) );
  CLKINVX2 U97 ( .A(a[0]), .Y(n158) );
  CLKINVX3 U98 ( .A(b[0]), .Y(n166) );
  CLKINVX3 U99 ( .A(b[1]), .Y(n165) );
  CLKINVX3 U100 ( .A(b[2]), .Y(n164) );
  CLKINVX3 U101 ( .A(b[3]), .Y(n163) );
  CLKINVX3 U102 ( .A(b[5]), .Y(n161) );
  CLKINVX3 U103 ( .A(b[4]), .Y(n162) );
  CLKINVX3 U104 ( .A(b[7]), .Y(n159) );
  CLKINVX3 U105 ( .A(b[6]), .Y(n160) );
  CLKINVX3 U106 ( .A(a[1]), .Y(n157) );
  CLKINVX3 U107 ( .A(a[3]), .Y(n155) );
  CLKINVX3 U108 ( .A(a[2]), .Y(n156) );
  CLKINVX3 U109 ( .A(a[5]), .Y(n153) );
  CLKINVX3 U110 ( .A(a[4]), .Y(n154) );
  NOR2X1 U111 ( .A(n158), .B(n166), .Y(product[0]) );
  NOR2X1 U112 ( .A(n166), .B(n157), .Y(n99) );
  NOR2X1 U113 ( .A(n157), .B(n165), .Y(n98) );
  NOR2X1 U114 ( .A(n157), .B(n164), .Y(n97) );
  NOR2X1 U115 ( .A(n157), .B(n163), .Y(n96) );
  NOR2X1 U116 ( .A(n157), .B(n162), .Y(n95) );
  NOR2X1 U117 ( .A(n157), .B(n161), .Y(n94) );
  NOR2X1 U118 ( .A(n157), .B(n160), .Y(n93) );
  NOR2X1 U119 ( .A(n157), .B(n159), .Y(n92) );
  NOR2X1 U120 ( .A(n166), .B(n156), .Y(n91) );
  NOR2X1 U121 ( .A(n165), .B(n156), .Y(n90) );
  NOR2X1 U122 ( .A(n164), .B(n156), .Y(n89) );
  NOR2X1 U123 ( .A(n163), .B(n156), .Y(n88) );
  NOR2X1 U124 ( .A(n162), .B(n156), .Y(n87) );
  NOR2X1 U125 ( .A(n161), .B(n156), .Y(n86) );
  NOR2X1 U126 ( .A(n160), .B(n156), .Y(n85) );
  NOR2X1 U127 ( .A(n159), .B(n156), .Y(n84) );
  NOR2X1 U128 ( .A(n166), .B(n155), .Y(n83) );
  NOR2X1 U129 ( .A(n165), .B(n155), .Y(n82) );
  NOR2X1 U130 ( .A(n164), .B(n155), .Y(n81) );
  NOR2X1 U131 ( .A(n163), .B(n155), .Y(n80) );
  NOR2X1 U132 ( .A(n162), .B(n155), .Y(n79) );
  NOR2X1 U133 ( .A(n161), .B(n155), .Y(n78) );
  NOR2X1 U134 ( .A(n160), .B(n155), .Y(n77) );
  NOR2X1 U135 ( .A(n159), .B(n155), .Y(n76) );
  NOR2X1 U136 ( .A(n166), .B(n154), .Y(n75) );
  NOR2X1 U137 ( .A(n165), .B(n154), .Y(n74) );
  NOR2X1 U138 ( .A(n164), .B(n154), .Y(n73) );
  NOR2X1 U139 ( .A(n163), .B(n154), .Y(n72) );
  NOR2X1 U140 ( .A(n162), .B(n154), .Y(n71) );
  NOR2X1 U141 ( .A(n161), .B(n154), .Y(n70) );
  NOR2X1 U142 ( .A(n160), .B(n154), .Y(n69) );
  NOR2X1 U143 ( .A(n159), .B(n154), .Y(n68) );
  NOR2X1 U144 ( .A(n166), .B(n153), .Y(n67) );
  NOR2X1 U145 ( .A(n165), .B(n153), .Y(n66) );
  NOR2X1 U146 ( .A(n164), .B(n153), .Y(n65) );
  NOR2X1 U147 ( .A(n163), .B(n153), .Y(n64) );
  NOR2X1 U148 ( .A(n162), .B(n153), .Y(n63) );
  NOR2X1 U149 ( .A(n161), .B(n153), .Y(n62) );
  NOR2X1 U150 ( .A(n160), .B(n153), .Y(n61) );
  NOR2X1 U151 ( .A(n159), .B(n153), .Y(n60) );
  NOR2X1 U152 ( .A(n158), .B(n165), .Y(n106) );
  NOR2X1 U153 ( .A(n158), .B(n164), .Y(n105) );
  NOR2X1 U154 ( .A(n158), .B(n163), .Y(n104) );
  NOR2X1 U155 ( .A(n158), .B(n162), .Y(n103) );
  NOR2X1 U156 ( .A(n158), .B(n161), .Y(n102) );
  NOR2X1 U157 ( .A(n158), .B(n160), .Y(n101) );
  NOR2X1 U158 ( .A(n158), .B(n159), .Y(n100) );
endmodule


module Equation_Implementation_DW01_add_144 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;

  wire   [15:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  XOR2X1 U1 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  AND2X2 U2 ( .A(A[14]), .B(carry[14]), .Y(SUM[15]) );
  AND2X1 U3 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module Equation_Implementation_DW01_add_151 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;
  assign SUM[0] = B[0];

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .Y(SUM[9]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X1 U1 ( .A(B[1]), .B(A[1]), .Y(carry[2]) );
  XOR2XL U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module Equation_Implementation_DW_mult_uns_12 ( a, b, product );
  input [31:0] a;
  input [9:0] b;
  output [41:0] product;
  wire   n19, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993;
  assign n19 = b[5];

  ADDFX2 U43 ( .A(n79), .B(n81), .CI(n43), .CO(n42), .S(product[30]) );
  ADDFX2 U44 ( .A(n82), .B(n84), .CI(n44), .CO(n43), .S(product[29]) );
  ADDFX2 U45 ( .A(n85), .B(n87), .CI(n45), .CO(n44), .S(product[28]) );
  ADDFX2 U46 ( .A(n88), .B(n90), .CI(n46), .CO(n45), .S(product[27]) );
  ADDFX2 U47 ( .A(n91), .B(n93), .CI(n47), .CO(n46), .S(product[26]) );
  ADDFX2 U48 ( .A(n94), .B(n96), .CI(n48), .CO(n47), .S(product[25]) );
  ADDFX2 U49 ( .A(n97), .B(n99), .CI(n49), .CO(n48), .S(product[24]) );
  ADDFX2 U50 ( .A(n100), .B(n102), .CI(n50), .CO(n49), .S(product[23]) );
  ADDFX2 U51 ( .A(n103), .B(n105), .CI(n51), .CO(n50), .S(product[22]) );
  ADDFX2 U52 ( .A(n106), .B(n108), .CI(n52), .CO(n51), .S(product[21]) );
  ADDFX2 U53 ( .A(n109), .B(n111), .CI(n53), .CO(n52), .S(product[20]) );
  ADDFX2 U54 ( .A(n112), .B(n114), .CI(n54), .CO(n53), .S(product[19]) );
  ADDFX2 U55 ( .A(n115), .B(n117), .CI(n55), .CO(n54), .S(product[18]) );
  ADDFX2 U56 ( .A(n118), .B(n120), .CI(n56), .CO(n55), .S(product[17]) );
  ADDFX2 U57 ( .A(n121), .B(n123), .CI(n57), .CO(n56), .S(product[16]) );
  ADDFX2 U58 ( .A(n124), .B(n126), .CI(n58), .CO(n57), .S(product[15]) );
  ADDFX2 U59 ( .A(n127), .B(n129), .CI(n59), .CO(n58), .S(product[14]) );
  ADDFX2 U60 ( .A(n130), .B(n132), .CI(n60), .CO(n59), .S(product[13]) );
  ADDFX2 U61 ( .A(n133), .B(n135), .CI(n61), .CO(n60), .S(product[12]) );
  ADDFX2 U62 ( .A(n136), .B(n138), .CI(n62), .CO(n61), .S(product[11]) );
  ADDFX2 U63 ( .A(n139), .B(n141), .CI(n63), .CO(n62), .S(product[10]) );
  ADDFX2 U64 ( .A(n142), .B(n143), .CI(n64), .CO(n63), .S(product[9]) );
  ADDFX2 U65 ( .A(n144), .B(n147), .CI(n65), .CO(n64), .S(product[8]) );
  ADDFX2 U66 ( .A(n148), .B(n151), .CI(n66), .CO(n65), .S(product[7]) );
  ADDFX2 U67 ( .A(n152), .B(n155), .CI(n67), .CO(n66), .S(product[6]) );
  ADDFX2 U68 ( .A(n156), .B(n157), .CI(n68), .CO(n67), .S(product[5]) );
  ADDFX2 U69 ( .A(n158), .B(n327), .CI(n69), .CO(n68), .S(product[4]) );
  ADDFX2 U70 ( .A(n160), .B(n357), .CI(n70), .CO(n69), .S(product[3]) );
  ADDHXL U71 ( .A(n358), .B(n71), .CO(n70), .S(product[2]) );
  ADDHXL U72 ( .A(n72), .B(n359), .CO(n71), .S(product[1]) );
  CMPR42X1 U78 ( .A(n275), .B(a[20]), .C(n330), .D(n301), .ICI(n80), .S(n79), 
        .ICO(n77), .CO(n78) );
  CMPR42X1 U79 ( .A(n276), .B(a[19]), .C(n331), .D(n302), .ICI(n83), .S(n82), 
        .ICO(n80), .CO(n81) );
  CMPR42X1 U80 ( .A(n277), .B(a[18]), .C(n332), .D(n303), .ICI(n86), .S(n85), 
        .ICO(n83), .CO(n84) );
  CMPR42X1 U81 ( .A(n278), .B(a[17]), .C(n333), .D(n304), .ICI(n89), .S(n88), 
        .ICO(n86), .CO(n87) );
  CMPR42X1 U82 ( .A(n279), .B(a[16]), .C(n334), .D(n305), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U83 ( .A(n280), .B(a[15]), .C(n335), .D(n306), .ICI(n95), .S(n94), 
        .ICO(n92), .CO(n93) );
  CMPR42X1 U84 ( .A(n281), .B(a[14]), .C(n336), .D(n307), .ICI(n98), .S(n97), 
        .ICO(n95), .CO(n96) );
  CMPR42X1 U85 ( .A(n282), .B(a[13]), .C(n337), .D(n308), .ICI(n101), .S(n100), 
        .ICO(n98), .CO(n99) );
  CMPR42X1 U86 ( .A(n283), .B(a[12]), .C(n338), .D(n309), .ICI(n104), .S(n103), 
        .ICO(n101), .CO(n102) );
  CMPR42X1 U87 ( .A(n284), .B(a[11]), .C(n107), .D(n310), .ICI(n339), .S(n106), 
        .ICO(n104), .CO(n105) );
  CMPR42X1 U88 ( .A(n285), .B(a[10]), .C(n110), .D(n311), .ICI(n340), .S(n109), 
        .ICO(n107), .CO(n108) );
  CMPR42X1 U89 ( .A(n286), .B(a[9]), .C(n113), .D(n312), .ICI(n341), .S(n112), 
        .ICO(n110), .CO(n111) );
  CMPR42X1 U90 ( .A(n287), .B(a[8]), .C(n116), .D(n313), .ICI(n342), .S(n115), 
        .ICO(n113), .CO(n114) );
  CMPR42X1 U91 ( .A(n288), .B(a[7]), .C(n119), .D(n314), .ICI(n343), .S(n118), 
        .ICO(n116), .CO(n117) );
  CMPR42X1 U92 ( .A(n289), .B(a[6]), .C(n122), .D(n315), .ICI(n344), .S(n121), 
        .ICO(n119), .CO(n120) );
  CMPR42X1 U93 ( .A(n290), .B(a[5]), .C(n125), .D(n316), .ICI(n345), .S(n124), 
        .ICO(n122), .CO(n123) );
  CMPR42X1 U94 ( .A(n291), .B(a[4]), .C(n128), .D(n317), .ICI(n346), .S(n127), 
        .ICO(n125), .CO(n126) );
  CMPR42X1 U95 ( .A(n292), .B(a[3]), .C(n131), .D(n318), .ICI(n347), .S(n130), 
        .ICO(n128), .CO(n129) );
  CMPR42X1 U96 ( .A(n293), .B(a[2]), .C(n134), .D(n319), .ICI(n348), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U97 ( .A(n294), .B(a[1]), .C(n137), .D(n320), .ICI(n349), .S(n136), 
        .ICO(n134), .CO(n135) );
  CMPR42X1 U98 ( .A(n295), .B(a[0]), .C(n140), .D(n321), .ICI(n350), .S(n139), 
        .ICO(n137), .CO(n138) );
  ADDFX2 U100 ( .A(n146), .B(n149), .CI(n352), .CO(n143), .S(n144) );
  ADDFX2 U102 ( .A(n150), .B(n298), .CI(n353), .CO(n147), .S(n148) );
  ADDHXL U103 ( .A(n324), .B(n153), .CO(n149), .S(n150) );
  ADDFX2 U104 ( .A(n154), .B(n325), .CI(n354), .CO(n151), .S(n152) );
  ADDHXL U106 ( .A(n326), .B(n355), .CO(n155), .S(n156) );
  ADDHXL U107 ( .A(n356), .B(n159), .CO(n157), .S(n158) );
  ADDHXL U108 ( .A(n19), .B(n328), .CO(n159), .S(n160) );
  ADDFX2 U509 ( .A(a[29]), .B(a[30]), .CI(n213), .CO(n212), .S(n243) );
  ADDFX2 U510 ( .A(a[28]), .B(a[29]), .CI(n214), .CO(n213), .S(n244) );
  ADDFX2 U511 ( .A(a[27]), .B(a[28]), .CI(n215), .CO(n214), .S(n245) );
  ADDFX2 U512 ( .A(a[26]), .B(a[27]), .CI(n216), .CO(n215), .S(n246) );
  ADDFX2 U513 ( .A(a[25]), .B(a[26]), .CI(n217), .CO(n216), .S(n247) );
  ADDFX2 U514 ( .A(a[24]), .B(a[25]), .CI(n218), .CO(n217), .S(n248) );
  ADDFX2 U515 ( .A(a[23]), .B(a[24]), .CI(n219), .CO(n218), .S(n249) );
  ADDFX2 U516 ( .A(a[22]), .B(a[23]), .CI(n220), .CO(n219), .S(n250) );
  ADDFX2 U517 ( .A(a[21]), .B(a[22]), .CI(n221), .CO(n220), .S(n251) );
  ADDFX2 U518 ( .A(a[20]), .B(a[21]), .CI(n222), .CO(n221), .S(n252) );
  ADDFX2 U519 ( .A(a[19]), .B(a[20]), .CI(n223), .CO(n222), .S(n253) );
  ADDFX2 U520 ( .A(a[18]), .B(a[19]), .CI(n224), .CO(n223), .S(n254) );
  ADDFX2 U521 ( .A(a[17]), .B(a[18]), .CI(n225), .CO(n224), .S(n255) );
  ADDFX2 U522 ( .A(a[16]), .B(a[17]), .CI(n226), .CO(n225), .S(n256) );
  ADDFX2 U523 ( .A(a[15]), .B(a[16]), .CI(n227), .CO(n226), .S(n257) );
  ADDFX2 U524 ( .A(a[14]), .B(a[15]), .CI(n228), .CO(n227), .S(n258) );
  ADDFX2 U525 ( .A(a[13]), .B(a[14]), .CI(n229), .CO(n228), .S(n259) );
  ADDFX2 U526 ( .A(a[12]), .B(a[13]), .CI(n230), .CO(n229), .S(n260) );
  ADDFX2 U527 ( .A(a[11]), .B(a[12]), .CI(n231), .CO(n230), .S(n261) );
  ADDFX2 U528 ( .A(a[10]), .B(a[11]), .CI(n232), .CO(n231), .S(n262) );
  ADDFX2 U529 ( .A(a[9]), .B(a[10]), .CI(n233), .CO(n232), .S(n263) );
  ADDFX2 U530 ( .A(a[8]), .B(a[9]), .CI(n234), .CO(n233), .S(n264) );
  ADDFX2 U531 ( .A(a[7]), .B(a[8]), .CI(n235), .CO(n234), .S(n265) );
  ADDFX2 U532 ( .A(a[6]), .B(a[7]), .CI(n236), .CO(n235), .S(n266) );
  ADDFX2 U533 ( .A(a[5]), .B(a[6]), .CI(n237), .CO(n236), .S(n267) );
  ADDFX2 U534 ( .A(a[4]), .B(a[5]), .CI(n238), .CO(n237), .S(n268) );
  ADDFX2 U535 ( .A(a[3]), .B(a[4]), .CI(n239), .CO(n238), .S(n269) );
  ADDFX2 U536 ( .A(a[2]), .B(a[3]), .CI(n240), .CO(n239), .S(n270) );
  ADDFX2 U537 ( .A(a[1]), .B(a[2]), .CI(n241), .CO(n240), .S(n271) );
  OR2X2 U541 ( .A(n19), .B(n943), .Y(n699) );
  OR2X2 U542 ( .A(n993), .B(n991), .Y(n700) );
  CMPR22X1 U543 ( .A(a[1]), .B(n707), .CO(n241), .S(n272) );
  CMPR22X1 U544 ( .A(n297), .B(n323), .CO(n145), .S(n146) );
  AOI222XL U545 ( .A0(n272), .A1(n802), .B0(a[1]), .B1(n738), .C0(a[0]), .C1(
        n720), .Y(n298) );
  XNOR2XL U546 ( .A(n889), .B(n19), .Y(n327) );
  AOI222XL U547 ( .A0(n709), .A1(n707), .B0(n733), .B1(a[1]), .C0(n732), .C1(
        n272), .Y(n889) );
  AOI222XL U548 ( .A0(n272), .A1(n704), .B0(a[1]), .B1(n717), .C0(n708), .C1(
        n714), .Y(n826) );
  INVX1 U549 ( .A(b[7]), .Y(n993) );
  XOR3X2 U550 ( .A(a[30]), .B(a[31]), .C(n212), .Y(n242) );
  BUFX4 U551 ( .A(n824), .Y(n705) );
  CLKINVX3 U552 ( .A(n732), .Y(n731) );
  CLKINVX3 U553 ( .A(n719), .Y(n718) );
  CLKINVX3 U554 ( .A(n985), .Y(n720) );
  CLKINVX3 U555 ( .A(n700), .Y(n738) );
  CLKINVX3 U556 ( .A(n713), .Y(n712) );
  CLKINVX3 U557 ( .A(n719), .Y(n717) );
  INVX1 U558 ( .A(n805), .Y(n719) );
  CLKINVX3 U559 ( .A(n700), .Y(n739) );
  CLKINVX3 U560 ( .A(n699), .Y(n733) );
  BUFX3 U561 ( .A(n806), .Y(n702) );
  CLKINVX3 U562 ( .A(n699), .Y(n734) );
  CLKINVX3 U563 ( .A(n716), .Y(n715) );
  INVX1 U564 ( .A(n729), .Y(n732) );
  BUFX3 U565 ( .A(n806), .Y(n703) );
  CLKINVX3 U566 ( .A(n985), .Y(n721) );
  INVX1 U567 ( .A(n944), .Y(n297) );
  INVX1 U568 ( .A(n948), .Y(n295) );
  INVX1 U569 ( .A(n950), .Y(n294) );
  INVX1 U570 ( .A(n952), .Y(n293) );
  INVX1 U571 ( .A(n954), .Y(n292) );
  INVX1 U572 ( .A(n956), .Y(n291) );
  INVX1 U573 ( .A(n958), .Y(n290) );
  INVX1 U574 ( .A(n960), .Y(n289) );
  INVX1 U575 ( .A(n962), .Y(n288) );
  INVX1 U576 ( .A(n964), .Y(n287) );
  INVX1 U577 ( .A(n966), .Y(n286) );
  INVX1 U578 ( .A(n968), .Y(n285) );
  INVX1 U579 ( .A(n970), .Y(n284) );
  XOR2X1 U580 ( .A(n740), .B(n741), .Y(n142) );
  XOR2XL U581 ( .A(n296), .B(n145), .Y(n740) );
  XOR2X1 U582 ( .A(n322), .B(n351), .Y(n741) );
  NAND3BX1 U583 ( .AN(n746), .B(n747), .C(n748), .Y(n141) );
  AND2X2 U584 ( .A(n351), .B(n322), .Y(n746) );
  MXI2XL U585 ( .A(n742), .B(n743), .S0(n145), .Y(n747) );
  INVX1 U586 ( .A(n268), .Y(n794) );
  INVX1 U587 ( .A(n264), .Y(n786) );
  AND2X1 U588 ( .A(n145), .B(n296), .Y(n140) );
  MXI2XL U589 ( .A(n744), .B(n745), .S0(n145), .Y(n748) );
  AND2X2 U590 ( .A(n351), .B(n296), .Y(n744) );
  NOR2BX1 U591 ( .AN(n351), .B(n296), .Y(n745) );
  INVX1 U592 ( .A(n269), .Y(n796) );
  INVX1 U593 ( .A(n153), .Y(n154) );
  INVX1 U594 ( .A(n267), .Y(n792) );
  INVX1 U595 ( .A(n266), .Y(n790) );
  INVX1 U596 ( .A(n265), .Y(n788) );
  INVX1 U597 ( .A(n263), .Y(n784) );
  INVX1 U598 ( .A(n262), .Y(n782) );
  INVX1 U599 ( .A(n261), .Y(n780) );
  INVX1 U600 ( .A(n260), .Y(n778) );
  INVX1 U601 ( .A(n259), .Y(n776) );
  INVX1 U602 ( .A(n258), .Y(n774) );
  INVX1 U603 ( .A(n257), .Y(n772) );
  INVX1 U604 ( .A(n256), .Y(n770) );
  INVX1 U605 ( .A(n255), .Y(n768) );
  INVX1 U606 ( .A(n254), .Y(n766) );
  INVX1 U607 ( .A(n253), .Y(n764) );
  INVX1 U608 ( .A(n252), .Y(n762) );
  INVX1 U609 ( .A(n270), .Y(n798) );
  NOR2BX1 U610 ( .AN(n322), .B(n296), .Y(n743) );
  INVX1 U611 ( .A(n271), .Y(n800) );
  AND2X2 U612 ( .A(n322), .B(n296), .Y(n742) );
  INVX1 U613 ( .A(n871), .Y(n805) );
  CLKINVX3 U614 ( .A(n716), .Y(n714) );
  INVX1 U615 ( .A(n804), .Y(n716) );
  CLKINVX3 U616 ( .A(n713), .Y(n711) );
  INVX1 U617 ( .A(n803), .Y(n713) );
  CLKINVX3 U618 ( .A(n737), .Y(n735) );
  INVX1 U619 ( .A(n705), .Y(n802) );
  CLKINVX3 U620 ( .A(n931), .Y(n709) );
  INVX1 U621 ( .A(n704), .Y(n806) );
  CLKINVX3 U622 ( .A(b[7]), .Y(n723) );
  INVX1 U623 ( .A(n730), .Y(n729) );
  CLKINVX3 U624 ( .A(n19), .Y(n725) );
  CLKINVX3 U625 ( .A(n931), .Y(n710) );
  CLKINVX3 U626 ( .A(n737), .Y(n736) );
  CLKINVX3 U627 ( .A(n728), .Y(n727) );
  CLKINVX3 U628 ( .A(n19), .Y(n724) );
  INVX1 U629 ( .A(n972), .Y(n283) );
  INVX1 U630 ( .A(n974), .Y(n282) );
  INVX1 U631 ( .A(n246), .Y(n753) );
  CLKINVX3 U632 ( .A(n946), .Y(n296) );
  INVX1 U633 ( .A(a[1]), .Y(n801) );
  INVX1 U634 ( .A(a[2]), .Y(n799) );
  INVX1 U635 ( .A(a[3]), .Y(n797) );
  INVX1 U636 ( .A(a[4]), .Y(n795) );
  INVX1 U637 ( .A(a[5]), .Y(n793) );
  INVX1 U638 ( .A(a[6]), .Y(n791) );
  INVX1 U639 ( .A(a[7]), .Y(n789) );
  INVX1 U640 ( .A(a[8]), .Y(n787) );
  INVX1 U641 ( .A(a[9]), .Y(n785) );
  INVX1 U642 ( .A(a[10]), .Y(n783) );
  INVX1 U643 ( .A(a[11]), .Y(n781) );
  INVX1 U644 ( .A(a[12]), .Y(n779) );
  INVX1 U645 ( .A(a[13]), .Y(n777) );
  INVX1 U646 ( .A(a[14]), .Y(n775) );
  INVX1 U647 ( .A(a[15]), .Y(n773) );
  INVX1 U648 ( .A(a[16]), .Y(n771) );
  INVX1 U649 ( .A(a[17]), .Y(n769) );
  INVX1 U650 ( .A(a[18]), .Y(n767) );
  INVX1 U651 ( .A(a[19]), .Y(n765) );
  INVX1 U652 ( .A(a[20]), .Y(n763) );
  CLKINVX3 U653 ( .A(a[21]), .Y(n761) );
  INVX1 U654 ( .A(n817), .Y(n803) );
  INVX1 U655 ( .A(n868), .Y(n804) );
  NAND2BXL U656 ( .AN(n991), .B(n993), .Y(n824) );
  INVX1 U657 ( .A(n823), .Y(n737) );
  BUFX3 U658 ( .A(n818), .Y(n704) );
  NOR2BX1 U659 ( .AN(b[0]), .B(n887), .Y(n818) );
  CLKINVX3 U660 ( .A(n728), .Y(n726) );
  INVX1 U661 ( .A(n819), .Y(n728) );
  INVX1 U662 ( .A(n820), .Y(n730) );
  CLKINVX3 U663 ( .A(b[7]), .Y(n722) );
  INVX1 U664 ( .A(n706), .Y(n707) );
  INVX1 U665 ( .A(a[30]), .Y(n749) );
  INVX1 U666 ( .A(n976), .Y(n281) );
  INVX1 U667 ( .A(n978), .Y(n280) );
  INVX1 U668 ( .A(n982), .Y(n278) );
  INVX1 U669 ( .A(n980), .Y(n279) );
  INVX1 U670 ( .A(n984), .Y(n277) );
  INVX1 U671 ( .A(n987), .Y(n276) );
  INVX1 U672 ( .A(n989), .Y(n275) );
  XOR2X1 U673 ( .A(n77), .B(n701), .Y(n810) );
  XOR2X1 U674 ( .A(n724), .B(b[2]), .Y(n701) );
  INVX1 U675 ( .A(n249), .Y(n758) );
  XOR2X1 U676 ( .A(n822), .B(n761), .Y(n811) );
  INVX1 U677 ( .A(n245), .Y(n751) );
  INVX1 U678 ( .A(n706), .Y(n708) );
  INVX1 U679 ( .A(a[22]), .Y(n760) );
  INVX1 U680 ( .A(a[24]), .Y(n757) );
  INVX1 U681 ( .A(a[26]), .Y(n754) );
  INVX1 U682 ( .A(a[27]), .Y(n752) );
  INVX1 U683 ( .A(a[29]), .Y(n750) );
  INVX1 U684 ( .A(a[0]), .Y(n706) );
  INVX1 U685 ( .A(n248), .Y(n756) );
  CLKINVX3 U686 ( .A(a[23]), .Y(n759) );
  INVX1 U687 ( .A(a[25]), .Y(n755) );
  XOR2X1 U688 ( .A(n807), .B(n808), .Y(product[31]) );
  XNOR2X1 U689 ( .A(n78), .B(n42), .Y(n808) );
  XOR2X1 U690 ( .A(n809), .B(n810), .Y(n807) );
  XOR2X1 U691 ( .A(n811), .B(n812), .Y(n809) );
  XOR2X1 U692 ( .A(n813), .B(n814), .Y(n812) );
  NAND2X1 U693 ( .A(n815), .B(n816), .Y(n814) );
  AOI22X1 U694 ( .A0(a[31]), .A1(n718), .B0(a[30]), .B1(n715), .Y(n816) );
  AOI22X1 U695 ( .A0(a[29]), .A1(n817), .B0(n242), .B1(n704), .Y(n815) );
  OAI221XL U696 ( .A0(n727), .A1(n754), .B0(n731), .B1(n751), .C0(n821), .Y(
        n813) );
  AOI22X1 U697 ( .A0(a[28]), .A1(n734), .B0(a[27]), .B1(n710), .Y(n821) );
  OAI221XL U698 ( .A0(n735), .A1(n759), .B0(n705), .B1(n756), .C0(n825), .Y(
        n822) );
  AOI22X1 U699 ( .A0(a[25]), .A1(n739), .B0(a[24]), .B1(n721), .Y(n825) );
  AOI221X1 U700 ( .A0(n708), .A1(n717), .B0(n708), .B1(n704), .C0(n723), .Y(
        n72) );
  XNOR2X1 U701 ( .A(b[2]), .B(n826), .Y(n359) );
  XNOR2X1 U702 ( .A(n827), .B(n722), .Y(n358) );
  OAI221XL U703 ( .A0(n712), .A1(n706), .B0(n702), .B1(n800), .C0(n828), .Y(
        n827) );
  AOI22X1 U704 ( .A0(a[2]), .A1(n717), .B0(a[1]), .B1(n714), .Y(n828) );
  XNOR2X1 U705 ( .A(n829), .B(n722), .Y(n357) );
  OAI221XL U706 ( .A0(n711), .A1(n801), .B0(n702), .B1(n798), .C0(n830), .Y(
        n829) );
  AOI22X1 U707 ( .A0(a[3]), .A1(n717), .B0(a[2]), .B1(n714), .Y(n830) );
  XNOR2X1 U708 ( .A(n831), .B(n722), .Y(n356) );
  OAI221XL U709 ( .A0(n711), .A1(n799), .B0(n702), .B1(n796), .C0(n832), .Y(
        n831) );
  AOI22X1 U710 ( .A0(a[4]), .A1(n717), .B0(a[3]), .B1(n714), .Y(n832) );
  XNOR2X1 U711 ( .A(n833), .B(n722), .Y(n355) );
  OAI221XL U712 ( .A0(n711), .A1(n797), .B0(n702), .B1(n794), .C0(n834), .Y(
        n833) );
  AOI22X1 U713 ( .A0(a[5]), .A1(n717), .B0(a[4]), .B1(n714), .Y(n834) );
  XNOR2X1 U714 ( .A(n835), .B(n722), .Y(n354) );
  OAI221XL U715 ( .A0(n711), .A1(n795), .B0(n702), .B1(n792), .C0(n836), .Y(
        n835) );
  AOI22X1 U716 ( .A0(a[6]), .A1(n717), .B0(a[5]), .B1(n714), .Y(n836) );
  XNOR2X1 U717 ( .A(n837), .B(n722), .Y(n353) );
  OAI221XL U718 ( .A0(n711), .A1(n793), .B0(n702), .B1(n790), .C0(n838), .Y(
        n837) );
  AOI22X1 U719 ( .A0(a[7]), .A1(n717), .B0(a[6]), .B1(n714), .Y(n838) );
  XNOR2X1 U720 ( .A(n839), .B(n722), .Y(n352) );
  OAI221XL U721 ( .A0(n711), .A1(n791), .B0(n702), .B1(n788), .C0(n840), .Y(
        n839) );
  AOI22X1 U722 ( .A0(a[8]), .A1(n717), .B0(a[7]), .B1(n714), .Y(n840) );
  XNOR2X1 U723 ( .A(n841), .B(n722), .Y(n351) );
  OAI221XL U724 ( .A0(n711), .A1(n789), .B0(n702), .B1(n786), .C0(n842), .Y(
        n841) );
  AOI22X1 U725 ( .A0(a[9]), .A1(n717), .B0(a[8]), .B1(n714), .Y(n842) );
  XNOR2X1 U726 ( .A(n843), .B(n722), .Y(n350) );
  OAI221XL U727 ( .A0(n711), .A1(n787), .B0(n702), .B1(n784), .C0(n844), .Y(
        n843) );
  AOI22X1 U728 ( .A0(a[10]), .A1(n717), .B0(a[9]), .B1(n715), .Y(n844) );
  XNOR2X1 U729 ( .A(n845), .B(n722), .Y(n349) );
  OAI221XL U730 ( .A0(n711), .A1(n785), .B0(n702), .B1(n782), .C0(n846), .Y(
        n845) );
  AOI22X1 U731 ( .A0(a[11]), .A1(n717), .B0(a[10]), .B1(n715), .Y(n846) );
  XNOR2X1 U732 ( .A(n847), .B(n722), .Y(n348) );
  OAI221XL U733 ( .A0(n711), .A1(n783), .B0(n702), .B1(n780), .C0(n848), .Y(
        n847) );
  AOI22X1 U734 ( .A0(a[12]), .A1(n717), .B0(a[11]), .B1(n715), .Y(n848) );
  XNOR2X1 U735 ( .A(n849), .B(n722), .Y(n347) );
  OAI221XL U736 ( .A0(n711), .A1(n781), .B0(n703), .B1(n778), .C0(n850), .Y(
        n849) );
  AOI22X1 U737 ( .A0(a[13]), .A1(n718), .B0(a[12]), .B1(n715), .Y(n850) );
  XNOR2X1 U738 ( .A(n851), .B(n722), .Y(n346) );
  OAI221XL U739 ( .A0(n711), .A1(n779), .B0(n703), .B1(n776), .C0(n852), .Y(
        n851) );
  AOI22X1 U740 ( .A0(a[14]), .A1(n718), .B0(a[13]), .B1(n715), .Y(n852) );
  XNOR2X1 U741 ( .A(n853), .B(n722), .Y(n345) );
  OAI221XL U742 ( .A0(n712), .A1(n777), .B0(n703), .B1(n774), .C0(n854), .Y(
        n853) );
  AOI22X1 U743 ( .A0(a[15]), .A1(n718), .B0(a[14]), .B1(n715), .Y(n854) );
  XNOR2X1 U744 ( .A(n855), .B(n722), .Y(n344) );
  OAI221XL U745 ( .A0(n712), .A1(n775), .B0(n703), .B1(n772), .C0(n856), .Y(
        n855) );
  AOI22X1 U746 ( .A0(a[16]), .A1(n718), .B0(a[15]), .B1(n715), .Y(n856) );
  XNOR2X1 U747 ( .A(n857), .B(n722), .Y(n343) );
  OAI221XL U748 ( .A0(n712), .A1(n773), .B0(n703), .B1(n770), .C0(n858), .Y(
        n857) );
  AOI22X1 U749 ( .A0(a[17]), .A1(n718), .B0(a[16]), .B1(n715), .Y(n858) );
  XNOR2X1 U750 ( .A(n859), .B(n993), .Y(n342) );
  OAI221XL U751 ( .A0(n712), .A1(n771), .B0(n703), .B1(n768), .C0(n860), .Y(
        n859) );
  AOI22X1 U752 ( .A0(a[18]), .A1(n718), .B0(a[17]), .B1(n715), .Y(n860) );
  XNOR2X1 U753 ( .A(n861), .B(n993), .Y(n341) );
  OAI221XL U754 ( .A0(n712), .A1(n769), .B0(n703), .B1(n766), .C0(n862), .Y(
        n861) );
  AOI22X1 U755 ( .A0(a[19]), .A1(n718), .B0(a[18]), .B1(n715), .Y(n862) );
  XNOR2X1 U756 ( .A(n863), .B(n723), .Y(n340) );
  OAI221XL U757 ( .A0(n712), .A1(n767), .B0(n703), .B1(n764), .C0(n864), .Y(
        n863) );
  AOI22X1 U758 ( .A0(a[20]), .A1(n718), .B0(a[19]), .B1(n715), .Y(n864) );
  XNOR2X1 U759 ( .A(n865), .B(n723), .Y(n339) );
  OAI221XL U760 ( .A0(n712), .A1(n765), .B0(n703), .B1(n762), .C0(n866), .Y(
        n865) );
  AOI22X1 U761 ( .A0(a[20]), .A1(n714), .B0(n718), .B1(a[21]), .Y(n866) );
  XNOR2X1 U762 ( .A(n867), .B(n723), .Y(n338) );
  OAI221XL U763 ( .A0(n712), .A1(n763), .B0(n761), .B1(n868), .C0(n869), .Y(
        n867) );
  AOI22X1 U764 ( .A0(n718), .A1(a[22]), .B0(n251), .B1(n704), .Y(n869) );
  XNOR2X1 U765 ( .A(n870), .B(n723), .Y(n337) );
  OAI221XL U766 ( .A0(n761), .A1(n712), .B0(n759), .B1(n871), .C0(n872), .Y(
        n870) );
  AOI22X1 U767 ( .A0(n714), .A1(a[22]), .B0(n250), .B1(n704), .Y(n872) );
  XNOR2X1 U768 ( .A(n873), .B(n723), .Y(n336) );
  OAI221XL U769 ( .A0(n760), .A1(n712), .B0(n703), .B1(n758), .C0(n874), .Y(
        n873) );
  AOI22X1 U770 ( .A0(n718), .A1(a[24]), .B0(n715), .B1(a[23]), .Y(n874) );
  XNOR2X1 U771 ( .A(n875), .B(n723), .Y(n335) );
  OAI221XL U772 ( .A0(n757), .A1(n868), .B0(n759), .B1(n711), .C0(n876), .Y(
        n875) );
  AOI22X1 U773 ( .A0(n718), .A1(a[25]), .B0(n704), .B1(n248), .Y(n876) );
  XNOR2X1 U774 ( .A(n877), .B(n723), .Y(n334) );
  OAI221XL U775 ( .A0(n757), .A1(n712), .B0(n754), .B1(n871), .C0(n878), .Y(
        n877) );
  AOI22X1 U776 ( .A0(n714), .A1(a[25]), .B0(n247), .B1(n704), .Y(n878) );
  XNOR2X1 U777 ( .A(n879), .B(n723), .Y(n333) );
  OAI221XL U778 ( .A0(n755), .A1(n712), .B0(n703), .B1(n753), .C0(n880), .Y(
        n879) );
  AOI22X1 U779 ( .A0(n718), .A1(a[27]), .B0(n715), .B1(a[26]), .Y(n880) );
  XNOR2X1 U780 ( .A(n881), .B(n723), .Y(n332) );
  OAI221XL U781 ( .A0(n752), .A1(n868), .B0(n754), .B1(n712), .C0(n882), .Y(
        n881) );
  AOI22X1 U782 ( .A0(n718), .A1(a[28]), .B0(n704), .B1(n245), .Y(n882) );
  XNOR2X1 U783 ( .A(n883), .B(n723), .Y(n331) );
  OAI221XL U784 ( .A0(n752), .A1(n711), .B0(n871), .B1(n750), .C0(n884), .Y(
        n883) );
  AOI22X1 U785 ( .A0(n714), .A1(a[28]), .B0(n244), .B1(n704), .Y(n884) );
  XNOR2X1 U786 ( .A(n885), .B(n723), .Y(n330) );
  OAI221XL U787 ( .A0(n871), .A1(n749), .B0(n868), .B1(n750), .C0(n886), .Y(
        n885) );
  AOI22X1 U788 ( .A0(n817), .A1(a[28]), .B0(n243), .B1(n704), .Y(n886) );
  NOR3X1 U789 ( .A(b[6]), .B(b[1]), .C(n887), .Y(n817) );
  NAND2BX1 U790 ( .AN(b[0]), .B(b[1]), .Y(n868) );
  NAND2X1 U791 ( .A(b[6]), .B(n887), .Y(n871) );
  XOR2X1 U792 ( .A(b[1]), .B(n723), .Y(n887) );
  XNOR2X1 U793 ( .A(n19), .B(n888), .Y(n328) );
  AOI22X1 U794 ( .A0(n708), .A1(n730), .B0(n708), .B1(n734), .Y(n888) );
  XNOR2X1 U795 ( .A(n890), .B(n724), .Y(n326) );
  OAI221XL U796 ( .A0(n726), .A1(n706), .B0(n731), .B1(n800), .C0(n891), .Y(
        n890) );
  AOI22X1 U797 ( .A0(a[2]), .A1(n733), .B0(a[1]), .B1(n709), .Y(n891) );
  XNOR2X1 U798 ( .A(n892), .B(n724), .Y(n325) );
  OAI221XL U799 ( .A0(n726), .A1(n801), .B0(n731), .B1(n798), .C0(n893), .Y(
        n892) );
  AOI22X1 U800 ( .A0(a[3]), .A1(n733), .B0(a[2]), .B1(n709), .Y(n893) );
  XNOR2X1 U801 ( .A(n894), .B(n725), .Y(n324) );
  OAI221XL U802 ( .A0(n726), .A1(n799), .B0(n731), .B1(n796), .C0(n895), .Y(
        n894) );
  AOI22X1 U803 ( .A0(a[4]), .A1(n733), .B0(a[3]), .B1(n709), .Y(n895) );
  XNOR2X1 U804 ( .A(n896), .B(n725), .Y(n323) );
  OAI221XL U805 ( .A0(n726), .A1(n797), .B0(n731), .B1(n794), .C0(n897), .Y(
        n896) );
  AOI22X1 U806 ( .A0(a[5]), .A1(n733), .B0(a[4]), .B1(n709), .Y(n897) );
  XNOR2X1 U807 ( .A(n898), .B(n725), .Y(n322) );
  OAI221XL U808 ( .A0(n726), .A1(n795), .B0(n731), .B1(n792), .C0(n899), .Y(
        n898) );
  AOI22X1 U809 ( .A0(a[6]), .A1(n733), .B0(a[5]), .B1(n709), .Y(n899) );
  XNOR2X1 U810 ( .A(n900), .B(n725), .Y(n321) );
  OAI221XL U811 ( .A0(n726), .A1(n793), .B0(n731), .B1(n790), .C0(n901), .Y(
        n900) );
  AOI22X1 U812 ( .A0(a[7]), .A1(n733), .B0(a[6]), .B1(n709), .Y(n901) );
  XNOR2X1 U813 ( .A(n902), .B(n725), .Y(n320) );
  OAI221XL U814 ( .A0(n726), .A1(n791), .B0(n731), .B1(n788), .C0(n903), .Y(
        n902) );
  AOI22X1 U815 ( .A0(a[8]), .A1(n733), .B0(a[7]), .B1(n709), .Y(n903) );
  XNOR2X1 U816 ( .A(n904), .B(n725), .Y(n319) );
  OAI221XL U817 ( .A0(n726), .A1(n789), .B0(n731), .B1(n786), .C0(n905), .Y(
        n904) );
  AOI22X1 U818 ( .A0(a[9]), .A1(n733), .B0(a[8]), .B1(n709), .Y(n905) );
  XNOR2X1 U819 ( .A(n906), .B(n725), .Y(n318) );
  OAI221XL U820 ( .A0(n726), .A1(n787), .B0(n731), .B1(n784), .C0(n907), .Y(
        n906) );
  AOI22X1 U821 ( .A0(a[10]), .A1(n733), .B0(a[9]), .B1(n710), .Y(n907) );
  XNOR2X1 U822 ( .A(n908), .B(n725), .Y(n317) );
  OAI221XL U823 ( .A0(n726), .A1(n785), .B0(n731), .B1(n782), .C0(n909), .Y(
        n908) );
  AOI22X1 U824 ( .A0(a[11]), .A1(n733), .B0(a[10]), .B1(n710), .Y(n909) );
  XNOR2X1 U825 ( .A(n910), .B(n725), .Y(n316) );
  OAI221XL U826 ( .A0(n726), .A1(n783), .B0(n729), .B1(n780), .C0(n911), .Y(
        n910) );
  AOI22X1 U827 ( .A0(a[12]), .A1(n733), .B0(a[11]), .B1(n710), .Y(n911) );
  XNOR2X1 U828 ( .A(n912), .B(n725), .Y(n315) );
  OAI221XL U829 ( .A0(n726), .A1(n781), .B0(n729), .B1(n778), .C0(n913), .Y(
        n912) );
  AOI22X1 U830 ( .A0(a[13]), .A1(n734), .B0(a[12]), .B1(n710), .Y(n913) );
  XNOR2X1 U831 ( .A(n914), .B(n725), .Y(n314) );
  OAI221XL U832 ( .A0(n727), .A1(n779), .B0(n729), .B1(n776), .C0(n915), .Y(
        n914) );
  AOI22X1 U833 ( .A0(a[14]), .A1(n734), .B0(a[13]), .B1(n710), .Y(n915) );
  XNOR2X1 U834 ( .A(n916), .B(n725), .Y(n313) );
  OAI221XL U835 ( .A0(n727), .A1(n777), .B0(n820), .B1(n774), .C0(n917), .Y(
        n916) );
  AOI22X1 U836 ( .A0(a[15]), .A1(n734), .B0(a[14]), .B1(n710), .Y(n917) );
  XNOR2X1 U837 ( .A(n918), .B(n724), .Y(n312) );
  OAI221XL U838 ( .A0(n727), .A1(n775), .B0(n820), .B1(n772), .C0(n919), .Y(
        n918) );
  AOI22X1 U839 ( .A0(a[16]), .A1(n734), .B0(a[15]), .B1(n710), .Y(n919) );
  XNOR2X1 U840 ( .A(n920), .B(n724), .Y(n311) );
  OAI221XL U841 ( .A0(n727), .A1(n773), .B0(n820), .B1(n770), .C0(n921), .Y(
        n920) );
  AOI22X1 U842 ( .A0(a[17]), .A1(n734), .B0(a[16]), .B1(n710), .Y(n921) );
  XNOR2X1 U843 ( .A(n922), .B(n724), .Y(n310) );
  OAI221XL U844 ( .A0(n727), .A1(n771), .B0(n820), .B1(n768), .C0(n923), .Y(
        n922) );
  AOI22X1 U845 ( .A0(a[18]), .A1(n734), .B0(a[17]), .B1(n710), .Y(n923) );
  XNOR2X1 U846 ( .A(n924), .B(n724), .Y(n309) );
  OAI221XL U847 ( .A0(n727), .A1(n769), .B0(n731), .B1(n766), .C0(n925), .Y(
        n924) );
  AOI22X1 U848 ( .A0(a[19]), .A1(n734), .B0(a[18]), .B1(n710), .Y(n925) );
  XNOR2X1 U849 ( .A(n926), .B(n724), .Y(n308) );
  OAI221XL U850 ( .A0(n727), .A1(n767), .B0(n731), .B1(n764), .C0(n927), .Y(
        n926) );
  AOI22X1 U851 ( .A0(a[20]), .A1(n734), .B0(a[19]), .B1(n710), .Y(n927) );
  XNOR2X1 U852 ( .A(n928), .B(n724), .Y(n307) );
  OAI221XL U853 ( .A0(n727), .A1(n765), .B0(n731), .B1(n762), .C0(n929), .Y(
        n928) );
  AOI22X1 U854 ( .A0(a[20]), .A1(n709), .B0(n733), .B1(a[21]), .Y(n929) );
  XNOR2X1 U855 ( .A(n930), .B(n724), .Y(n306) );
  OAI221XL U856 ( .A0(n727), .A1(n763), .B0(n761), .B1(n931), .C0(n932), .Y(
        n930) );
  AOI22X1 U857 ( .A0(n734), .A1(a[22]), .B0(n251), .B1(n730), .Y(n932) );
  XNOR2X1 U858 ( .A(n933), .B(n724), .Y(n305) );
  OAI221XL U859 ( .A0(n761), .A1(n727), .B0(n759), .B1(n699), .C0(n934), .Y(
        n933) );
  AOI22X1 U860 ( .A0(n709), .A1(a[22]), .B0(n250), .B1(n730), .Y(n934) );
  XNOR2X1 U861 ( .A(n935), .B(n724), .Y(n304) );
  OAI221XL U862 ( .A0(n760), .A1(n727), .B0(n731), .B1(n758), .C0(n936), .Y(
        n935) );
  AOI22X1 U863 ( .A0(n734), .A1(a[24]), .B0(n710), .B1(a[23]), .Y(n936) );
  XNOR2X1 U864 ( .A(n937), .B(n724), .Y(n303) );
  OAI221XL U865 ( .A0(n757), .A1(n931), .B0(n759), .B1(n727), .C0(n938), .Y(
        n937) );
  AOI22X1 U866 ( .A0(n734), .A1(a[25]), .B0(n730), .B1(n248), .Y(n938) );
  XNOR2X1 U867 ( .A(n939), .B(n724), .Y(n302) );
  OAI221XL U868 ( .A0(n757), .A1(n727), .B0(n699), .B1(n754), .C0(n940), .Y(
        n939) );
  AOI22X1 U869 ( .A0(n709), .A1(a[25]), .B0(n247), .B1(n732), .Y(n940) );
  XNOR2X1 U870 ( .A(n941), .B(n724), .Y(n301) );
  OAI221XL U871 ( .A0(n755), .A1(n727), .B0(n731), .B1(n753), .C0(n942), .Y(
        n941) );
  AOI22X1 U872 ( .A0(a[27]), .A1(n733), .B0(a[26]), .B1(n709), .Y(n942) );
  NAND2X1 U873 ( .A(n943), .B(b[3]), .Y(n931) );
  NAND2BX1 U874 ( .AN(n943), .B(n19), .Y(n820) );
  NAND3BX1 U875 ( .AN(b[3]), .B(n943), .C(n19), .Y(n819) );
  XNOR2X1 U876 ( .A(b[3]), .B(b[2]), .Y(n943) );
  AOI22X1 U877 ( .A0(a[0]), .A1(n802), .B0(a[0]), .B1(n739), .Y(n153) );
  OAI221XL U878 ( .A0(n735), .A1(n706), .B0(n705), .B1(n800), .C0(n945), .Y(
        n944) );
  AOI22X1 U879 ( .A0(a[2]), .A1(n738), .B0(a[1]), .B1(n720), .Y(n945) );
  OAI221XL U880 ( .A0(n735), .A1(n801), .B0(n705), .B1(n798), .C0(n947), .Y(
        n946) );
  AOI22X1 U881 ( .A0(a[3]), .A1(n738), .B0(a[2]), .B1(n720), .Y(n947) );
  OAI221XL U882 ( .A0(n735), .A1(n799), .B0(n705), .B1(n796), .C0(n949), .Y(
        n948) );
  AOI22X1 U883 ( .A0(a[4]), .A1(n738), .B0(a[3]), .B1(n720), .Y(n949) );
  OAI221XL U884 ( .A0(n735), .A1(n797), .B0(n705), .B1(n794), .C0(n951), .Y(
        n950) );
  AOI22X1 U885 ( .A0(a[5]), .A1(n738), .B0(a[4]), .B1(n720), .Y(n951) );
  OAI221XL U886 ( .A0(n735), .A1(n795), .B0(n705), .B1(n792), .C0(n953), .Y(
        n952) );
  AOI22X1 U887 ( .A0(a[6]), .A1(n738), .B0(a[5]), .B1(n720), .Y(n953) );
  OAI221XL U888 ( .A0(n735), .A1(n793), .B0(n705), .B1(n790), .C0(n955), .Y(
        n954) );
  AOI22X1 U889 ( .A0(a[7]), .A1(n738), .B0(a[6]), .B1(n720), .Y(n955) );
  OAI221XL U890 ( .A0(n735), .A1(n791), .B0(n705), .B1(n788), .C0(n957), .Y(
        n956) );
  AOI22X1 U891 ( .A0(a[8]), .A1(n738), .B0(a[7]), .B1(n720), .Y(n957) );
  OAI221XL U892 ( .A0(n735), .A1(n789), .B0(n705), .B1(n786), .C0(n959), .Y(
        n958) );
  AOI22X1 U893 ( .A0(a[9]), .A1(n738), .B0(a[8]), .B1(n720), .Y(n959) );
  OAI221XL U894 ( .A0(n735), .A1(n787), .B0(n705), .B1(n784), .C0(n961), .Y(
        n960) );
  AOI22X1 U895 ( .A0(a[10]), .A1(n738), .B0(a[9]), .B1(n720), .Y(n961) );
  OAI221XL U896 ( .A0(n735), .A1(n785), .B0(n705), .B1(n782), .C0(n963), .Y(
        n962) );
  AOI22X1 U897 ( .A0(a[11]), .A1(n738), .B0(a[10]), .B1(n721), .Y(n963) );
  OAI221XL U898 ( .A0(n735), .A1(n783), .B0(n705), .B1(n780), .C0(n965), .Y(
        n964) );
  AOI22X1 U899 ( .A0(a[12]), .A1(n739), .B0(a[11]), .B1(n721), .Y(n965) );
  OAI221XL U900 ( .A0(n736), .A1(n781), .B0(n705), .B1(n778), .C0(n967), .Y(
        n966) );
  AOI22X1 U901 ( .A0(a[13]), .A1(n739), .B0(a[12]), .B1(n721), .Y(n967) );
  OAI221XL U902 ( .A0(n736), .A1(n779), .B0(n705), .B1(n776), .C0(n969), .Y(
        n968) );
  AOI22X1 U903 ( .A0(a[14]), .A1(n739), .B0(a[13]), .B1(n721), .Y(n969) );
  OAI221XL U904 ( .A0(n736), .A1(n777), .B0(n705), .B1(n774), .C0(n971), .Y(
        n970) );
  AOI22X1 U905 ( .A0(a[15]), .A1(n739), .B0(a[14]), .B1(n721), .Y(n971) );
  OAI221XL U906 ( .A0(n736), .A1(n775), .B0(n705), .B1(n772), .C0(n973), .Y(
        n972) );
  AOI22X1 U907 ( .A0(a[16]), .A1(n739), .B0(a[15]), .B1(n721), .Y(n973) );
  OAI221XL U908 ( .A0(n736), .A1(n773), .B0(n705), .B1(n770), .C0(n975), .Y(
        n974) );
  AOI22X1 U909 ( .A0(a[17]), .A1(n739), .B0(a[16]), .B1(n721), .Y(n975) );
  OAI221XL U910 ( .A0(n736), .A1(n771), .B0(n705), .B1(n768), .C0(n977), .Y(
        n976) );
  AOI22X1 U911 ( .A0(a[18]), .A1(n739), .B0(a[17]), .B1(n721), .Y(n977) );
  OAI221XL U912 ( .A0(n736), .A1(n769), .B0(n705), .B1(n766), .C0(n979), .Y(
        n978) );
  AOI22X1 U913 ( .A0(a[19]), .A1(n739), .B0(a[18]), .B1(n721), .Y(n979) );
  OAI221XL U914 ( .A0(n736), .A1(n767), .B0(n705), .B1(n764), .C0(n981), .Y(
        n980) );
  AOI22X1 U915 ( .A0(a[20]), .A1(n739), .B0(a[19]), .B1(n721), .Y(n981) );
  OAI221XL U916 ( .A0(n736), .A1(n765), .B0(n705), .B1(n762), .C0(n983), .Y(
        n982) );
  AOI22X1 U917 ( .A0(a[20]), .A1(n720), .B0(n739), .B1(a[21]), .Y(n983) );
  OAI221XL U918 ( .A0(n736), .A1(n763), .B0(n761), .B1(n985), .C0(n986), .Y(
        n984) );
  AOI22X1 U919 ( .A0(n739), .A1(a[22]), .B0(n251), .B1(n802), .Y(n986) );
  OAI221XL U920 ( .A0(n761), .A1(n736), .B0(n700), .B1(n759), .C0(n988), .Y(
        n987) );
  AOI22X1 U921 ( .A0(n720), .A1(a[22]), .B0(n250), .B1(n802), .Y(n988) );
  OAI221XL U922 ( .A0(n760), .A1(n736), .B0(n705), .B1(n758), .C0(n990), .Y(
        n989) );
  AOI22X1 U923 ( .A0(a[24]), .A1(n738), .B0(a[23]), .B1(n720), .Y(n990) );
  NAND2X1 U924 ( .A(n991), .B(n992), .Y(n985) );
  NAND3BX1 U925 ( .AN(n992), .B(n991), .C(n993), .Y(n823) );
  XNOR2X1 U926 ( .A(b[6]), .B(n19), .Y(n991) );
  XOR2X1 U927 ( .A(b[6]), .B(b[7]), .Y(n992) );
endmodule


module Equation_Implementation_DW01_sub_8 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7;
  wire   [7:0] carry;

  ADDFX2 U2_1 ( .A(A[1]), .B(n6), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n3), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFX2 U2_3 ( .A(A[3]), .B(n4), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFX2 U2_2 ( .A(A[2]), .B(n5), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFX2 U2_5 ( .A(A[5]), .B(n2), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  INVXL U1 ( .A(B[0]), .Y(n7) );
  INVX1 U2 ( .A(carry[6]), .Y(DIFF[6]) );
  INVX1 U3 ( .A(B[5]), .Y(n2) );
  INVX1 U4 ( .A(B[2]), .Y(n5) );
  INVX1 U5 ( .A(B[3]), .Y(n4) );
  INVX1 U6 ( .A(B[4]), .Y(n3) );
  INVX1 U7 ( .A(B[1]), .Y(n6) );
  OR2X2 U8 ( .A(A[0]), .B(n7), .Y(carry[1]) );
  XNOR2X1 U9 ( .A(n7), .B(A[0]), .Y(DIFF[0]) );
endmodule


module Equation_Implementation_DW_mult_uns_10 ( a, b, product );
  input [31:0] a;
  input [9:0] b;
  output [41:0] product;
  wire   n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n173, n174, n175, n176, n177, n240, n241, \product[29] ,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262;
  assign product[28] = \product[29] ;
  assign product[24] = \product[29] ;
  assign product[22] = \product[29] ;
  assign product[18] = \product[29] ;
  assign product[19] = \product[29] ;
  assign product[31] = \product[29] ;
  assign product[21] = \product[29] ;
  assign product[25] = \product[29] ;
  assign product[27] = \product[29] ;
  assign product[30] = \product[29] ;
  assign product[17] = \product[29] ;
  assign product[16] = \product[29] ;
  assign product[20] = \product[29] ;
  assign product[29] = \product[29] ;

  ADDFX2 U28 ( .A(n35), .B(n109), .CI(n21), .CO(n20), .S(product[15]) );
  ADDFX2 U29 ( .A(n38), .B(n36), .CI(n22), .CO(n21), .S(product[14]) );
  ADDFX2 U30 ( .A(n39), .B(n41), .CI(n23), .CO(n22), .S(product[13]) );
  ADDFX2 U31 ( .A(n42), .B(n46), .CI(n24), .CO(n23), .S(product[12]) );
  ADDFX2 U32 ( .A(n47), .B(n52), .CI(n25), .CO(n24), .S(product[11]) );
  ADDFX2 U33 ( .A(n53), .B(n60), .CI(n26), .CO(n25), .S(product[10]) );
  ADDFX2 U34 ( .A(n61), .B(n68), .CI(n27), .CO(n26), .S(product[9]) );
  ADDFX2 U35 ( .A(n69), .B(n76), .CI(n28), .CO(n27), .S(product[8]) );
  ADDFX2 U36 ( .A(n77), .B(n84), .CI(n29), .CO(n28), .S(product[7]) );
  ADDFX2 U37 ( .A(n85), .B(n92), .CI(n30), .CO(n29), .S(product[6]) );
  ADDFX2 U38 ( .A(n93), .B(n99), .CI(n31), .CO(n30), .S(product[5]) );
  ADDFX2 U39 ( .A(n100), .B(n103), .CI(n32), .CO(n31), .S(product[4]) );
  ADDFX2 U40 ( .A(n104), .B(n106), .CI(n33), .CO(n32), .S(product[3]) );
  ADDFX2 U41 ( .A(n34), .B(n164), .CI(n108), .CO(n33), .S(product[2]) );
  ADDHXL U42 ( .A(n171), .B(n177), .CO(n34), .S(product[1]) );
  ADDFX2 U43 ( .A(n110), .B(n116), .CI(n37), .CO(n35), .S(n36) );
  CMPR42X1 U44 ( .A(n117), .B(n123), .C(n43), .D(n111), .ICI(n40), .S(n39), 
        .ICO(n37), .CO(n38) );
  CMPR42X1 U45 ( .A(n48), .B(n112), .C(n49), .D(n44), .ICI(n45), .S(n42), 
        .ICO(n40), .CO(n41) );
  ADDFX2 U46 ( .A(n118), .B(n130), .CI(n124), .CO(n43), .S(n44) );
  CMPR42X1 U47 ( .A(n57), .B(n54), .C(n55), .D(n50), .ICI(n51), .S(n47), .ICO(
        n45), .CO(n46) );
  CMPR42X1 U48 ( .A(n119), .B(n137), .C(n113), .D(n125), .ICI(n131), .S(n50), 
        .ICO(n48), .CO(n49) );
  CMPR42X1 U49 ( .A(n58), .B(n65), .C(n56), .D(n63), .ICI(n59), .S(n53), .ICO(
        n51), .CO(n52) );
  CMPR42X1 U50 ( .A(n138), .B(n120), .C(n114), .D(n132), .ICI(n62), .S(n56), 
        .ICO(n54), .CO(n55) );
  ADDHXL U51 ( .A(n144), .B(n126), .CO(n57), .S(n58) );
  CMPR42X1 U52 ( .A(n66), .B(n73), .C(n64), .D(n71), .ICI(n67), .S(n61), .ICO(
        n59), .CO(n60) );
  CMPR42X1 U53 ( .A(n145), .B(n127), .C(n115), .D(n139), .ICI(n70), .S(n64), 
        .ICO(n62), .CO(n63) );
  ADDFX2 U54 ( .A(n121), .B(n151), .CI(n133), .CO(n65), .S(n66) );
  CMPR42X1 U55 ( .A(n74), .B(n81), .C(n72), .D(n79), .ICI(n75), .S(n69), .ICO(
        n67), .CO(n68) );
  CMPR42X1 U56 ( .A(n152), .B(n134), .C(n122), .D(n146), .ICI(n78), .S(n72), 
        .ICO(n70), .CO(n71) );
  ADDFX2 U57 ( .A(n128), .B(n158), .CI(n140), .CO(n73), .S(n74) );
  CMPR42X1 U58 ( .A(n82), .B(n86), .C(n80), .D(n87), .ICI(n83), .S(n77), .ICO(
        n75), .CO(n76) );
  CMPR42X1 U59 ( .A(n129), .B(n153), .C(n141), .D(n147), .ICI(n89), .S(n80), 
        .ICO(n78), .CO(n79) );
  ADDFX2 U60 ( .A(n135), .B(n165), .CI(n159), .CO(n81), .S(n82) );
  CMPR42X1 U61 ( .A(n94), .B(n96), .C(n90), .D(n88), .ICI(n91), .S(n85), .ICO(
        n83), .CO(n84) );
  CMPR42X1 U62 ( .A(n136), .B(n166), .C(n154), .D(n148), .ICI(n160), .S(n88), 
        .ICO(n86), .CO(n87) );
  CMPR42X1 U65 ( .A(n101), .B(n167), .C(n97), .D(n95), .ICI(n98), .S(n93), 
        .ICO(n91), .CO(n92) );
  ADDFX2 U66 ( .A(n155), .B(n173), .CI(n161), .CO(n94), .S(n95) );
  ADDHXL U67 ( .A(n149), .B(n143), .CO(n96), .S(n97) );
  CMPR42X1 U68 ( .A(n162), .B(n174), .C(n105), .D(n168), .ICI(n102), .S(n100), 
        .ICO(n98), .CO(n99) );
  ADDHXL U69 ( .A(n156), .B(n150), .CO(n101), .S(n102) );
  ADDFX2 U70 ( .A(n169), .B(n175), .CI(n107), .CO(n103), .S(n104) );
  ADDHXL U71 ( .A(n163), .B(n157), .CO(n105), .S(n106) );
  ADDHXL U72 ( .A(n176), .B(n170), .CO(n107), .S(n108) );
  BUFX3 U162 ( .A(a[6]), .Y(n241) );
  CLKINVX3 U163 ( .A(a[2]), .Y(n249) );
  CLKINVX3 U164 ( .A(a[5]), .Y(n246) );
  CLKINVX3 U165 ( .A(a[4]), .Y(n247) );
  CLKINVX3 U166 ( .A(a[3]), .Y(n248) );
  BUFX3 U167 ( .A(n250), .Y(n240) );
  INVX1 U168 ( .A(a[1]), .Y(n250) );
  CLKINVX3 U169 ( .A(n243), .Y(\product[29] ) );
  INVX1 U170 ( .A(n245), .Y(n243) );
  INVX1 U171 ( .A(n20), .Y(n245) );
  CLKINVX3 U172 ( .A(a[0]), .Y(n251) );
  CLKINVX3 U173 ( .A(b[2]), .Y(n259) );
  CLKINVX3 U174 ( .A(b[1]), .Y(n260) );
  CLKINVX3 U175 ( .A(b[6]), .Y(n255) );
  CLKINVX3 U176 ( .A(b[3]), .Y(n258) );
  CLKINVX3 U177 ( .A(b[4]), .Y(n257) );
  INVX1 U178 ( .A(b[5]), .Y(n256) );
  CLKINVX3 U179 ( .A(b[0]), .Y(n244) );
  CLKINVX3 U180 ( .A(b[7]), .Y(n254) );
  CLKINVX3 U181 ( .A(b[9]), .Y(n252) );
  CLKINVX3 U182 ( .A(b[8]), .Y(n253) );
  NOR2X1 U183 ( .A(n251), .B(n244), .Y(product[0]) );
  XNOR2X1 U184 ( .A(n261), .B(n262), .Y(n90) );
  NAND2X1 U185 ( .A(n262), .B(n261), .Y(n89) );
  NAND2X1 U186 ( .A(b[5]), .B(a[1]), .Y(n261) );
  NOR2BX1 U187 ( .AN(n241), .B(n244), .Y(n262) );
  NOR2X1 U188 ( .A(n244), .B(n240), .Y(n177) );
  NOR2X1 U189 ( .A(n244), .B(n249), .Y(n176) );
  NOR2X1 U190 ( .A(n244), .B(n248), .Y(n175) );
  NOR2X1 U191 ( .A(n244), .B(n247), .Y(n174) );
  NOR2X1 U192 ( .A(n244), .B(n246), .Y(n173) );
  NOR2X1 U193 ( .A(n251), .B(n260), .Y(n171) );
  NOR2X1 U194 ( .A(n240), .B(n260), .Y(n170) );
  NOR2X1 U195 ( .A(n249), .B(n260), .Y(n169) );
  NOR2X1 U196 ( .A(n248), .B(n260), .Y(n168) );
  NOR2X1 U197 ( .A(n247), .B(n260), .Y(n167) );
  NOR2X1 U198 ( .A(n246), .B(n260), .Y(n166) );
  NAND2X1 U199 ( .A(b[1]), .B(n241), .Y(n165) );
  NOR2X1 U200 ( .A(n251), .B(n259), .Y(n164) );
  NOR2X1 U201 ( .A(n240), .B(n259), .Y(n163) );
  NOR2X1 U202 ( .A(n249), .B(n259), .Y(n162) );
  NOR2X1 U203 ( .A(n248), .B(n259), .Y(n161) );
  NOR2X1 U204 ( .A(n247), .B(n259), .Y(n160) );
  NOR2X1 U205 ( .A(n246), .B(n259), .Y(n159) );
  NAND2X1 U206 ( .A(b[2]), .B(n241), .Y(n158) );
  NOR2X1 U207 ( .A(n251), .B(n258), .Y(n157) );
  NOR2X1 U208 ( .A(n240), .B(n258), .Y(n156) );
  NOR2X1 U209 ( .A(n249), .B(n258), .Y(n155) );
  NOR2X1 U210 ( .A(n248), .B(n258), .Y(n154) );
  NOR2X1 U211 ( .A(n247), .B(n258), .Y(n153) );
  NOR2X1 U212 ( .A(n246), .B(n258), .Y(n152) );
  NAND2X1 U213 ( .A(b[3]), .B(n241), .Y(n151) );
  NOR2X1 U214 ( .A(n251), .B(n257), .Y(n150) );
  NOR2X1 U215 ( .A(n240), .B(n257), .Y(n149) );
  NOR2X1 U216 ( .A(n249), .B(n257), .Y(n148) );
  NOR2X1 U217 ( .A(n248), .B(n257), .Y(n147) );
  NOR2X1 U218 ( .A(n247), .B(n257), .Y(n146) );
  NOR2X1 U219 ( .A(n246), .B(n257), .Y(n145) );
  NAND2X1 U220 ( .A(b[4]), .B(n241), .Y(n144) );
  NOR2X1 U221 ( .A(n251), .B(n256), .Y(n143) );
  NOR2X1 U222 ( .A(n256), .B(n249), .Y(n141) );
  NOR2X1 U223 ( .A(n256), .B(n248), .Y(n140) );
  NOR2X1 U224 ( .A(n256), .B(n247), .Y(n139) );
  NOR2X1 U225 ( .A(n256), .B(n246), .Y(n138) );
  NAND2X1 U226 ( .A(n241), .B(b[5]), .Y(n137) );
  NOR2X1 U227 ( .A(n251), .B(n255), .Y(n136) );
  NOR2X1 U228 ( .A(n240), .B(n255), .Y(n135) );
  NOR2X1 U229 ( .A(n249), .B(n255), .Y(n134) );
  NOR2X1 U230 ( .A(n248), .B(n255), .Y(n133) );
  NOR2X1 U231 ( .A(n247), .B(n255), .Y(n132) );
  NOR2X1 U232 ( .A(n246), .B(n255), .Y(n131) );
  NAND2X1 U233 ( .A(b[6]), .B(n241), .Y(n130) );
  NOR2X1 U234 ( .A(n251), .B(n254), .Y(n129) );
  NOR2X1 U235 ( .A(n240), .B(n254), .Y(n128) );
  NOR2X1 U236 ( .A(n249), .B(n254), .Y(n127) );
  NOR2X1 U237 ( .A(n248), .B(n254), .Y(n126) );
  NOR2X1 U238 ( .A(n247), .B(n254), .Y(n125) );
  NOR2X1 U239 ( .A(n246), .B(n254), .Y(n124) );
  NAND2X1 U240 ( .A(b[7]), .B(n241), .Y(n123) );
  NOR2X1 U241 ( .A(n251), .B(n253), .Y(n122) );
  NOR2X1 U242 ( .A(n240), .B(n253), .Y(n121) );
  NOR2X1 U243 ( .A(n249), .B(n253), .Y(n120) );
  NOR2X1 U244 ( .A(n248), .B(n253), .Y(n119) );
  NOR2X1 U245 ( .A(n247), .B(n253), .Y(n118) );
  NOR2X1 U246 ( .A(n246), .B(n253), .Y(n117) );
  NAND2X1 U247 ( .A(b[8]), .B(n241), .Y(n116) );
  NOR2X1 U248 ( .A(n251), .B(n252), .Y(n115) );
  NOR2X1 U249 ( .A(n240), .B(n252), .Y(n114) );
  NOR2X1 U250 ( .A(n249), .B(n252), .Y(n113) );
  NOR2X1 U251 ( .A(n248), .B(n252), .Y(n112) );
  NOR2X1 U252 ( .A(n247), .B(n252), .Y(n111) );
  NOR2X1 U253 ( .A(n246), .B(n252), .Y(n110) );
  NAND2X1 U254 ( .A(b[9]), .B(n241), .Y(n109) );
endmodule


module Equation_Implementation_DW_mult_uns_9 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n74, n79, n80, n81, n88, n89, n94, n95, n96, n98, n100,
         n101, n102, n108, n109, n114, n115, n116, n118, n120, n121, n122,
         n127, n128, n129, n130, n132, n134, n135, n136, n138, n140, n141,
         n142, n143, n144, n147, n148, n149, n150, n151, n152, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n167,
         n168, n169, n170, n171, n172, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n187, n188, n189, n190, n191,
         n192, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n706, n708, n709, n710, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103;
  assign n79 = a[29];
  assign n132 = a[20];
  assign n706 = a[17];
  assign n708 = a[11];
  assign n709 = a[8];
  assign n710 = a[5];

  ADDFX2 U34 ( .A(n880), .B(n81), .CI(n37), .CO(n36), .S(product[30]) );
  ADDFX2 U35 ( .A(n876), .B(n88), .CI(n38), .CO(n37), .S(product[29]) );
  ADDFX2 U36 ( .A(n95), .B(n89), .CI(n39), .CO(n38), .S(product[28]) );
  ADDFX2 U37 ( .A(n96), .B(n101), .CI(n40), .CO(n39), .S(product[27]) );
  ADDFX2 U38 ( .A(n102), .B(n108), .CI(n41), .CO(n40), .S(product[26]) );
  ADDFX2 U39 ( .A(n115), .B(n109), .CI(n42), .CO(n41), .S(product[25]) );
  ADDFX2 U40 ( .A(n116), .B(n121), .CI(n43), .CO(n42), .S(product[24]) );
  ADDFX2 U41 ( .A(n122), .B(n128), .CI(n44), .CO(n43), .S(product[23]) );
  ADDFX2 U42 ( .A(n135), .B(n129), .CI(n45), .CO(n44), .S(product[22]) );
  ADDFX2 U43 ( .A(n136), .B(n141), .CI(n46), .CO(n45), .S(product[21]) );
  ADDFX2 U44 ( .A(n142), .B(n148), .CI(n47), .CO(n46), .S(product[20]) );
  ADDFX2 U45 ( .A(n155), .B(n149), .CI(n48), .CO(n47), .S(product[19]) );
  ADDFX2 U46 ( .A(n156), .B(n161), .CI(n49), .CO(n48), .S(product[18]) );
  ADDFX2 U47 ( .A(n162), .B(n168), .CI(n50), .CO(n49), .S(product[17]) );
  ADDFX2 U48 ( .A(n175), .B(n169), .CI(n51), .CO(n50), .S(product[16]) );
  ADDFX2 U49 ( .A(n176), .B(n181), .CI(n52), .CO(n51), .S(product[15]) );
  ADDFX2 U50 ( .A(n182), .B(n188), .CI(n53), .CO(n52), .S(product[14]) );
  ADDFX2 U51 ( .A(n189), .B(n195), .CI(n54), .CO(n53), .S(product[13]) );
  ADDFX2 U52 ( .A(n196), .B(n202), .CI(n55), .CO(n54), .S(product[12]) );
  ADDFX2 U53 ( .A(n203), .B(n207), .CI(n56), .CO(n55), .S(product[11]) );
  ADDFX2 U54 ( .A(n208), .B(n212), .CI(n57), .CO(n56), .S(product[10]) );
  ADDFX2 U55 ( .A(n213), .B(n372), .CI(n58), .CO(n57), .S(product[9]) );
  ADDFX2 U56 ( .A(n217), .B(n373), .CI(n59), .CO(n58), .S(product[8]) );
  ADDFX2 U57 ( .A(n221), .B(n224), .CI(n60), .CO(n59), .S(product[7]) );
  ADDFX2 U58 ( .A(n225), .B(n228), .CI(n61), .CO(n60), .S(product[6]) );
  ADDFX2 U59 ( .A(n229), .B(n230), .CI(n62), .CO(n61), .S(product[5]) );
  ADDFX2 U60 ( .A(n231), .B(n367), .CI(n63), .CO(n62), .S(product[4]) );
  ADDFX2 U61 ( .A(n233), .B(n378), .CI(n64), .CO(n63), .S(product[3]) );
  ADDHXL U62 ( .A(n379), .B(n65), .CO(n64), .S(product[2]) );
  ADDHXL U63 ( .A(n66), .B(n380), .CO(n65), .S(product[1]) );
  CMPR42X1 U71 ( .A(n876), .B(a[27]), .C(a[23]), .D(a[27]), .ICI(n80), .CO(n74) );
  CMPR42X1 U74 ( .A(n875), .B(n130), .C(n130), .D(a[23]), .ICI(a[28]), .ICO(
        n80), .CO(n81) );
  CMPR42X1 U77 ( .A(a[26]), .B(n875), .C(n132), .D(n98), .ICI(n94), .S(n89), 
        .CO(n88) );
  CMPR42X1 U80 ( .A(n309), .B(a[27]), .C(n132), .D(a[30]), .ICI(n100), .S(n96), 
        .ICO(n94), .CO(n95) );
  CMPR42X1 U81 ( .A(n130), .B(n130), .C(a[30]), .D(a[28]), .ICI(n309), .CO(n98) );
  CMPR42X1 U82 ( .A(n872), .B(n130), .C(n310), .D(a[26]), .ICI(n311), .S(n102), 
        .ICO(n100), .CO(n101) );
  CMPR42X1 U85 ( .A(n132), .B(n872), .C(n311), .D(n118), .ICI(n114), .S(n109), 
        .CO(n108) );
  CMPR42X1 U88 ( .A(n320), .B(a[23]), .C(n312), .D(a[31]), .ICI(n120), .S(n116), .ICO(n114), .CO(n115) );
  CMPR42X1 U89 ( .A(n130), .B(a[31]), .C(a[30]), .D(a[28]), .ICI(n320), .CO(
        n118) );
  CMPR42X1 U90 ( .A(n872), .B(n130), .C(n321), .D(n313), .ICI(n127), .S(n122), 
        .ICO(n120), .CO(n121) );
  CMPR42X1 U93 ( .A(n314), .B(n876), .C(n322), .D(n138), .ICI(n134), .S(n129), 
        .ICO(n127), .CO(n128) );
  CMPR42X1 U96 ( .A(n331), .B(n315), .C(n323), .D(n143), .ICI(n140), .S(n136), 
        .ICO(n134), .CO(n135) );
  CMPR42X1 U97 ( .A(n130), .B(a[31]), .C(a[23]), .D(a[23]), .ICI(n331), .CO(
        n138) );
  CMPR42X1 U98 ( .A(n144), .B(n150), .C(n332), .D(n324), .ICI(n147), .S(n142), 
        .ICO(n140), .CO(n141) );
  ADDFX2 U99 ( .A(n316), .B(n152), .CI(n876), .CO(n143), .S(n144) );
  CMPR42X1 U101 ( .A(n325), .B(n881), .C(n333), .D(n151), .ICI(n154), .S(n149), 
        .ICO(n147), .CO(n148) );
  ADDFX2 U102 ( .A(n157), .B(n130), .CI(n158), .CO(n150), .S(n151) );
  CMPR42X1 U104 ( .A(n159), .B(n326), .C(n334), .D(n163), .ICI(n160), .S(n156), 
        .ICO(n154), .CO(n155) );
  CMPR42X1 U105 ( .A(n130), .B(a[26]), .C(n317), .D(n165), .ICI(n343), .S(n159), .ICO(n157), .CO(n158) );
  CMPR42X1 U106 ( .A(n164), .B(n170), .C(n344), .D(n335), .ICI(n167), .S(n162), 
        .ICO(n160), .CO(n161) );
  ADDFX2 U107 ( .A(n327), .B(n172), .CI(n882), .CO(n163), .S(n164) );
  CMPR42X1 U109 ( .A(n336), .B(n889), .C(n345), .D(n171), .ICI(n174), .S(n169), 
        .ICO(n167), .CO(n168) );
  ADDFX2 U110 ( .A(n177), .B(n318), .CI(n178), .CO(n170), .S(n171) );
  CMPR42X1 U112 ( .A(n179), .B(n337), .C(n346), .D(n183), .ICI(n180), .S(n176), 
        .ICO(n174), .CO(n175) );
  CMPR42X1 U113 ( .A(n319), .B(n874), .C(n328), .D(n185), .ICI(n356), .S(n179), 
        .ICO(n177), .CO(n178) );
  CMPR42X1 U114 ( .A(n190), .B(n184), .C(n357), .D(n347), .ICI(n187), .S(n182), 
        .ICO(n180), .CO(n181) );
  ADDFX2 U115 ( .A(n338), .B(n192), .CI(n888), .CO(n183), .S(n184) );
  CMPR42X1 U117 ( .A(n197), .B(n348), .C(n358), .D(n191), .ICI(n194), .S(n189), 
        .ICO(n187), .CO(n188) );
  ADDFX2 U118 ( .A(n329), .B(n199), .CI(n894), .CO(n190), .S(n191) );
  CMPR42X1 U120 ( .A(n204), .B(n200), .C(n359), .D(n198), .ICI(n201), .S(n196), 
        .ICO(n194), .CO(n195) );
  ADDFX2 U121 ( .A(n339), .B(n369), .CI(n349), .CO(n197), .S(n198) );
  CMPR42X1 U124 ( .A(n205), .B(n209), .C(n206), .D(n360), .ICI(n370), .S(n203), 
        .ICO(n201), .CO(n202) );
  ADDHXL U125 ( .A(n340), .B(n350), .CO(n204), .S(n205) );
  CMPR42X1 U126 ( .A(n210), .B(n341), .C(n211), .D(n361), .ICI(n371), .S(n208), 
        .ICO(n206), .CO(n207) );
  ADDHXL U127 ( .A(n351), .B(n214), .CO(n209), .S(n210) );
  CMPR42X1 U128 ( .A(n215), .B(n352), .C(n218), .D(n362), .ICI(n216), .S(n213), 
        .ICO(n211), .CO(n212) );
  ADDHXL U129 ( .A(n864), .B(n342), .CO(n214), .S(n215) );
  ADDFX2 U130 ( .A(n219), .B(n222), .CI(n220), .CO(n216), .S(n217) );
  ADDHXL U131 ( .A(n353), .B(n363), .CO(n218), .S(n219) );
  ADDFX2 U132 ( .A(n223), .B(n354), .CI(n374), .CO(n220), .S(n221) );
  ADDHXL U133 ( .A(n364), .B(n226), .CO(n222), .S(n223) );
  ADDFX2 U134 ( .A(n227), .B(n365), .CI(n375), .CO(n224), .S(n225) );
  ADDHXL U135 ( .A(n863), .B(n355), .CO(n226), .S(n227) );
  ADDHXL U136 ( .A(n366), .B(n376), .CO(n228), .S(n229) );
  ADDHXL U137 ( .A(n377), .B(n232), .CO(n230), .S(n231) );
  ADDHXL U138 ( .A(n862), .B(n368), .CO(n232), .S(n233) );
  ADDFX2 U648 ( .A(n859), .B(b[31]), .CI(n256), .CO(n265), .S(n266) );
  ADDFX2 U649 ( .A(b[8]), .B(n859), .CI(n257), .CO(n256), .S(n267) );
  ADDFX2 U650 ( .A(n858), .B(b[8]), .CI(n258), .CO(n257), .S(n268) );
  ADDFX2 U651 ( .A(n857), .B(n858), .CI(n259), .CO(n258), .S(n269) );
  ADDFX2 U652 ( .A(n856), .B(n857), .CI(n260), .CO(n259), .S(n270) );
  ADDFX2 U653 ( .A(b[4]), .B(n856), .CI(n261), .CO(n260), .S(n271) );
  ADDFX2 U654 ( .A(n855), .B(b[4]), .CI(n262), .CO(n261), .S(n272) );
  ADDFX2 U655 ( .A(n854), .B(n855), .CI(n263), .CO(n262), .S(n273) );
  ADDFX2 U656 ( .A(n853), .B(n854), .CI(n264), .CO(n263), .S(n274) );
  XNOR2X1 U660 ( .A(n867), .B(n932), .Y(product[31]) );
  AOI222X1 U661 ( .A0(n897), .A1(n275), .B0(n1024), .B1(n853), .C0(n846), .C1(
        n878), .Y(n1025) );
  CMPR22X1 U662 ( .A(n853), .B(n878), .CO(n264), .S(n275) );
  NAND2X2 U663 ( .A(n1097), .B(n1098), .Y(n1054) );
  CLKINVX3 U664 ( .A(n998), .Y(n900) );
  NAND2X2 U665 ( .A(n1020), .B(n1022), .Y(n998) );
  CLKINVX3 U666 ( .A(n967), .Y(n905) );
  NAND2X2 U667 ( .A(n989), .B(n991), .Y(n967) );
  CLKINVX3 U668 ( .A(n937), .Y(n910) );
  NAND2X2 U669 ( .A(a[0]), .B(n960), .Y(n937) );
  CLKINVX3 U670 ( .A(n1024), .Y(n896) );
  NOR2BX2 U671 ( .AN(n1090), .B(n1091), .Y(n1024) );
  AOI22XL U672 ( .A0(n846), .A1(b[4]), .B0(n897), .B1(n271), .Y(n1033) );
  AOI22XL U673 ( .A0(n1024), .A1(n859), .B0(n846), .B1(n860), .Y(n1042) );
  AOI22XL U674 ( .A0(n1024), .A1(n860), .B0(n846), .B1(n859), .Y(n1044) );
  AOI221XL U675 ( .A0(n905), .A1(b[28]), .B0(n842), .B1(n860), .C0(n988), .Y(
        n987) );
  AOI21XL U676 ( .A0(n899), .A1(n896), .B0(n917), .Y(n1046) );
  AOI22XL U677 ( .A0(n914), .A1(n856), .B0(n270), .B1(n910), .Y(n947) );
  AOI222XL U678 ( .A0(n910), .A1(n275), .B0(n839), .B1(n853), .C0(n914), .C1(
        n878), .Y(n934) );
  AOI22XL U679 ( .A0(n842), .A1(n856), .B0(n905), .B1(n271), .Y(n974) );
  AOI22XL U680 ( .A0(n842), .A1(b[4]), .B0(n840), .B1(n855), .Y(n972) );
  AOI22XL U681 ( .A0(n840), .A1(n856), .B0(n905), .B1(n270), .Y(n976) );
  AOI22XL U682 ( .A0(n845), .A1(n856), .B0(n900), .B1(n271), .Y(n1005) );
  AOI222XL U683 ( .A0(n905), .A1(n275), .B0(n842), .B1(n853), .C0(n840), .C1(
        n878), .Y(n963) );
  AOI22XL U684 ( .A0(n845), .A1(b[4]), .B0(n843), .B1(n855), .Y(n1003) );
  AOI22XL U685 ( .A0(n843), .A1(n856), .B0(n900), .B1(n270), .Y(n1007) );
  AOI22XL U686 ( .A0(n900), .A1(n878), .B0(n845), .B1(n878), .Y(n992) );
  AOI22XL U687 ( .A0(n905), .A1(n878), .B0(n842), .B1(n878), .Y(n961) );
  AOI22XL U688 ( .A0(n1024), .A1(n858), .B0(n846), .B1(n857), .Y(n1038) );
  AOI22XL U689 ( .A0(n897), .A1(n878), .B0(n1024), .B1(n878), .Y(n1023) );
  AOI221XL U690 ( .A0(n839), .A1(n878), .B0(n910), .B1(n878), .C0(n913), .Y(
        n66) );
  AOI22XL U691 ( .A0(n1024), .A1(b[9]), .B0(n846), .B1(n858), .Y(n1040) );
  AOI221XL U692 ( .A0(n897), .A1(n859), .B0(n1024), .B1(n860), .C0(n1048), .Y(
        n1047) );
  AOI22XL U693 ( .A0(n839), .A1(n856), .B0(n271), .B1(n910), .Y(n945) );
  AOI22XL U694 ( .A0(n839), .A1(b[4]), .B0(n914), .B1(n855), .Y(n942) );
  AOI222XL U695 ( .A0(n900), .A1(n275), .B0(n845), .B1(n853), .C0(n843), .C1(
        n878), .Y(n994) );
  CLKINVX3 U696 ( .A(n879), .Y(n878) );
  INVX1 U697 ( .A(b[0]), .Y(n879) );
  INVX1 U698 ( .A(n266), .Y(n918) );
  INVX1 U699 ( .A(n267), .Y(n919) );
  CLKINVX3 U700 ( .A(n860), .Y(n917) );
  INVX1 U701 ( .A(n269), .Y(n922) );
  INVX1 U702 ( .A(n272), .Y(n926) );
  INVX1 U703 ( .A(n268), .Y(n920) );
  INVX1 U704 ( .A(n841), .Y(n907) );
  CLKINVX3 U705 ( .A(b[4]), .Y(n925) );
  CLKINVX3 U706 ( .A(n857), .Y(n923) );
  INVX1 U707 ( .A(b[0]), .Y(n877) );
  INVX1 U708 ( .A(n273), .Y(n928) );
  BUFX3 U709 ( .A(b[10]), .Y(n860) );
  INVX1 U710 ( .A(n844), .Y(n902) );
  INVX1 U711 ( .A(n274), .Y(n930) );
  INVX1 U712 ( .A(n847), .Y(n895) );
  CLKINVX3 U713 ( .A(n1037), .Y(n897) );
  INVX1 U714 ( .A(n870), .Y(n869) );
  INVX1 U715 ( .A(n843), .Y(n904) );
  CLKINVX3 U716 ( .A(n868), .Y(n130) );
  INVX1 U717 ( .A(n845), .Y(n901) );
  INVX1 U718 ( .A(n840), .Y(n909) );
  INVX1 U719 ( .A(n842), .Y(n906) );
  INVX1 U720 ( .A(n846), .Y(n899) );
  INVX1 U721 ( .A(n80), .Y(n880) );
  BUFX4 U722 ( .A(b[9]), .Y(n859) );
  BUFX3 U723 ( .A(b[6]), .Y(n857) );
  INVX1 U724 ( .A(n185), .Y(n888) );
  INVX1 U725 ( .A(n192), .Y(n894) );
  CLKINVX3 U726 ( .A(n856), .Y(n924) );
  CLKINVX3 U727 ( .A(n854), .Y(n929) );
  CLKINVX3 U728 ( .A(n855), .Y(n927) );
  INVX1 U729 ( .A(n858), .Y(n921) );
  CLKINVX2 U730 ( .A(n1054), .Y(n892) );
  INVX1 U731 ( .A(n853), .Y(n931) );
  INVX1 U732 ( .A(n849), .Y(n891) );
  BUFX3 U733 ( .A(n993), .Y(n845) );
  NOR2BX1 U734 ( .AN(n1020), .B(n1022), .Y(n993) );
  BUFX3 U735 ( .A(n997), .Y(n844) );
  NAND3BX1 U736 ( .AN(n1020), .B(n1022), .C(n1021), .Y(n997) );
  BUFX3 U737 ( .A(n1028), .Y(n847) );
  NAND3BX1 U738 ( .AN(n1090), .B(n1091), .C(n1092), .Y(n1028) );
  BUFX3 U739 ( .A(n962), .Y(n842) );
  NOR2BX1 U740 ( .AN(n989), .B(n991), .Y(n962) );
  INVX1 U741 ( .A(n850), .Y(n890) );
  BUFX3 U742 ( .A(n1026), .Y(n846) );
  NOR2X1 U743 ( .A(n1090), .B(n1092), .Y(n1026) );
  BUFX3 U744 ( .A(n966), .Y(n841) );
  NAND3BX1 U745 ( .AN(n989), .B(n991), .C(n990), .Y(n966) );
  BUFX3 U746 ( .A(n995), .Y(n843) );
  NOR2X1 U747 ( .A(n1020), .B(n1021), .Y(n995) );
  INVX1 U748 ( .A(n873), .Y(n870) );
  INVX1 U749 ( .A(n863), .Y(n903) );
  INVX1 U750 ( .A(n864), .Y(n898) );
  INVX1 U751 ( .A(n848), .Y(n893) );
  BUFX3 U752 ( .A(n964), .Y(n840) );
  NOR2X1 U753 ( .A(n989), .B(n990), .Y(n964) );
  INVX1 U754 ( .A(n871), .Y(n868) );
  INVX1 U755 ( .A(n872), .Y(n871) );
  INVX1 U756 ( .A(n862), .Y(n908) );
  INVX1 U757 ( .A(n839), .Y(n911) );
  INVX1 U758 ( .A(n838), .Y(n912) );
  BUFX3 U759 ( .A(b[5]), .Y(n856) );
  BUFX3 U760 ( .A(b[7]), .Y(n858) );
  BUFX3 U761 ( .A(b[3]), .Y(n855) );
  BUFX3 U762 ( .A(b[1]), .Y(n853) );
  BUFX3 U763 ( .A(b[2]), .Y(n854) );
  INVX1 U764 ( .A(n172), .Y(n889) );
  BUFX3 U765 ( .A(n708), .Y(n864) );
  INVX1 U766 ( .A(n152), .Y(n881) );
  INVX1 U767 ( .A(n165), .Y(n882) );
  BUFX3 U768 ( .A(n709), .Y(n863) );
  XNOR2X1 U769 ( .A(n1076), .B(n874), .Y(n317) );
  OAI21XL U770 ( .A0(n923), .A1(n886), .B0(n1080), .Y(n1079) );
  BUFX3 U771 ( .A(n710), .Y(n862) );
  XNOR2X1 U772 ( .A(n1082), .B(n874), .Y(n313) );
  BUFX3 U773 ( .A(n1050), .Y(n850) );
  NOR2BX1 U774 ( .AN(n1097), .B(n1098), .Y(n1050) );
  INVX1 U775 ( .A(n861), .Y(n913) );
  BUFX3 U776 ( .A(n1053), .Y(n849) );
  NAND3BX1 U777 ( .AN(n1097), .B(n1098), .C(n1099), .Y(n1053) );
  BUFX3 U778 ( .A(n1051), .Y(n848) );
  NOR2X1 U779 ( .A(n1097), .B(n1099), .Y(n1051) );
  INVX1 U780 ( .A(n866), .Y(n873) );
  BUFX3 U781 ( .A(n933), .Y(n839) );
  NOR2X1 U782 ( .A(n960), .B(n916), .Y(n933) );
  BUFX3 U783 ( .A(n936), .Y(n838) );
  CLKINVX3 U784 ( .A(n944), .Y(n914) );
  INVX1 U785 ( .A(n1085), .Y(n883) );
  INVX1 U786 ( .A(n865), .Y(n887) );
  INVX1 U787 ( .A(n866), .Y(n872) );
  AOI22X1 U788 ( .A0(n852), .A1(n853), .B0(n851), .B1(n878), .Y(n1074) );
  BUFX3 U789 ( .A(a[14]), .Y(n865) );
  XNOR2X1 U790 ( .A(n1083), .B(n874), .Y(n312) );
  BUFX3 U791 ( .A(a[2]), .Y(n861) );
  OAI21XL U792 ( .A0(n925), .A1(n886), .B0(n1102), .Y(n1101) );
  NAND2X1 U793 ( .A(n851), .B(n855), .Y(n1102) );
  INVX1 U794 ( .A(a[1]), .Y(n915) );
  OAI21XL U795 ( .A0(n925), .A1(n884), .B0(n1078), .Y(n1077) );
  NAND2X1 U796 ( .A(n852), .B(n856), .Y(n1078) );
  XNOR2X1 U797 ( .A(n1100), .B(n874), .Y(n165) );
  INVX1 U798 ( .A(n867), .Y(n866) );
  INVX1 U799 ( .A(n79), .Y(n867) );
  XNOR2X1 U800 ( .A(n1084), .B(n874), .Y(n311) );
  INVX1 U801 ( .A(n1081), .Y(n885) );
  NAND2X1 U802 ( .A(n878), .B(n852), .Y(n1072) );
  NAND2X1 U803 ( .A(n851), .B(n856), .Y(n1080) );
  CLKINVX3 U804 ( .A(n875), .Y(n874) );
  INVX1 U805 ( .A(n706), .Y(n875) );
  INVX1 U806 ( .A(a[0]), .Y(n916) );
  INVX1 U807 ( .A(n851), .Y(n884) );
  INVX1 U808 ( .A(n132), .Y(n876) );
  INVX1 U809 ( .A(n852), .Y(n886) );
  BUFX3 U810 ( .A(n1075), .Y(n851) );
  NOR2X1 U811 ( .A(n852), .B(n1103), .Y(n1075) );
  BUFX3 U812 ( .A(n1073), .Y(n852) );
  XOR2X1 U813 ( .A(a[15]), .B(n865), .Y(n1073) );
  XNOR2X1 U814 ( .A(n74), .B(n36), .Y(n932) );
  XOR2X1 U815 ( .A(n913), .B(n934), .Y(n380) );
  XOR2X1 U816 ( .A(n935), .B(n861), .Y(n379) );
  OAI221XL U817 ( .A0(n879), .A1(n838), .B0(n930), .B1(n937), .C0(n938), .Y(
        n935) );
  AOI22X1 U818 ( .A0(n839), .A1(n854), .B0(n914), .B1(n853), .Y(n938) );
  XOR2X1 U819 ( .A(n939), .B(n861), .Y(n378) );
  OAI221XL U820 ( .A0(n931), .A1(n838), .B0(n937), .B1(n928), .C0(n940), .Y(
        n939) );
  AOI22X1 U821 ( .A0(n839), .A1(n855), .B0(n914), .B1(n854), .Y(n940) );
  XOR2X1 U822 ( .A(n941), .B(n861), .Y(n377) );
  OAI221XL U823 ( .A0(n929), .A1(n838), .B0(n926), .B1(n937), .C0(n942), .Y(
        n941) );
  XOR2X1 U824 ( .A(n943), .B(n861), .Y(n376) );
  OAI221XL U825 ( .A0(n925), .A1(n944), .B0(n927), .B1(n838), .C0(n945), .Y(
        n943) );
  XOR2X1 U826 ( .A(n946), .B(n861), .Y(n375) );
  OAI221XL U827 ( .A0(n925), .A1(n838), .B0(n923), .B1(n911), .C0(n947), .Y(
        n946) );
  XOR2X1 U828 ( .A(n948), .B(n861), .Y(n374) );
  OAI221XL U829 ( .A0(n924), .A1(n838), .B0(n922), .B1(n937), .C0(n949), .Y(
        n948) );
  AOI22X1 U830 ( .A0(n839), .A1(n858), .B0(n914), .B1(n857), .Y(n949) );
  XOR2X1 U831 ( .A(n950), .B(n861), .Y(n373) );
  OAI221XL U832 ( .A0(n923), .A1(n838), .B0(n937), .B1(n920), .C0(n951), .Y(
        n950) );
  AOI22X1 U833 ( .A0(n839), .A1(b[8]), .B0(n914), .B1(n858), .Y(n951) );
  XOR2X1 U834 ( .A(n952), .B(n861), .Y(n372) );
  OAI221XL U835 ( .A0(n921), .A1(n838), .B0(n937), .B1(n919), .C0(n953), .Y(
        n952) );
  AOI22X1 U836 ( .A0(n839), .A1(n859), .B0(n914), .B1(n859), .Y(n953) );
  XOR2X1 U837 ( .A(n954), .B(n861), .Y(n371) );
  OAI221XL U838 ( .A0(n917), .A1(n838), .B0(n918), .B1(n937), .C0(n955), .Y(
        n954) );
  AOI22X1 U839 ( .A0(n839), .A1(b[30]), .B0(n914), .B1(n859), .Y(n955) );
  XOR2X1 U840 ( .A(n913), .B(n956), .Y(n370) );
  AOI221X1 U841 ( .A0(n265), .A1(n910), .B0(n912), .B1(n859), .C0(n957), .Y(
        n956) );
  AOI21X1 U842 ( .A0(n944), .A1(n911), .B0(n917), .Y(n957) );
  XOR2X1 U843 ( .A(n861), .B(n958), .Y(n369) );
  AOI221X1 U844 ( .A0(n910), .A1(n860), .B0(n839), .B1(b[29]), .C0(n959), .Y(
        n958) );
  AOI21X1 U845 ( .A0(n838), .A1(n944), .B0(n917), .Y(n959) );
  NAND2X1 U846 ( .A(a[1]), .B(n916), .Y(n944) );
  NAND3X1 U847 ( .A(n916), .B(n915), .C(n960), .Y(n936) );
  XOR2X1 U848 ( .A(n915), .B(n913), .Y(n960) );
  XOR2X1 U849 ( .A(n908), .B(n961), .Y(n368) );
  XOR2X1 U850 ( .A(n908), .B(n963), .Y(n367) );
  XOR2X1 U851 ( .A(n965), .B(n862), .Y(n366) );
  OAI221XL U852 ( .A0(n877), .A1(n841), .B0(n930), .B1(n967), .C0(n968), .Y(
        n965) );
  AOI22X1 U853 ( .A0(n842), .A1(n854), .B0(n840), .B1(n853), .Y(n968) );
  XOR2X1 U854 ( .A(n969), .B(n862), .Y(n365) );
  OAI221XL U855 ( .A0(n931), .A1(n841), .B0(n928), .B1(n967), .C0(n970), .Y(
        n969) );
  AOI22X1 U856 ( .A0(n842), .A1(n855), .B0(n840), .B1(n854), .Y(n970) );
  XOR2X1 U857 ( .A(n971), .B(n862), .Y(n364) );
  OAI221XL U858 ( .A0(n929), .A1(n841), .B0(n926), .B1(n967), .C0(n972), .Y(
        n971) );
  XOR2X1 U859 ( .A(n973), .B(n862), .Y(n363) );
  OAI221XL U860 ( .A0(n925), .A1(n909), .B0(n927), .B1(n841), .C0(n974), .Y(
        n973) );
  XOR2X1 U861 ( .A(n975), .B(n862), .Y(n362) );
  OAI221XL U862 ( .A0(n925), .A1(n841), .B0(n923), .B1(n906), .C0(n976), .Y(
        n975) );
  XOR2X1 U863 ( .A(n977), .B(n862), .Y(n361) );
  OAI221XL U864 ( .A0(n924), .A1(n841), .B0(n922), .B1(n967), .C0(n978), .Y(
        n977) );
  AOI22X1 U865 ( .A0(n842), .A1(n858), .B0(n840), .B1(n857), .Y(n978) );
  XOR2X1 U866 ( .A(n979), .B(n862), .Y(n360) );
  OAI221XL U867 ( .A0(n923), .A1(n841), .B0(n920), .B1(n967), .C0(n980), .Y(
        n979) );
  AOI22X1 U868 ( .A0(n842), .A1(b[8]), .B0(n840), .B1(n858), .Y(n980) );
  XOR2X1 U869 ( .A(n981), .B(n862), .Y(n359) );
  OAI221XL U870 ( .A0(n921), .A1(n841), .B0(n919), .B1(n967), .C0(n982), .Y(
        n981) );
  AOI22X1 U871 ( .A0(n842), .A1(n859), .B0(n840), .B1(b[8]), .Y(n982) );
  XOR2X1 U872 ( .A(n983), .B(n862), .Y(n358) );
  OAI221XL U873 ( .A0(n917), .A1(n841), .B0(n918), .B1(n967), .C0(n984), .Y(
        n983) );
  AOI22X1 U874 ( .A0(n842), .A1(n860), .B0(n840), .B1(n859), .Y(n984) );
  XOR2X1 U875 ( .A(n908), .B(n985), .Y(n357) );
  AOI221X1 U876 ( .A0(n905), .A1(n265), .B0(n907), .B1(n859), .C0(n986), .Y(
        n985) );
  AOI21X1 U877 ( .A0(n909), .A1(n906), .B0(n917), .Y(n986) );
  XOR2X1 U878 ( .A(n862), .B(n987), .Y(n356) );
  AOI21X1 U879 ( .A0(n841), .A1(n909), .B0(n917), .Y(n988) );
  XNOR2X1 U880 ( .A(a[3]), .B(a[4]), .Y(n990) );
  XOR2X1 U881 ( .A(a[4]), .B(n862), .Y(n991) );
  XOR2X1 U882 ( .A(a[3]), .B(n861), .Y(n989) );
  XOR2X1 U883 ( .A(n903), .B(n992), .Y(n355) );
  XOR2X1 U884 ( .A(n903), .B(n994), .Y(n354) );
  XOR2X1 U885 ( .A(n996), .B(n863), .Y(n353) );
  OAI221XL U886 ( .A0(n877), .A1(n844), .B0(n930), .B1(n998), .C0(n999), .Y(
        n996) );
  AOI22X1 U887 ( .A0(n845), .A1(n854), .B0(n843), .B1(n853), .Y(n999) );
  XOR2X1 U888 ( .A(n1000), .B(n863), .Y(n352) );
  OAI221XL U889 ( .A0(n931), .A1(n844), .B0(n928), .B1(n998), .C0(n1001), .Y(
        n1000) );
  AOI22X1 U890 ( .A0(n845), .A1(n855), .B0(n843), .B1(n854), .Y(n1001) );
  XOR2X1 U891 ( .A(n1002), .B(n863), .Y(n351) );
  OAI221XL U892 ( .A0(n929), .A1(n844), .B0(n926), .B1(n998), .C0(n1003), .Y(
        n1002) );
  XOR2X1 U893 ( .A(n1004), .B(n863), .Y(n350) );
  OAI221XL U894 ( .A0(n925), .A1(n904), .B0(n927), .B1(n844), .C0(n1005), .Y(
        n1004) );
  XOR2X1 U895 ( .A(n1006), .B(n863), .Y(n349) );
  OAI221XL U896 ( .A0(n925), .A1(n844), .B0(n923), .B1(n901), .C0(n1007), .Y(
        n1006) );
  XOR2X1 U897 ( .A(n1008), .B(n863), .Y(n348) );
  OAI221XL U898 ( .A0(n924), .A1(n844), .B0(n922), .B1(n998), .C0(n1009), .Y(
        n1008) );
  AOI22X1 U899 ( .A0(n845), .A1(n858), .B0(n843), .B1(n857), .Y(n1009) );
  XOR2X1 U900 ( .A(n1010), .B(n863), .Y(n347) );
  OAI221XL U901 ( .A0(n923), .A1(n844), .B0(n920), .B1(n998), .C0(n1011), .Y(
        n1010) );
  AOI22X1 U902 ( .A0(n845), .A1(b[9]), .B0(n843), .B1(n858), .Y(n1011) );
  XOR2X1 U903 ( .A(n1012), .B(n863), .Y(n346) );
  OAI221XL U904 ( .A0(n921), .A1(n844), .B0(n919), .B1(n998), .C0(n1013), .Y(
        n1012) );
  AOI22X1 U905 ( .A0(n845), .A1(n859), .B0(n843), .B1(b[9]), .Y(n1013) );
  XOR2X1 U906 ( .A(n1014), .B(n863), .Y(n345) );
  OAI221XL U907 ( .A0(n917), .A1(n844), .B0(n918), .B1(n998), .C0(n1015), .Y(
        n1014) );
  AOI22X1 U908 ( .A0(n845), .A1(n860), .B0(n843), .B1(n859), .Y(n1015) );
  XOR2X1 U909 ( .A(n903), .B(n1016), .Y(n344) );
  AOI221X1 U910 ( .A0(n900), .A1(n265), .B0(n902), .B1(n859), .C0(n1017), .Y(
        n1016) );
  AOI21X1 U911 ( .A0(n904), .A1(n901), .B0(n917), .Y(n1017) );
  XOR2X1 U912 ( .A(n863), .B(n1018), .Y(n343) );
  AOI221X1 U913 ( .A0(n900), .A1(n860), .B0(n845), .B1(n860), .C0(n1019), .Y(
        n1018) );
  AOI21X1 U914 ( .A0(n844), .A1(n904), .B0(n917), .Y(n1019) );
  XNOR2X1 U915 ( .A(a[6]), .B(a[7]), .Y(n1021) );
  XOR2X1 U916 ( .A(a[7]), .B(n863), .Y(n1022) );
  XOR2X1 U917 ( .A(a[6]), .B(n862), .Y(n1020) );
  XOR2X1 U918 ( .A(n898), .B(n1023), .Y(n342) );
  XOR2X1 U919 ( .A(n898), .B(n1025), .Y(n341) );
  XOR2X1 U920 ( .A(n1027), .B(n864), .Y(n340) );
  OAI221XL U921 ( .A0(n877), .A1(n847), .B0(n929), .B1(n896), .C0(n1029), .Y(
        n1027) );
  AOI22X1 U922 ( .A0(n846), .A1(n853), .B0(n897), .B1(n274), .Y(n1029) );
  XOR2X1 U923 ( .A(n1030), .B(n864), .Y(n339) );
  OAI221XL U924 ( .A0(n931), .A1(n847), .B0(n927), .B1(n896), .C0(n1031), .Y(
        n1030) );
  AOI22X1 U925 ( .A0(n846), .A1(n854), .B0(n897), .B1(n273), .Y(n1031) );
  XOR2X1 U926 ( .A(n1032), .B(n864), .Y(n338) );
  OAI221XL U927 ( .A0(n927), .A1(n847), .B0(n924), .B1(n896), .C0(n1033), .Y(
        n1032) );
  XOR2X1 U928 ( .A(n1034), .B(n864), .Y(n337) );
  OAI221XL U929 ( .A0(n925), .A1(n847), .B0(n923), .B1(n896), .C0(n1035), .Y(
        n1034) );
  AOI22X1 U930 ( .A0(n846), .A1(n856), .B0(n897), .B1(n270), .Y(n1035) );
  XOR2X1 U931 ( .A(n1036), .B(n864), .Y(n336) );
  OAI221XL U932 ( .A0(n924), .A1(n847), .B0(n922), .B1(n1037), .C0(n1038), .Y(
        n1036) );
  XOR2X1 U933 ( .A(n1039), .B(n864), .Y(n335) );
  OAI221XL U934 ( .A0(n923), .A1(n847), .B0(n920), .B1(n1037), .C0(n1040), .Y(
        n1039) );
  XOR2X1 U935 ( .A(n1041), .B(n864), .Y(n334) );
  OAI221XL U936 ( .A0(n921), .A1(n847), .B0(n919), .B1(n1037), .C0(n1042), .Y(
        n1041) );
  XOR2X1 U937 ( .A(n1043), .B(n864), .Y(n333) );
  OAI221XL U938 ( .A0(n917), .A1(n847), .B0(n918), .B1(n1037), .C0(n1044), .Y(
        n1043) );
  XOR2X1 U939 ( .A(n898), .B(n1045), .Y(n332) );
  AOI221X1 U940 ( .A0(n897), .A1(n265), .B0(n895), .B1(n859), .C0(n1046), .Y(
        n1045) );
  XOR2X1 U941 ( .A(n864), .B(n1047), .Y(n331) );
  AOI21X1 U942 ( .A0(n847), .A1(n899), .B0(n917), .Y(n1048) );
  XOR2X1 U943 ( .A(n887), .B(n1049), .Y(n329) );
  AOI222X1 U944 ( .A0(n892), .A1(n275), .B0(n850), .B1(n853), .C0(n848), .C1(
        n878), .Y(n1049) );
  XOR2X1 U945 ( .A(n1052), .B(n865), .Y(n328) );
  OAI221XL U946 ( .A0(n931), .A1(n849), .B0(n928), .B1(n1054), .C0(n1055), .Y(
        n1052) );
  AOI22X1 U947 ( .A0(n848), .A1(n854), .B0(n850), .B1(n855), .Y(n1055) );
  XOR2X1 U948 ( .A(n1056), .B(n865), .Y(n327) );
  OAI221XL U949 ( .A0(n925), .A1(n893), .B0(n927), .B1(n849), .C0(n1057), .Y(
        n1056) );
  AOI22X1 U950 ( .A0(n850), .A1(n856), .B0(n892), .B1(n271), .Y(n1057) );
  XOR2X1 U951 ( .A(n1058), .B(n865), .Y(n326) );
  OAI221XL U952 ( .A0(n925), .A1(n849), .B0(n923), .B1(n890), .C0(n1059), .Y(
        n1058) );
  AOI22X1 U953 ( .A0(n848), .A1(n856), .B0(n892), .B1(n270), .Y(n1059) );
  XOR2X1 U954 ( .A(n1060), .B(n865), .Y(n325) );
  OAI221XL U955 ( .A0(n924), .A1(n849), .B0(n922), .B1(n1054), .C0(n1061), .Y(
        n1060) );
  AOI22X1 U956 ( .A0(n850), .A1(n858), .B0(n848), .B1(n857), .Y(n1061) );
  XOR2X1 U957 ( .A(n1062), .B(n865), .Y(n324) );
  OAI221XL U958 ( .A0(n923), .A1(n849), .B0(n920), .B1(n1054), .C0(n1063), .Y(
        n1062) );
  AOI22X1 U959 ( .A0(n850), .A1(b[9]), .B0(n848), .B1(n858), .Y(n1063) );
  XOR2X1 U960 ( .A(n1064), .B(n865), .Y(n323) );
  OAI221XL U961 ( .A0(n921), .A1(n849), .B0(n919), .B1(n1054), .C0(n1065), .Y(
        n1064) );
  AOI22X1 U962 ( .A0(n850), .A1(n859), .B0(n848), .B1(n860), .Y(n1065) );
  XOR2X1 U963 ( .A(n1066), .B(n865), .Y(n322) );
  OAI221XL U964 ( .A0(n917), .A1(n849), .B0(n918), .B1(n1054), .C0(n1067), .Y(
        n1066) );
  AOI22X1 U965 ( .A0(n850), .A1(n860), .B0(n848), .B1(n859), .Y(n1067) );
  XOR2X1 U966 ( .A(n887), .B(n1068), .Y(n321) );
  AOI221X1 U967 ( .A0(n892), .A1(n265), .B0(n891), .B1(n859), .C0(n1069), .Y(
        n1068) );
  AOI21X1 U968 ( .A0(n893), .A1(n890), .B0(n917), .Y(n1069) );
  XOR2X1 U969 ( .A(n865), .B(n1070), .Y(n320) );
  AOI221X1 U970 ( .A0(n892), .A1(n860), .B0(n850), .B1(n859), .C0(n1071), .Y(
        n1070) );
  AOI21X1 U971 ( .A0(n849), .A1(n893), .B0(n917), .Y(n1071) );
  XOR2X1 U972 ( .A(n869), .B(n1072), .Y(n319) );
  XOR2X1 U973 ( .A(n869), .B(n1074), .Y(n318) );
  AOI22X1 U974 ( .A0(n851), .A1(n854), .B0(n852), .B1(n855), .Y(n1076) );
  XOR2X1 U975 ( .A(n1077), .B(n874), .Y(n316) );
  XOR2X1 U976 ( .A(n1079), .B(n874), .Y(n315) );
  XOR2X1 U977 ( .A(n885), .B(n874), .Y(n314) );
  AOI22X1 U978 ( .A0(n852), .A1(n858), .B0(n851), .B1(n857), .Y(n1081) );
  AOI22X1 U979 ( .A0(n852), .A1(n860), .B0(n851), .B1(n858), .Y(n1082) );
  AOI22X1 U980 ( .A0(n852), .A1(n859), .B0(n851), .B1(n860), .Y(n1083) );
  AOI22X1 U981 ( .A0(n852), .A1(n860), .B0(n851), .B1(n859), .Y(n1084) );
  XOR2X1 U982 ( .A(n875), .B(n883), .Y(n310) );
  XOR2X1 U983 ( .A(n874), .B(n883), .Y(n309) );
  AOI21X1 U984 ( .A0(n884), .A1(n886), .B0(n917), .Y(n1085) );
  XOR2X1 U985 ( .A(n865), .B(n1086), .Y(n200) );
  NAND2X1 U986 ( .A(n1086), .B(n887), .Y(n199) );
  XOR2X1 U987 ( .A(n865), .B(n1087), .Y(n1086) );
  AOI22X1 U988 ( .A0(n892), .A1(n878), .B0(n850), .B1(b[0]), .Y(n1087) );
  XOR2X1 U989 ( .A(n1088), .B(n864), .Y(n192) );
  OAI221XL U990 ( .A0(n929), .A1(n847), .B0(n925), .B1(n896), .C0(n1089), .Y(
        n1088) );
  AOI22X1 U991 ( .A0(n846), .A1(n855), .B0(n897), .B1(n272), .Y(n1089) );
  NAND2X1 U992 ( .A(n1090), .B(n1091), .Y(n1037) );
  XNOR2X1 U993 ( .A(a[10]), .B(a[9]), .Y(n1092) );
  XOR2X1 U994 ( .A(a[10]), .B(n864), .Y(n1091) );
  XOR2X1 U995 ( .A(a[9]), .B(n863), .Y(n1090) );
  XOR2X1 U996 ( .A(n1093), .B(n865), .Y(n185) );
  OAI221XL U997 ( .A0(n877), .A1(n849), .B0(n930), .B1(n1054), .C0(n1094), .Y(
        n1093) );
  AOI22X1 U998 ( .A0(n850), .A1(n854), .B0(n848), .B1(n853), .Y(n1094) );
  XOR2X1 U999 ( .A(n1095), .B(n865), .Y(n172) );
  OAI221XL U1000 ( .A0(n925), .A1(n890), .B0(n929), .B1(n849), .C0(n1096), .Y(
        n1095) );
  AOI22X1 U1001 ( .A0(n848), .A1(n855), .B0(n892), .B1(n272), .Y(n1096) );
  XNOR2X1 U1002 ( .A(a[12]), .B(a[13]), .Y(n1099) );
  XOR2X1 U1003 ( .A(a[13]), .B(n865), .Y(n1098) );
  XOR2X1 U1004 ( .A(a[12]), .B(n864), .Y(n1097) );
  AOI22X1 U1005 ( .A0(n852), .A1(n854), .B0(n851), .B1(n853), .Y(n1100) );
  XOR2X1 U1006 ( .A(n1101), .B(n874), .Y(n152) );
  XNOR2X1 U1007 ( .A(a[15]), .B(a[16]), .Y(n1103) );
endmodule


module Equation_Implementation_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  ADDFX2 U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFX2 U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFX2 U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFX2 U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFX2 U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  INVX1 U1 ( .A(carry[7]), .Y(DIFF[7]) );
  XNOR2X2 U2 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
  INVX1 U3 ( .A(B[3]), .Y(n5) );
  INVX1 U4 ( .A(B[2]), .Y(n6) );
  INVX1 U5 ( .A(B[0]), .Y(n8) );
  INVX1 U6 ( .A(B[1]), .Y(n7) );
  OR2X2 U7 ( .A(A[0]), .B(n8), .Y(carry[1]) );
  INVX1 U8 ( .A(B[5]), .Y(n3) );
  INVX1 U9 ( .A(B[6]), .Y(n2) );
  INVX1 U10 ( .A(B[4]), .Y(n4) );
endmodule


module Equation_Implementation_DW_mult_uns_3 ( a, b, product );
  input [11:0] a;
  input [9:0] b;
  output [21:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, \a[0] , \a[1] , n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105;
  assign product[3] = \a[0] ;
  assign \a[0]  = a[0];
  assign product[4] = \a[1] ;
  assign \a[1]  = a[1];

  ADDFX2 U3 ( .A(n103), .B(a[9]), .CI(n3), .CO(n2), .S(product[20]) );
  ADDFX2 U4 ( .A(n102), .B(a[8]), .CI(n4), .CO(n3), .S(product[19]) );
  ADDFX2 U5 ( .A(n101), .B(a[7]), .CI(n5), .CO(n4), .S(product[18]) );
  ADDFX2 U6 ( .A(n100), .B(n27), .CI(n6), .CO(n5), .S(product[17]) );
  ADDFX2 U7 ( .A(n28), .B(n29), .CI(n7), .CO(n6), .S(product[16]) );
  ADDFX2 U8 ( .A(n30), .B(n31), .CI(n8), .CO(n7), .S(product[15]) );
  ADDFX2 U9 ( .A(n32), .B(n33), .CI(n9), .CO(n8), .S(product[14]) );
  ADDFX2 U10 ( .A(n34), .B(n35), .CI(n10), .CO(n9), .S(product[13]) );
  ADDFX2 U11 ( .A(n36), .B(n37), .CI(n11), .CO(n10), .S(product[12]) );
  ADDFX2 U12 ( .A(n38), .B(n39), .CI(n12), .CO(n11), .S(product[11]) );
  ADDFX2 U13 ( .A(n40), .B(n98), .CI(n13), .CO(n12), .S(product[10]) );
  ADDFX2 U14 ( .A(n97), .B(a[6]), .CI(n14), .CO(n13), .S(product[9]) );
  ADDFX2 U15 ( .A(n96), .B(a[5]), .CI(n15), .CO(n14), .S(product[8]) );
  ADDFX2 U16 ( .A(n95), .B(a[4]), .CI(n16), .CO(n15), .S(product[7]) );
  ADDFX2 U17 ( .A(n94), .B(a[3]), .CI(n17), .CO(n16), .S(product[6]) );
  ADDHXL U25 ( .A(a[6]), .B(n104), .CO(n27), .S(n28) );
  ADDHXL U26 ( .A(a[5]), .B(n103), .CO(n29), .S(n30) );
  ADDFX2 U27 ( .A(a[4]), .B(a[11]), .CI(n102), .CO(n31), .S(n32) );
  ADDFX2 U28 ( .A(a[3]), .B(a[10]), .CI(n101), .CO(n33), .S(n34) );
  ADDFX2 U29 ( .A(a[2]), .B(a[9]), .CI(n100), .CO(n35), .S(n36) );
  ADDFX2 U30 ( .A(\a[1] ), .B(a[8]), .CI(n99), .CO(n37), .S(n38) );
  ADDHXL U31 ( .A(a[7]), .B(\a[0] ), .CO(n39), .S(n40) );
  INVXL U48 ( .A(\a[1] ), .Y(n94) );
  INVX1 U49 ( .A(a[3]), .Y(n96) );
  INVX1 U50 ( .A(a[4]), .Y(n97) );
  INVX1 U51 ( .A(a[5]), .Y(n98) );
  INVX1 U52 ( .A(a[2]), .Y(n95) );
  INVX1 U53 ( .A(a[6]), .Y(n99) );
  INVX1 U54 ( .A(a[7]), .Y(n100) );
  INVX1 U55 ( .A(a[10]), .Y(n103) );
  INVX1 U56 ( .A(a[8]), .Y(n101) );
  INVX1 U57 ( .A(a[9]), .Y(n102) );
  INVX1 U58 ( .A(a[11]), .Y(n104) );
  XOR2X1 U59 ( .A(a[2]), .B(\a[0] ), .Y(product[5]) );
  XOR2X1 U60 ( .A(n103), .B(n105), .Y(product[21]) );
  XOR2X1 U61 ( .A(n2), .B(a[11]), .Y(n105) );
  NAND2X1 U62 ( .A(\a[0] ), .B(n95), .Y(n17) );
endmodule


module Equation_Implementation_DW_mult_uns_2 ( a, b, product );
  input [12:0] a;
  input [9:0] b;
  output [22:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, \a[1] , \a[2] , n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106;
  assign product[4] = \a[1] ;
  assign \a[1]  = a[1];
  assign product[5] = \a[2] ;
  assign \a[2]  = a[2];

  ADDFX2 U3 ( .A(n96), .B(a[10]), .CI(n3), .CO(n2), .S(product[21]) );
  ADDFX2 U4 ( .A(n97), .B(a[9]), .CI(n4), .CO(n3), .S(product[20]) );
  ADDFX2 U5 ( .A(n98), .B(a[8]), .CI(n5), .CO(n4), .S(product[19]) );
  ADDFX2 U6 ( .A(n99), .B(n27), .CI(n6), .CO(n5), .S(product[18]) );
  ADDFX2 U7 ( .A(n28), .B(n29), .CI(n7), .CO(n6), .S(product[17]) );
  ADDFX2 U8 ( .A(n30), .B(n31), .CI(n8), .CO(n7), .S(product[16]) );
  ADDFX2 U9 ( .A(n32), .B(n33), .CI(n9), .CO(n8), .S(product[15]) );
  ADDFX2 U10 ( .A(n34), .B(n35), .CI(n10), .CO(n9), .S(product[14]) );
  ADDFX2 U11 ( .A(n36), .B(n37), .CI(n11), .CO(n10), .S(product[13]) );
  ADDFX2 U12 ( .A(n38), .B(n39), .CI(n12), .CO(n11), .S(product[12]) );
  ADDFX2 U13 ( .A(n40), .B(n101), .CI(n13), .CO(n12), .S(product[11]) );
  ADDFX2 U14 ( .A(n102), .B(a[7]), .CI(n14), .CO(n13), .S(product[10]) );
  ADDFX2 U15 ( .A(n103), .B(a[6]), .CI(n15), .CO(n14), .S(product[9]) );
  ADDFX2 U16 ( .A(n104), .B(a[5]), .CI(n16), .CO(n15), .S(product[8]) );
  ADDFX2 U17 ( .A(n105), .B(a[4]), .CI(n17), .CO(n16), .S(product[7]) );
  ADDHXL U25 ( .A(a[7]), .B(n95), .CO(n27), .S(n28) );
  ADDHXL U26 ( .A(a[6]), .B(n96), .CO(n29), .S(n30) );
  ADDFX2 U27 ( .A(a[5]), .B(a[12]), .CI(n97), .CO(n31), .S(n32) );
  ADDFX2 U28 ( .A(a[4]), .B(a[11]), .CI(n98), .CO(n33), .S(n34) );
  ADDFX2 U29 ( .A(a[3]), .B(a[10]), .CI(n99), .CO(n35), .S(n36) );
  ADDFX2 U30 ( .A(\a[2] ), .B(a[9]), .CI(n100), .CO(n37), .S(n38) );
  ADDHXL U31 ( .A(a[8]), .B(\a[1] ), .CO(n39), .S(n40) );
  XOR2XL U48 ( .A(n2), .B(a[12]), .Y(n106) );
  INVX1 U49 ( .A(\a[2] ), .Y(n105) );
  INVXL U50 ( .A(a[4]), .Y(n103) );
  INVXL U51 ( .A(a[5]), .Y(n102) );
  INVXL U52 ( .A(a[6]), .Y(n101) );
  INVXL U53 ( .A(a[3]), .Y(n104) );
  INVXL U54 ( .A(a[7]), .Y(n100) );
  INVXL U55 ( .A(a[9]), .Y(n98) );
  INVXL U56 ( .A(a[8]), .Y(n99) );
  INVX1 U57 ( .A(a[11]), .Y(n96) );
  INVXL U58 ( .A(a[10]), .Y(n97) );
  INVXL U59 ( .A(a[12]), .Y(n95) );
  XOR2X1 U60 ( .A(a[3]), .B(\a[1] ), .Y(product[6]) );
  XOR2X1 U61 ( .A(n96), .B(n106), .Y(product[22]) );
  NAND2X1 U62 ( .A(\a[1] ), .B(n104), .Y(n17) );
endmodule


module Equation_Implementation_DW_mult_uns_0 ( a, b, product );
  input [31:0] a;
  input [9:0] b;
  output [41:0] product;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n49, n51, n53, n55, n57, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n70, \a[1] , \a[2] , \product[22] , n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182;
  assign n70 = a[7];
  assign product[4] = \a[1] ;
  assign \a[1]  = a[1];
  assign product[5] = \a[2] ;
  assign \a[2]  = a[2];
  assign product[30] = \product[22] ;
  assign product[29] = \product[22] ;
  assign product[28] = \product[22] ;
  assign product[27] = \product[22] ;
  assign product[26] = \product[22] ;
  assign product[25] = \product[22] ;
  assign product[24] = \product[22] ;
  assign product[23] = \product[22] ;
  assign product[22] = \product[22] ;

  ADDFX2 U12 ( .A(n171), .B(n49), .CI(n12), .CO(n11), .S(product[21]) );
  ADDFX2 U13 ( .A(n172), .B(n51), .CI(n13), .CO(n12), .S(product[20]) );
  ADDFX2 U14 ( .A(n173), .B(n53), .CI(n14), .CO(n13), .S(product[19]) );
  ADDFX2 U15 ( .A(n174), .B(n55), .CI(n15), .CO(n14), .S(product[18]) );
  ADDFX2 U16 ( .A(n175), .B(n57), .CI(n16), .CO(n15), .S(product[17]) );
  ADDFX2 U17 ( .A(n176), .B(n59), .CI(n17), .CO(n16), .S(product[16]) );
  ADDFX2 U18 ( .A(n60), .B(n61), .CI(n18), .CO(n17), .S(product[15]) );
  ADDFX2 U19 ( .A(n62), .B(n63), .CI(n19), .CO(n18), .S(product[14]) );
  ADDFX2 U20 ( .A(n64), .B(n65), .CI(n20), .CO(n19), .S(product[13]) );
  ADDFX2 U21 ( .A(n66), .B(n67), .CI(n21), .CO(n20), .S(product[12]) );
  ADDFX2 U23 ( .A(n70), .B(n177), .CI(n23), .CO(n22), .S(product[10]) );
  ADDFX2 U24 ( .A(n178), .B(a[6]), .CI(n24), .CO(n23), .S(product[9]) );
  ADDFX2 U25 ( .A(n179), .B(a[5]), .CI(n25), .CO(n24), .S(product[8]) );
  ADDFX2 U26 ( .A(n180), .B(a[4]), .CI(n26), .CO(n25), .S(product[7]) );
  ADDFX2 U41 ( .A(a[10]), .B(a[17]), .CI(n171), .CO(n49) );
  ADDFX2 U42 ( .A(a[9]), .B(a[16]), .CI(n171), .CO(n51) );
  ADDFX2 U43 ( .A(a[8]), .B(a[15]), .CI(n171), .CO(n53) );
  ADDFX2 U44 ( .A(n70), .B(a[14]), .CI(n171), .CO(n55) );
  ADDFX2 U45 ( .A(a[6]), .B(a[13]), .CI(n171), .CO(n57) );
  ADDFX2 U46 ( .A(a[5]), .B(a[12]), .CI(n172), .CO(n59), .S(n60) );
  ADDFX2 U47 ( .A(a[4]), .B(a[11]), .CI(n173), .CO(n61), .S(n62) );
  ADDFX2 U48 ( .A(a[3]), .B(a[10]), .CI(n174), .CO(n63), .S(n64) );
  ADDFX2 U49 ( .A(\a[2] ), .B(a[9]), .CI(n175), .CO(n65), .S(n66) );
  ADDFX2 U50 ( .A(\a[1] ), .B(a[8]), .CI(n176), .CO(n67), .S(n68) );
  OR2XL U83 ( .A(a[3]), .B(n181), .Y(n26) );
  INVX8 U84 ( .A(n11), .Y(\product[22] ) );
  INVX1 U85 ( .A(a[5]), .Y(n177) );
  INVXL U86 ( .A(a[3]), .Y(n179) );
  INVX1 U87 ( .A(a[4]), .Y(n178) );
  INVX1 U88 ( .A(n70), .Y(n175) );
  INVX1 U89 ( .A(a[6]), .Y(n176) );
  INVX1 U90 ( .A(a[8]), .Y(n174) );
  INVX1 U91 ( .A(a[10]), .Y(n172) );
  INVX1 U92 ( .A(a[9]), .Y(n173) );
  CLKINVX3 U93 ( .A(a[27]), .Y(n171) );
  INVX1 U94 ( .A(\a[2] ), .Y(n180) );
  INVX1 U95 ( .A(\a[1] ), .Y(n181) );
  AND2X1 U96 ( .A(n68), .B(n22), .Y(n21) );
  XOR2X1 U97 ( .A(n68), .B(n22), .Y(product[11]) );
  XNOR2X1 U98 ( .A(n181), .B(a[3]), .Y(product[6]) );
  XOR2X1 U99 ( .A(n182), .B(a[28]), .Y(product[31]) );
  XNOR2X1 U100 ( .A(a[27]), .B(n11), .Y(n182) );
endmodule


module Equation_Implementation_DW_mult_uns_8 ( a, b, product );
  input [2:0] a;
  input [8:0] b;
  output [11:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n92, n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121;
  assign n12 = a[1];

  ADDFX2 U3 ( .A(n15), .B(n96), .CI(n3), .CO(n2), .S(product[10]) );
  ADDFX2 U4 ( .A(n16), .B(n24), .CI(n4), .CO(n3), .S(product[9]) );
  ADDFX2 U5 ( .A(n17), .B(n25), .CI(n5), .CO(n4), .S(product[8]) );
  ADDFX2 U6 ( .A(n18), .B(n26), .CI(n6), .CO(n5), .S(product[7]) );
  ADDFX2 U7 ( .A(n19), .B(n27), .CI(n7), .CO(n6), .S(product[6]) );
  ADDFX2 U8 ( .A(n20), .B(n28), .CI(n8), .CO(n7), .S(product[5]) );
  ADDFX2 U9 ( .A(n21), .B(n29), .CI(n9), .CO(n8), .S(product[4]) );
  ADDFX2 U10 ( .A(n22), .B(n30), .CI(n10), .CO(n9), .S(product[3]) );
  ADDFX2 U11 ( .A(n31), .B(n23), .CI(n11), .CO(n10), .S(product[2]) );
  ADDHXL U12 ( .A(n13), .B(n32), .CO(n11), .S(product[1]) );
  OR2X2 U68 ( .A(n98), .B(n108), .Y(n92) );
  CLKINVX3 U69 ( .A(a[0]), .Y(n98) );
  INVX1 U70 ( .A(n92), .Y(product[0]) );
  INVX1 U71 ( .A(b[8]), .Y(n100) );
  BUFX3 U72 ( .A(n112), .Y(n95) );
  NAND2X1 U73 ( .A(n96), .B(n98), .Y(n112) );
  INVX1 U74 ( .A(n96), .Y(n99) );
  INVX1 U75 ( .A(b[0]), .Y(n108) );
  INVX1 U76 ( .A(b[1]), .Y(n107) );
  INVX1 U77 ( .A(b[4]), .Y(n104) );
  INVX1 U78 ( .A(b[5]), .Y(n103) );
  INVX1 U79 ( .A(b[2]), .Y(n106) );
  INVX1 U80 ( .A(b[3]), .Y(n105) );
  INVX1 U81 ( .A(b[7]), .Y(n101) );
  INVX1 U82 ( .A(b[6]), .Y(n102) );
  BUFX3 U83 ( .A(n12), .Y(n96) );
  BUFX3 U84 ( .A(n121), .Y(n94) );
  XNOR2X1 U85 ( .A(a[2]), .B(n96), .Y(n121) );
  BUFX3 U86 ( .A(n111), .Y(n93) );
  NAND2X1 U87 ( .A(n94), .B(a[2]), .Y(n111) );
  XOR2X1 U88 ( .A(n109), .B(n110), .Y(product[11]) );
  XNOR2X1 U89 ( .A(n96), .B(n2), .Y(n110) );
  NAND2BX1 U90 ( .AN(n93), .B(b[8]), .Y(n109) );
  OAI22X1 U91 ( .A0(b[0]), .A1(n95), .B0(n113), .B1(n98), .Y(n32) );
  OAI22X1 U92 ( .A0(n113), .A1(n95), .B0(n114), .B1(n98), .Y(n31) );
  XNOR2X1 U93 ( .A(b[1]), .B(n96), .Y(n113) );
  OAI22X1 U94 ( .A0(n114), .A1(n95), .B0(n115), .B1(n98), .Y(n30) );
  XNOR2X1 U95 ( .A(b[2]), .B(n96), .Y(n114) );
  OAI22X1 U96 ( .A0(n115), .A1(n95), .B0(n116), .B1(n98), .Y(n29) );
  XNOR2X1 U97 ( .A(b[3]), .B(n96), .Y(n115) );
  OAI22X1 U98 ( .A0(n116), .A1(n95), .B0(n117), .B1(n98), .Y(n28) );
  XNOR2X1 U99 ( .A(b[4]), .B(n96), .Y(n116) );
  OAI22X1 U100 ( .A0(n117), .A1(n95), .B0(n118), .B1(n98), .Y(n27) );
  XNOR2X1 U101 ( .A(b[5]), .B(n96), .Y(n117) );
  OAI22X1 U102 ( .A0(n118), .A1(n95), .B0(n119), .B1(n98), .Y(n26) );
  XNOR2X1 U103 ( .A(b[6]), .B(n96), .Y(n118) );
  OAI22X1 U104 ( .A0(n119), .A1(n95), .B0(n120), .B1(n98), .Y(n25) );
  XNOR2X1 U105 ( .A(b[7]), .B(n96), .Y(n119) );
  OAI22X1 U106 ( .A0(n120), .A1(n95), .B0(n99), .B1(n98), .Y(n24) );
  XNOR2X1 U107 ( .A(b[8]), .B(n96), .Y(n120) );
  NOR2X1 U108 ( .A(n94), .B(n108), .Y(n23) );
  OAI22X1 U109 ( .A0(n93), .A1(n108), .B0(n94), .B1(n107), .Y(n22) );
  OAI22X1 U110 ( .A0(n93), .A1(n107), .B0(n94), .B1(n106), .Y(n21) );
  OAI22X1 U111 ( .A0(n93), .A1(n106), .B0(n94), .B1(n105), .Y(n20) );
  OAI22X1 U112 ( .A0(n93), .A1(n105), .B0(n94), .B1(n104), .Y(n19) );
  OAI22X1 U113 ( .A0(n93), .A1(n104), .B0(n94), .B1(n103), .Y(n18) );
  OAI22X1 U114 ( .A0(n93), .A1(n103), .B0(n94), .B1(n102), .Y(n17) );
  OAI22X1 U115 ( .A0(n93), .A1(n102), .B0(n94), .B1(n101), .Y(n16) );
  OAI22X1 U116 ( .A0(n93), .A1(n101), .B0(n94), .B1(n100), .Y(n15) );
  OAI21XL U117 ( .A0(b[0]), .A1(n99), .B0(n95), .Y(n13) );
endmodule


module Equation_Implementation_DW_div_uns_13 ( a, b, quotient, remainder, 
        divide_by_0 );
  input [31:0] a;
  input [9:0] b;
  output [31:0] quotient;
  output [9:0] remainder;
  output divide_by_0;
  wire   \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] , \u_div/SumTmp[1][3] ,
         \u_div/SumTmp[1][4] , \u_div/SumTmp[1][5] , \u_div/SumTmp[1][6] ,
         \u_div/SumTmp[1][7] , \u_div/SumTmp[1][8] , \u_div/SumTmp[1][9] ,
         \u_div/SumTmp[2][1] , \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] ,
         \u_div/SumTmp[2][4] , \u_div/SumTmp[2][5] , \u_div/SumTmp[2][6] ,
         \u_div/SumTmp[2][7] , \u_div/SumTmp[2][8] , \u_div/SumTmp[2][9] ,
         \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[3][5] , \u_div/SumTmp[3][6] ,
         \u_div/SumTmp[3][7] , \u_div/SumTmp[3][8] , \u_div/SumTmp[3][9] ,
         \u_div/SumTmp[4][0] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[4][5] ,
         \u_div/SumTmp[4][6] , \u_div/SumTmp[4][7] , \u_div/SumTmp[4][8] ,
         \u_div/SumTmp[4][9] , \u_div/SumTmp[5][0] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[5][5] , \u_div/SumTmp[5][6] , \u_div/SumTmp[5][7] ,
         \u_div/SumTmp[5][8] , \u_div/SumTmp[5][9] , \u_div/SumTmp[6][0] ,
         \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[6][5] , \u_div/SumTmp[6][6] ,
         \u_div/SumTmp[6][7] , \u_div/SumTmp[6][8] , \u_div/SumTmp[6][9] ,
         \u_div/SumTmp[7][0] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[7][5] ,
         \u_div/SumTmp[7][6] , \u_div/SumTmp[7][7] , \u_div/SumTmp[7][8] ,
         \u_div/SumTmp[7][9] , \u_div/SumTmp[8][0] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[8][5] , \u_div/SumTmp[8][6] , \u_div/SumTmp[8][7] ,
         \u_div/SumTmp[8][8] , \u_div/SumTmp[8][9] , \u_div/SumTmp[9][0] ,
         \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[9][5] , \u_div/SumTmp[9][6] ,
         \u_div/SumTmp[9][7] , \u_div/SumTmp[9][8] , \u_div/SumTmp[9][9] ,
         \u_div/SumTmp[10][0] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[10][5] ,
         \u_div/SumTmp[10][6] , \u_div/SumTmp[10][7] , \u_div/SumTmp[10][8] ,
         \u_div/SumTmp[10][9] , \u_div/SumTmp[11][0] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[11][5] , \u_div/SumTmp[11][6] , \u_div/SumTmp[11][7] ,
         \u_div/SumTmp[11][8] , \u_div/SumTmp[11][9] , \u_div/SumTmp[12][0] ,
         \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[12][4] , \u_div/SumTmp[12][5] , \u_div/SumTmp[12][6] ,
         \u_div/SumTmp[12][7] , \u_div/SumTmp[12][8] , \u_div/SumTmp[12][9] ,
         \u_div/SumTmp[13][0] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[13][5] ,
         \u_div/SumTmp[13][6] , \u_div/SumTmp[13][7] , \u_div/SumTmp[13][8] ,
         \u_div/SumTmp[13][9] , \u_div/SumTmp[14][0] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[14][5] , \u_div/SumTmp[14][6] , \u_div/SumTmp[14][7] ,
         \u_div/SumTmp[14][8] , \u_div/SumTmp[14][9] , \u_div/SumTmp[15][0] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[15][5] , \u_div/SumTmp[15][6] ,
         \u_div/SumTmp[15][7] , \u_div/SumTmp[15][8] , \u_div/SumTmp[15][9] ,
         \u_div/SumTmp[16][0] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[16][5] ,
         \u_div/SumTmp[16][6] , \u_div/SumTmp[16][7] , \u_div/SumTmp[16][8] ,
         \u_div/SumTmp[16][9] , \u_div/SumTmp[17][0] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[17][5] , \u_div/SumTmp[17][6] , \u_div/SumTmp[17][7] ,
         \u_div/SumTmp[17][8] , \u_div/SumTmp[17][9] , \u_div/SumTmp[18][0] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[18][5] , \u_div/SumTmp[18][6] ,
         \u_div/SumTmp[18][7] , \u_div/SumTmp[18][8] , \u_div/SumTmp[18][9] ,
         \u_div/SumTmp[19][0] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] , \u_div/SumTmp[19][5] ,
         \u_div/SumTmp[19][6] , \u_div/SumTmp[19][7] , \u_div/SumTmp[19][8] ,
         \u_div/SumTmp[19][9] , \u_div/SumTmp[20][0] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[20][5] , \u_div/SumTmp[20][6] , \u_div/SumTmp[20][7] ,
         \u_div/SumTmp[20][8] , \u_div/SumTmp[20][9] , \u_div/SumTmp[21][0] ,
         \u_div/SumTmp[21][1] , \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] ,
         \u_div/SumTmp[21][4] , \u_div/SumTmp[21][5] , \u_div/SumTmp[21][6] ,
         \u_div/SumTmp[21][7] , \u_div/SumTmp[21][8] , \u_div/SumTmp[21][9] ,
         \u_div/SumTmp[22][0] , \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] ,
         \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] , \u_div/SumTmp[22][5] ,
         \u_div/SumTmp[22][6] , \u_div/SumTmp[22][7] , \u_div/SumTmp[22][8] ,
         \u_div/SumTmp[22][9] , \u_div/SumTmp[23][0] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[23][5] , \u_div/SumTmp[23][6] , \u_div/SumTmp[23][7] ,
         \u_div/SumTmp[23][8] , \u_div/SumTmp[24][0] , \u_div/SumTmp[24][1] ,
         \u_div/SumTmp[24][2] , \u_div/SumTmp[24][3] , \u_div/SumTmp[24][4] ,
         \u_div/SumTmp[24][5] , \u_div/SumTmp[24][6] , \u_div/SumTmp[24][7] ,
         \u_div/SumTmp[25][0] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[25][5] ,
         \u_div/SumTmp[25][6] , \u_div/SumTmp[26][0] , \u_div/SumTmp[26][1] ,
         \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] , \u_div/SumTmp[26][4] ,
         \u_div/SumTmp[26][5] , \u_div/SumTmp[27][0] , \u_div/SumTmp[27][1] ,
         \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] , \u_div/SumTmp[27][4] ,
         \u_div/SumTmp[28][0] , \u_div/SumTmp[28][1] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][3] , \u_div/SumTmp[29][0] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[30][0] , \u_div/SumTmp[30][1] ,
         \u_div/SumTmp[31][0] , \u_div/CryTmp[0][2] , \u_div/CryTmp[0][3] ,
         \u_div/CryTmp[0][4] , \u_div/CryTmp[0][5] , \u_div/CryTmp[0][6] ,
         \u_div/CryTmp[0][7] , \u_div/CryTmp[0][8] , \u_div/CryTmp[0][9] ,
         \u_div/CryTmp[0][10] , \u_div/CryTmp[1][2] , \u_div/CryTmp[1][3] ,
         \u_div/CryTmp[1][4] , \u_div/CryTmp[1][5] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[1][7] , \u_div/CryTmp[1][8] , \u_div/CryTmp[1][9] ,
         \u_div/CryTmp[1][10] , \u_div/CryTmp[2][2] , \u_div/CryTmp[2][3] ,
         \u_div/CryTmp[2][4] , \u_div/CryTmp[2][5] , \u_div/CryTmp[2][6] ,
         \u_div/CryTmp[2][7] , \u_div/CryTmp[2][8] , \u_div/CryTmp[2][9] ,
         \u_div/CryTmp[2][10] , \u_div/CryTmp[3][1] , \u_div/CryTmp[3][2] ,
         \u_div/CryTmp[3][3] , \u_div/CryTmp[3][4] , \u_div/CryTmp[3][5] ,
         \u_div/CryTmp[3][6] , \u_div/CryTmp[3][7] , \u_div/CryTmp[3][8] ,
         \u_div/CryTmp[3][9] , \u_div/CryTmp[3][10] , \u_div/CryTmp[4][1] ,
         \u_div/CryTmp[4][2] , \u_div/CryTmp[4][3] , \u_div/CryTmp[4][4] ,
         \u_div/CryTmp[4][5] , \u_div/CryTmp[4][6] , \u_div/CryTmp[4][7] ,
         \u_div/CryTmp[4][8] , \u_div/CryTmp[4][9] , \u_div/CryTmp[4][10] ,
         \u_div/CryTmp[5][1] , \u_div/CryTmp[5][2] , \u_div/CryTmp[5][3] ,
         \u_div/CryTmp[5][4] , \u_div/CryTmp[5][5] , \u_div/CryTmp[5][6] ,
         \u_div/CryTmp[5][7] , \u_div/CryTmp[5][8] , \u_div/CryTmp[5][9] ,
         \u_div/CryTmp[5][10] , \u_div/CryTmp[6][1] , \u_div/CryTmp[6][2] ,
         \u_div/CryTmp[6][3] , \u_div/CryTmp[6][4] , \u_div/CryTmp[6][5] ,
         \u_div/CryTmp[6][6] , \u_div/CryTmp[6][7] , \u_div/CryTmp[6][8] ,
         \u_div/CryTmp[6][9] , \u_div/CryTmp[6][10] , \u_div/CryTmp[7][1] ,
         \u_div/CryTmp[7][2] , \u_div/CryTmp[7][3] , \u_div/CryTmp[7][4] ,
         \u_div/CryTmp[7][5] , \u_div/CryTmp[7][6] , \u_div/CryTmp[7][7] ,
         \u_div/CryTmp[7][8] , \u_div/CryTmp[7][9] , \u_div/CryTmp[7][10] ,
         \u_div/CryTmp[8][1] , \u_div/CryTmp[8][2] , \u_div/CryTmp[8][3] ,
         \u_div/CryTmp[8][4] , \u_div/CryTmp[8][5] , \u_div/CryTmp[8][6] ,
         \u_div/CryTmp[8][7] , \u_div/CryTmp[8][8] , \u_div/CryTmp[8][9] ,
         \u_div/CryTmp[8][10] , \u_div/CryTmp[9][1] , \u_div/CryTmp[9][2] ,
         \u_div/CryTmp[9][3] , \u_div/CryTmp[9][4] , \u_div/CryTmp[9][5] ,
         \u_div/CryTmp[9][6] , \u_div/CryTmp[9][7] , \u_div/CryTmp[9][8] ,
         \u_div/CryTmp[9][9] , \u_div/CryTmp[9][10] , \u_div/CryTmp[10][1] ,
         \u_div/CryTmp[10][2] , \u_div/CryTmp[10][3] , \u_div/CryTmp[10][4] ,
         \u_div/CryTmp[10][5] , \u_div/CryTmp[10][6] , \u_div/CryTmp[10][7] ,
         \u_div/CryTmp[10][8] , \u_div/CryTmp[10][9] , \u_div/CryTmp[10][10] ,
         \u_div/CryTmp[11][1] , \u_div/CryTmp[11][2] , \u_div/CryTmp[11][3] ,
         \u_div/CryTmp[11][4] , \u_div/CryTmp[11][5] , \u_div/CryTmp[11][6] ,
         \u_div/CryTmp[11][7] , \u_div/CryTmp[11][8] , \u_div/CryTmp[11][9] ,
         \u_div/CryTmp[11][10] , \u_div/CryTmp[12][1] , \u_div/CryTmp[12][2] ,
         \u_div/CryTmp[12][3] , \u_div/CryTmp[12][4] , \u_div/CryTmp[12][5] ,
         \u_div/CryTmp[12][6] , \u_div/CryTmp[12][7] , \u_div/CryTmp[12][8] ,
         \u_div/CryTmp[12][9] , \u_div/CryTmp[12][10] , \u_div/CryTmp[13][1] ,
         \u_div/CryTmp[13][2] , \u_div/CryTmp[13][3] , \u_div/CryTmp[13][4] ,
         \u_div/CryTmp[13][5] , \u_div/CryTmp[13][6] , \u_div/CryTmp[13][7] ,
         \u_div/CryTmp[13][8] , \u_div/CryTmp[13][9] , \u_div/CryTmp[13][10] ,
         \u_div/CryTmp[14][1] , \u_div/CryTmp[14][2] , \u_div/CryTmp[14][3] ,
         \u_div/CryTmp[14][4] , \u_div/CryTmp[14][5] , \u_div/CryTmp[14][6] ,
         \u_div/CryTmp[14][7] , \u_div/CryTmp[14][8] , \u_div/CryTmp[14][9] ,
         \u_div/CryTmp[14][10] , \u_div/CryTmp[15][1] , \u_div/CryTmp[15][2] ,
         \u_div/CryTmp[15][3] , \u_div/CryTmp[15][4] , \u_div/CryTmp[15][5] ,
         \u_div/CryTmp[15][6] , \u_div/CryTmp[15][7] , \u_div/CryTmp[15][8] ,
         \u_div/CryTmp[15][9] , \u_div/CryTmp[15][10] , \u_div/CryTmp[16][1] ,
         \u_div/CryTmp[16][2] , \u_div/CryTmp[16][3] , \u_div/CryTmp[16][4] ,
         \u_div/CryTmp[16][5] , \u_div/CryTmp[16][6] , \u_div/CryTmp[16][7] ,
         \u_div/CryTmp[16][8] , \u_div/CryTmp[16][9] , \u_div/CryTmp[16][10] ,
         \u_div/CryTmp[17][1] , \u_div/CryTmp[17][2] , \u_div/CryTmp[17][3] ,
         \u_div/CryTmp[17][4] , \u_div/CryTmp[17][5] , \u_div/CryTmp[17][6] ,
         \u_div/CryTmp[17][7] , \u_div/CryTmp[17][8] , \u_div/CryTmp[17][9] ,
         \u_div/CryTmp[17][10] , \u_div/CryTmp[18][1] , \u_div/CryTmp[18][2] ,
         \u_div/CryTmp[18][3] , \u_div/CryTmp[18][4] , \u_div/CryTmp[18][5] ,
         \u_div/CryTmp[18][6] , \u_div/CryTmp[18][7] , \u_div/CryTmp[18][8] ,
         \u_div/CryTmp[18][9] , \u_div/CryTmp[18][10] , \u_div/CryTmp[19][1] ,
         \u_div/CryTmp[19][2] , \u_div/CryTmp[19][3] , \u_div/CryTmp[19][4] ,
         \u_div/CryTmp[19][5] , \u_div/CryTmp[19][6] , \u_div/CryTmp[19][7] ,
         \u_div/CryTmp[19][8] , \u_div/CryTmp[19][9] , \u_div/CryTmp[19][10] ,
         \u_div/CryTmp[20][1] , \u_div/CryTmp[20][2] , \u_div/CryTmp[20][3] ,
         \u_div/CryTmp[20][4] , \u_div/CryTmp[20][5] , \u_div/CryTmp[20][6] ,
         \u_div/CryTmp[20][7] , \u_div/CryTmp[20][8] , \u_div/CryTmp[20][9] ,
         \u_div/CryTmp[20][10] , \u_div/CryTmp[21][1] , \u_div/CryTmp[21][2] ,
         \u_div/CryTmp[21][3] , \u_div/CryTmp[21][4] , \u_div/CryTmp[21][5] ,
         \u_div/CryTmp[21][6] , \u_div/CryTmp[21][7] , \u_div/CryTmp[21][8] ,
         \u_div/CryTmp[21][9] , \u_div/CryTmp[21][10] , \u_div/CryTmp[22][1] ,
         \u_div/CryTmp[22][2] , \u_div/CryTmp[22][3] , \u_div/CryTmp[22][4] ,
         \u_div/CryTmp[22][5] , \u_div/CryTmp[22][6] , \u_div/CryTmp[22][7] ,
         \u_div/CryTmp[22][8] , \u_div/CryTmp[22][9] , \u_div/CryTmp[23][1] ,
         \u_div/CryTmp[23][2] , \u_div/CryTmp[23][3] , \u_div/CryTmp[23][4] ,
         \u_div/CryTmp[23][5] , \u_div/CryTmp[23][6] , \u_div/CryTmp[23][7] ,
         \u_div/CryTmp[23][8] , \u_div/CryTmp[23][9] , \u_div/CryTmp[24][1] ,
         \u_div/CryTmp[24][2] , \u_div/CryTmp[24][3] , \u_div/CryTmp[24][4] ,
         \u_div/CryTmp[24][5] , \u_div/CryTmp[24][6] , \u_div/CryTmp[24][7] ,
         \u_div/CryTmp[24][8] , \u_div/CryTmp[25][1] , \u_div/CryTmp[25][2] ,
         \u_div/CryTmp[25][3] , \u_div/CryTmp[25][4] , \u_div/CryTmp[25][5] ,
         \u_div/CryTmp[25][6] , \u_div/CryTmp[25][7] , \u_div/CryTmp[26][1] ,
         \u_div/CryTmp[26][2] , \u_div/CryTmp[26][3] , \u_div/CryTmp[26][4] ,
         \u_div/CryTmp[26][5] , \u_div/CryTmp[26][6] , \u_div/CryTmp[27][1] ,
         \u_div/CryTmp[27][2] , \u_div/CryTmp[27][3] , \u_div/CryTmp[27][4] ,
         \u_div/CryTmp[27][5] , \u_div/CryTmp[28][1] , \u_div/CryTmp[28][2] ,
         \u_div/CryTmp[28][3] , \u_div/CryTmp[28][4] , \u_div/CryTmp[29][1] ,
         \u_div/CryTmp[29][2] , \u_div/CryTmp[29][3] , \u_div/CryTmp[30][1] ,
         \u_div/CryTmp[30][2] , \u_div/PartRem[1][2] , \u_div/PartRem[1][3] ,
         \u_div/PartRem[1][4] , \u_div/PartRem[1][5] , \u_div/PartRem[1][6] ,
         \u_div/PartRem[1][7] , \u_div/PartRem[1][8] , \u_div/PartRem[1][9] ,
         \u_div/PartRem[2][1] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[2][4] , \u_div/PartRem[2][5] , \u_div/PartRem[2][6] ,
         \u_div/PartRem[2][7] , \u_div/PartRem[2][8] , \u_div/PartRem[2][9] ,
         \u_div/PartRem[3][9] , \u_div/PartRem[4][9] , \u_div/PartRem[5][9] ,
         \u_div/PartRem[6][9] , \u_div/PartRem[7][9] , \u_div/PartRem[8][9] ,
         \u_div/PartRem[9][9] , \u_div/PartRem[10][9] , \u_div/PartRem[11][9] ,
         \u_div/PartRem[12][9] , \u_div/PartRem[13][9] ,
         \u_div/PartRem[14][9] , \u_div/PartRem[15][9] ,
         \u_div/PartRem[16][9] , \u_div/PartRem[17][9] ,
         \u_div/PartRem[18][9] , \u_div/PartRem[19][9] ,
         \u_div/PartRem[20][9] , \u_div/PartRem[21][9] ,
         \u_div/PartRem[22][9] , \u_div/PartRem[23][9] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304;
  wire   [9:0] \u_div/BInv ;

  ADDFX2 \u_div/u_fa_PartRem_0_20_9  ( .A(\u_div/PartRem[21][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[20][9] ), .CO(
        \u_div/CryTmp[20][10] ), .S(\u_div/SumTmp[20][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_9  ( .A(\u_div/PartRem[22][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[21][9] ), .CO(
        \u_div/CryTmp[21][10] ), .S(\u_div/SumTmp[21][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_9  ( .A(\u_div/PartRem[20][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[19][9] ), .CO(
        \u_div/CryTmp[19][10] ), .S(\u_div/SumTmp[19][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_9  ( .A(\u_div/PartRem[19][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[18][9] ), .CO(
        \u_div/CryTmp[18][10] ), .S(\u_div/SumTmp[18][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_9  ( .A(\u_div/PartRem[18][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[17][9] ), .CO(
        \u_div/CryTmp[17][10] ), .S(\u_div/SumTmp[17][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_9  ( .A(\u_div/PartRem[17][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[16][9] ), .CO(
        \u_div/CryTmp[16][10] ), .S(\u_div/SumTmp[16][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_9  ( .A(\u_div/PartRem[16][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[15][9] ), .CO(
        \u_div/CryTmp[15][10] ), .S(\u_div/SumTmp[15][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_9  ( .A(\u_div/PartRem[15][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[14][9] ), .CO(
        \u_div/CryTmp[14][10] ), .S(\u_div/SumTmp[14][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_9  ( .A(\u_div/PartRem[14][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[13][9] ), .CO(
        \u_div/CryTmp[13][10] ), .S(\u_div/SumTmp[13][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_9  ( .A(\u_div/PartRem[13][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[12][9] ), .CO(
        \u_div/CryTmp[12][10] ), .S(\u_div/SumTmp[12][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_9  ( .A(\u_div/PartRem[12][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[11][9] ), .CO(
        \u_div/CryTmp[11][10] ), .S(\u_div/SumTmp[11][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_9  ( .A(\u_div/PartRem[11][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[10][9] ), .CO(
        \u_div/CryTmp[10][10] ), .S(\u_div/SumTmp[10][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_9  ( .A(\u_div/PartRem[10][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[9][9] ), .CO(\u_div/CryTmp[9][10] ), .S(\u_div/SumTmp[9][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_9  ( .A(\u_div/PartRem[9][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[8][9] ), .CO(\u_div/CryTmp[8][10] ), .S(\u_div/SumTmp[8][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_9  ( .A(\u_div/PartRem[8][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[7][9] ), .CO(\u_div/CryTmp[7][10] ), .S(\u_div/SumTmp[7][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_9  ( .A(\u_div/PartRem[7][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[6][9] ), .CO(\u_div/CryTmp[6][10] ), .S(\u_div/SumTmp[6][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_9  ( .A(\u_div/PartRem[6][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[5][9] ), .CO(\u_div/CryTmp[5][10] ), .S(\u_div/SumTmp[5][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_9  ( .A(\u_div/PartRem[3][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[2][9] ), .CO(\u_div/CryTmp[2][10] ), .S(\u_div/SumTmp[2][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_9  ( .A(\u_div/PartRem[5][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[4][9] ), .CO(\u_div/CryTmp[4][10] ), .S(\u_div/SumTmp[4][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_9  ( .A(\u_div/PartRem[4][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[3][9] ), .CO(\u_div/CryTmp[3][10] ), .S(\u_div/SumTmp[3][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_9  ( .A(\u_div/PartRem[2][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[1][9] ), .CO(\u_div/CryTmp[1][10] ), .S(\u_div/SumTmp[1][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_22_8  ( .A(n227), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[22][8] ), .CO(\u_div/CryTmp[22][9] ), .S(
        \u_div/SumTmp[22][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_8  ( .A(n212), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[20][8] ), .CO(\u_div/CryTmp[20][9] ), .S(
        \u_div/SumTmp[20][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_8  ( .A(n210), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[21][8] ), .CO(\u_div/CryTmp[21][9] ), .S(
        \u_div/SumTmp[21][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_8  ( .A(n175), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[19][8] ), .CO(\u_div/CryTmp[19][9] ), .S(
        \u_div/SumTmp[19][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_8  ( .A(n207), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[18][8] ), .CO(\u_div/CryTmp[18][9] ), .S(
        \u_div/SumTmp[18][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_8  ( .A(n206), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[17][8] ), .CO(\u_div/CryTmp[17][9] ), .S(
        \u_div/SumTmp[17][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_8  ( .A(n205), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[16][8] ), .CO(\u_div/CryTmp[16][9] ), .S(
        \u_div/SumTmp[16][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_8  ( .A(n204), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[15][8] ), .CO(\u_div/CryTmp[15][9] ), .S(
        \u_div/SumTmp[15][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_8  ( .A(n202), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[14][8] ), .CO(\u_div/CryTmp[14][9] ), .S(
        \u_div/SumTmp[14][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_8  ( .A(n200), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[13][8] ), .CO(\u_div/CryTmp[13][9] ), .S(
        \u_div/SumTmp[13][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_8  ( .A(n198), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[12][8] ), .CO(\u_div/CryTmp[12][9] ), .S(
        \u_div/SumTmp[12][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_8  ( .A(n196), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[11][8] ), .CO(\u_div/CryTmp[11][9] ), .S(
        \u_div/SumTmp[11][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_8  ( .A(n194), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[10][8] ), .CO(\u_div/CryTmp[10][9] ), .S(
        \u_div/SumTmp[10][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_8  ( .A(n192), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[9][8] ), .CO(\u_div/CryTmp[9][9] ), .S(
        \u_div/SumTmp[9][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_8  ( .A(n190), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[8][8] ), .CO(\u_div/CryTmp[8][9] ), .S(
        \u_div/SumTmp[8][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_8  ( .A(n188), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[7][8] ), .CO(\u_div/CryTmp[7][9] ), .S(
        \u_div/SumTmp[7][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_8  ( .A(n186), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[6][8] ), .CO(\u_div/CryTmp[6][9] ), .S(
        \u_div/SumTmp[6][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_8  ( .A(n184), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[5][8] ), .CO(\u_div/CryTmp[5][9] ), .S(
        \u_div/SumTmp[5][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_8  ( .A(n183), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[4][8] ), .CO(\u_div/CryTmp[4][9] ), .S(
        \u_div/SumTmp[4][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_8  ( .A(n181), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[3][8] ), .CO(\u_div/CryTmp[3][9] ), .S(
        \u_div/SumTmp[3][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_7  ( .A(\u_div/PartRem[1][7] ), .B(
        \u_div/BInv [7]), .CI(\u_div/CryTmp[0][7] ), .CO(\u_div/CryTmp[0][8] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_8  ( .A(\u_div/PartRem[1][8] ), .B(
        \u_div/BInv [8]), .CI(\u_div/CryTmp[0][8] ), .CO(\u_div/CryTmp[0][9] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_8  ( .A(\u_div/PartRem[2][8] ), .B(
        \u_div/BInv [8]), .CI(\u_div/CryTmp[1][8] ), .CO(\u_div/CryTmp[1][9] ), 
        .S(\u_div/SumTmp[1][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_8  ( .A(n208), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[2][8] ), .CO(\u_div/CryTmp[2][9] ), .S(
        \u_div/SumTmp[2][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_23_7  ( .A(n213), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[23][7] ), .CO(\u_div/CryTmp[23][8] ), .S(
        \u_div/SumTmp[23][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_7  ( .A(n209), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[21][7] ), .CO(\u_div/CryTmp[21][8] ), .S(
        \u_div/SumTmp[21][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_22_7  ( .A(n226), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[22][7] ), .CO(\u_div/CryTmp[22][8] ), .S(
        \u_div/SumTmp[22][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_7  ( .A(n211), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[20][7] ), .CO(\u_div/CryTmp[20][8] ), .S(
        \u_div/SumTmp[20][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_7  ( .A(n174), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[19][7] ), .CO(\u_div/CryTmp[19][8] ), .S(
        \u_div/SumTmp[19][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_7  ( .A(n203), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[18][7] ), .CO(\u_div/CryTmp[18][8] ), .S(
        \u_div/SumTmp[18][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_7  ( .A(n201), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[17][7] ), .CO(\u_div/CryTmp[17][8] ), .S(
        \u_div/SumTmp[17][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_7  ( .A(n199), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[16][7] ), .CO(\u_div/CryTmp[16][8] ), .S(
        \u_div/SumTmp[16][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_7  ( .A(n197), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[15][7] ), .CO(\u_div/CryTmp[15][8] ), .S(
        \u_div/SumTmp[15][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_7  ( .A(n195), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[14][7] ), .CO(\u_div/CryTmp[14][8] ), .S(
        \u_div/SumTmp[14][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_7  ( .A(n193), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[13][7] ), .CO(\u_div/CryTmp[13][8] ), .S(
        \u_div/SumTmp[13][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_7  ( .A(n191), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[12][7] ), .CO(\u_div/CryTmp[12][8] ), .S(
        \u_div/SumTmp[12][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_7  ( .A(n189), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[11][7] ), .CO(\u_div/CryTmp[11][8] ), .S(
        \u_div/SumTmp[11][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_7  ( .A(n187), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[10][7] ), .CO(\u_div/CryTmp[10][8] ), .S(
        \u_div/SumTmp[10][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_7  ( .A(n185), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[9][7] ), .CO(\u_div/CryTmp[9][8] ), .S(
        \u_div/SumTmp[9][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_7  ( .A(n182), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[8][7] ), .CO(\u_div/CryTmp[8][8] ), .S(
        \u_div/SumTmp[8][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_7  ( .A(n180), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[7][7] ), .CO(\u_div/CryTmp[7][8] ), .S(
        \u_div/SumTmp[7][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_7  ( .A(n179), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[6][7] ), .CO(\u_div/CryTmp[6][8] ), .S(
        \u_div/SumTmp[6][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_7  ( .A(n178), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[5][7] ), .CO(\u_div/CryTmp[5][8] ), .S(
        \u_div/SumTmp[5][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_7  ( .A(n177), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[4][7] ), .CO(\u_div/CryTmp[4][8] ), .S(
        \u_div/SumTmp[4][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_7  ( .A(\u_div/PartRem[2][7] ), .B(
        \u_div/BInv [7]), .CI(\u_div/CryTmp[1][7] ), .CO(\u_div/CryTmp[1][8] ), 
        .S(\u_div/SumTmp[1][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_7  ( .A(n158), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[2][7] ), .CO(\u_div/CryTmp[2][8] ), .S(
        \u_div/SumTmp[2][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_7  ( .A(n176), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[3][7] ), .CO(\u_div/CryTmp[3][8] ), .S(
        \u_div/SumTmp[3][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_22_6  ( .A(n222), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[22][6] ), .CO(\u_div/CryTmp[22][7] ), .S(
        \u_div/SumTmp[22][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_23_6  ( .A(n167), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[23][6] ), .CO(\u_div/CryTmp[23][7] ), .S(
        \u_div/SumTmp[23][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_6  ( .A(n161), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[21][6] ), .CO(\u_div/CryTmp[21][7] ), .S(
        \u_div/SumTmp[21][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_6  ( .A(n164), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[20][6] ), .CO(\u_div/CryTmp[20][7] ), .S(
        \u_div/SumTmp[20][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_24_6  ( .A(n225), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[24][6] ), .CO(\u_div/CryTmp[24][7] ), .S(
        \u_div/SumTmp[24][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_6  ( .A(n107), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[19][6] ), .CO(\u_div/CryTmp[19][7] ), .S(
        \u_div/SumTmp[19][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_6  ( .A(n155), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[18][6] ), .CO(\u_div/CryTmp[18][7] ), .S(
        \u_div/SumTmp[18][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_6  ( .A(n154), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[17][6] ), .CO(\u_div/CryTmp[17][7] ), .S(
        \u_div/SumTmp[17][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_6  ( .A(n153), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[16][6] ), .CO(\u_div/CryTmp[16][7] ), .S(
        \u_div/SumTmp[16][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_6  ( .A(n152), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[15][6] ), .CO(\u_div/CryTmp[15][7] ), .S(
        \u_div/SumTmp[15][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_6  ( .A(n150), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[14][6] ), .CO(\u_div/CryTmp[14][7] ), .S(
        \u_div/SumTmp[14][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_6  ( .A(n148), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[13][6] ), .CO(\u_div/CryTmp[13][7] ), .S(
        \u_div/SumTmp[13][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_6  ( .A(n146), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[12][6] ), .CO(\u_div/CryTmp[12][7] ), .S(
        \u_div/SumTmp[12][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_6  ( .A(n144), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[11][6] ), .CO(\u_div/CryTmp[11][7] ), .S(
        \u_div/SumTmp[11][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_6  ( .A(n141), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[10][6] ), .CO(\u_div/CryTmp[10][7] ), .S(
        \u_div/SumTmp[10][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_6  ( .A(n138), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[9][6] ), .CO(\u_div/CryTmp[9][7] ), .S(
        \u_div/SumTmp[9][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_6  ( .A(n135), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[8][6] ), .CO(\u_div/CryTmp[8][7] ), .S(
        \u_div/SumTmp[8][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_6  ( .A(n132), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[7][6] ), .CO(\u_div/CryTmp[7][7] ), .S(
        \u_div/SumTmp[7][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_6  ( .A(n131), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[6][6] ), .CO(\u_div/CryTmp[6][7] ), .S(
        \u_div/SumTmp[6][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_5  ( .A(\u_div/PartRem[1][5] ), .B(
        \u_div/BInv [5]), .CI(\u_div/CryTmp[0][5] ), .CO(\u_div/CryTmp[0][6] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_6  ( .A(\u_div/PartRem[1][6] ), .B(
        \u_div/BInv [6]), .CI(\u_div/CryTmp[0][6] ), .CO(\u_div/CryTmp[0][7] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_5_6  ( .A(n128), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[5][6] ), .CO(\u_div/CryTmp[5][7] ), .S(
        \u_div/SumTmp[5][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_6  ( .A(\u_div/PartRem[2][6] ), .B(
        \u_div/BInv [6]), .CI(\u_div/CryTmp[1][6] ), .CO(\u_div/CryTmp[1][7] ), 
        .S(\u_div/SumTmp[1][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_6  ( .A(n157), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[2][6] ), .CO(\u_div/CryTmp[2][7] ), .S(
        \u_div/SumTmp[2][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_6  ( .A(n116), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[3][6] ), .CO(\u_div/CryTmp[3][7] ), .S(
        \u_div/SumTmp[3][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_6  ( .A(n114), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[4][6] ), .CO(\u_div/CryTmp[4][7] ), .S(
        \u_div/SumTmp[4][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_23_5  ( .A(n166), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[23][5] ), .CO(\u_div/CryTmp[23][6] ), .S(
        \u_div/SumTmp[23][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_24_5  ( .A(n224), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[24][5] ), .CO(\u_div/CryTmp[24][6] ), .S(
        \u_div/SumTmp[24][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_22_5  ( .A(n221), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[22][5] ), .CO(\u_div/CryTmp[22][6] ), .S(
        \u_div/SumTmp[22][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_5  ( .A(n160), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[21][5] ), .CO(\u_div/CryTmp[21][6] ), .S(
        \u_div/SumTmp[21][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_5  ( .A(n163), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[20][5] ), .CO(\u_div/CryTmp[20][6] ), .S(
        \u_div/SumTmp[20][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_5  ( .A(n106), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[19][5] ), .CO(\u_div/CryTmp[19][6] ), .S(
        \u_div/SumTmp[19][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_5  ( .A(n151), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[18][5] ), .CO(\u_div/CryTmp[18][6] ), .S(
        \u_div/SumTmp[18][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_5  ( .A(n149), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[17][5] ), .CO(\u_div/CryTmp[17][6] ), .S(
        \u_div/SumTmp[17][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_25_5  ( .A(n169), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[25][5] ), .CO(\u_div/CryTmp[25][6] ), .S(
        \u_div/SumTmp[25][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_5  ( .A(n147), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[16][5] ), .CO(\u_div/CryTmp[16][6] ), .S(
        \u_div/SumTmp[16][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_5  ( .A(n145), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[15][5] ), .CO(\u_div/CryTmp[15][6] ), .S(
        \u_div/SumTmp[15][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_5  ( .A(n142), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[14][5] ), .CO(\u_div/CryTmp[14][6] ), .S(
        \u_div/SumTmp[14][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_5  ( .A(n139), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[13][5] ), .CO(\u_div/CryTmp[13][6] ), .S(
        \u_div/SumTmp[13][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_5  ( .A(n136), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[12][5] ), .CO(\u_div/CryTmp[12][6] ), .S(
        \u_div/SumTmp[12][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_5  ( .A(n133), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[11][5] ), .CO(\u_div/CryTmp[11][6] ), .S(
        \u_div/SumTmp[11][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_5  ( .A(n129), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[10][5] ), .CO(\u_div/CryTmp[10][6] ), .S(
        \u_div/SumTmp[10][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_5  ( .A(n126), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[9][5] ), .CO(\u_div/CryTmp[9][6] ), .S(
        \u_div/SumTmp[9][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_5  ( .A(n124), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[8][5] ), .CO(\u_div/CryTmp[8][6] ), .S(
        \u_div/SumTmp[8][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_5  ( .A(n123), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[7][5] ), .CO(\u_div/CryTmp[7][6] ), .S(
        \u_div/SumTmp[7][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_5  ( .A(\u_div/PartRem[2][5] ), .B(
        \u_div/BInv [5]), .CI(\u_div/CryTmp[1][5] ), .CO(\u_div/CryTmp[1][6] ), 
        .S(\u_div/SumTmp[1][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_5  ( .A(n121), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[6][5] ), .CO(\u_div/CryTmp[6][6] ), .S(
        \u_div/SumTmp[6][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_5  ( .A(n156), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[2][5] ), .CO(\u_div/CryTmp[2][6] ), .S(
        \u_div/SumTmp[2][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_5  ( .A(n115), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[3][5] ), .CO(\u_div/CryTmp[3][6] ), .S(
        \u_div/SumTmp[3][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_5  ( .A(n112), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[4][5] ), .CO(\u_div/CryTmp[4][6] ), .S(
        \u_div/SumTmp[4][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_5  ( .A(n110), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[5][5] ), .CO(\u_div/CryTmp[5][6] ), .S(
        \u_div/SumTmp[5][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_24_4  ( .A(n223), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[24][4] ), .CO(\u_div/CryTmp[24][5] ), .S(
        \u_div/SumTmp[24][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_23_4  ( .A(n165), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[23][4] ), .CO(\u_div/CryTmp[23][5] ), .S(
        \u_div/SumTmp[23][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_22_4  ( .A(n220), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[22][4] ), .CO(\u_div/CryTmp[22][5] ), .S(
        \u_div/SumTmp[22][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_4  ( .A(n159), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[21][4] ), .CO(\u_div/CryTmp[21][5] ), .S(
        \u_div/SumTmp[21][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_4  ( .A(n162), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[20][4] ), .CO(\u_div/CryTmp[20][5] ), .S(
        \u_div/SumTmp[20][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_25_4  ( .A(n168), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[25][4] ), .CO(\u_div/CryTmp[25][5] ), .S(
        \u_div/SumTmp[25][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_4  ( .A(n105), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[19][4] ), .CO(\u_div/CryTmp[19][5] ), .S(
        \u_div/SumTmp[19][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_4  ( .A(n143), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[18][4] ), .CO(\u_div/CryTmp[18][5] ), .S(
        \u_div/SumTmp[18][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_26_4  ( .A(n171), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[26][4] ), .CO(\u_div/CryTmp[26][5] ), .S(
        \u_div/SumTmp[26][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_4  ( .A(n140), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[17][4] ), .CO(\u_div/CryTmp[17][5] ), .S(
        \u_div/SumTmp[17][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_4  ( .A(n137), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[16][4] ), .CO(\u_div/CryTmp[16][5] ), .S(
        \u_div/SumTmp[16][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_4  ( .A(n134), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[15][4] ), .CO(\u_div/CryTmp[15][5] ), .S(
        \u_div/SumTmp[15][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_4  ( .A(n130), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[14][4] ), .CO(\u_div/CryTmp[14][5] ), .S(
        \u_div/SumTmp[14][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_4  ( .A(n127), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[13][4] ), .CO(\u_div/CryTmp[13][5] ), .S(
        \u_div/SumTmp[13][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_3  ( .A(\u_div/PartRem[1][3] ), .B(
        \u_div/BInv [3]), .CI(\u_div/CryTmp[0][3] ), .CO(\u_div/CryTmp[0][4] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_4  ( .A(\u_div/PartRem[1][4] ), .B(
        \u_div/BInv [4]), .CI(\u_div/CryTmp[0][4] ), .CO(\u_div/CryTmp[0][5] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_12_4  ( .A(n125), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[12][4] ), .CO(\u_div/CryTmp[12][5] ), .S(
        \u_div/SumTmp[12][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_4  ( .A(n122), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[11][4] ), .CO(\u_div/CryTmp[11][5] ), .S(
        \u_div/SumTmp[11][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/BInv [4]), .CI(\u_div/CryTmp[1][4] ), .CO(\u_div/CryTmp[1][5] ), 
        .S(\u_div/SumTmp[1][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_4  ( .A(n120), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[10][4] ), .CO(\u_div/CryTmp[10][5] ), .S(
        \u_div/SumTmp[10][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_4  ( .A(n119), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[9][4] ), .CO(\u_div/CryTmp[9][5] ), .S(
        \u_div/SumTmp[9][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_4  ( .A(n118), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[8][4] ), .CO(\u_div/CryTmp[8][5] ), .S(
        \u_div/SumTmp[8][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_4  ( .A(n117), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[7][4] ), .CO(\u_div/CryTmp[7][5] ), .S(
        \u_div/SumTmp[7][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_4  ( .A(n89), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[2][4] ), .CO(\u_div/CryTmp[2][5] ), .S(
        \u_div/SumTmp[2][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_4  ( .A(n113), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[3][4] ), .CO(\u_div/CryTmp[3][5] ), .S(
        \u_div/SumTmp[3][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_4  ( .A(n111), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[4][4] ), .CO(\u_div/CryTmp[4][5] ), .S(
        \u_div/SumTmp[4][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_4  ( .A(n109), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[5][4] ), .CO(\u_div/CryTmp[5][5] ), .S(
        \u_div/SumTmp[5][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_4  ( .A(n108), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[6][4] ), .CO(\u_div/CryTmp[6][5] ), .S(
        \u_div/SumTmp[6][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_24_3  ( .A(n218), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[24][3] ), .CO(\u_div/CryTmp[24][4] ), .S(
        \u_div/SumTmp[24][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_23_3  ( .A(n95), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[23][3] ), .CO(\u_div/CryTmp[23][4] ), .S(
        \u_div/SumTmp[23][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_25_3  ( .A(n97), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[25][3] ), .CO(\u_div/CryTmp[25][4] ), .S(
        \u_div/SumTmp[25][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_22_3  ( .A(n216), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[22][3] ), .CO(\u_div/CryTmp[22][4] ), .S(
        \u_div/SumTmp[22][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_3  ( .A(n91), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[21][3] ), .CO(\u_div/CryTmp[21][4] ), .S(
        \u_div/SumTmp[21][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_26_3  ( .A(n99), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[26][3] ), .CO(\u_div/CryTmp[26][4] ), .S(
        \u_div/SumTmp[26][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_3  ( .A(n93), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[20][3] ), .CO(\u_div/CryTmp[20][4] ), .S(
        \u_div/SumTmp[20][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_3  ( .A(n54), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[19][3] ), .CO(\u_div/CryTmp[19][4] ), .S(
        \u_div/SumTmp[19][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_27_3  ( .A(n101), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[27][3] ), .CO(\u_div/CryTmp[27][4] ), .S(
        \u_div/SumTmp[27][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_3  ( .A(n86), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[18][3] ), .CO(\u_div/CryTmp[18][4] ), .S(
        \u_div/SumTmp[18][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_3  ( .A(n85), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[17][3] ), .CO(\u_div/CryTmp[17][4] ), .S(
        \u_div/SumTmp[17][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_3  ( .A(n84), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[16][3] ), .CO(\u_div/CryTmp[16][4] ), .S(
        \u_div/SumTmp[16][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_3  ( .A(n83), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[15][3] ), .CO(\u_div/CryTmp[15][4] ), .S(
        \u_div/SumTmp[15][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_3  ( .A(n81), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[14][3] ), .CO(\u_div/CryTmp[14][4] ), .S(
        \u_div/SumTmp[14][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/BInv [3]), .CI(\u_div/CryTmp[1][3] ), .CO(\u_div/CryTmp[1][4] ), 
        .S(\u_div/SumTmp[1][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_3  ( .A(n79), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[13][3] ), .CO(\u_div/CryTmp[13][4] ), .S(
        \u_div/SumTmp[13][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_3  ( .A(n77), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[12][3] ), .CO(\u_div/CryTmp[12][4] ), .S(
        \u_div/SumTmp[12][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_3  ( .A(n75), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[11][3] ), .CO(\u_div/CryTmp[11][4] ), .S(
        \u_div/SumTmp[11][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_3  ( .A(n88), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[2][3] ), .CO(\u_div/CryTmp[2][4] ), .S(
        \u_div/SumTmp[2][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_3  ( .A(n73), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[10][3] ), .CO(\u_div/CryTmp[10][4] ), .S(
        \u_div/SumTmp[10][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_3  ( .A(n72), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[9][3] ), .CO(\u_div/CryTmp[9][4] ), .S(
        \u_div/SumTmp[9][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_3  ( .A(n70), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[8][3] ), .CO(\u_div/CryTmp[8][4] ), .S(
        \u_div/SumTmp[8][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_3  ( .A(n69), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[3][3] ), .CO(\u_div/CryTmp[3][4] ), .S(
        \u_div/SumTmp[3][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_3  ( .A(n64), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[4][3] ), .CO(\u_div/CryTmp[4][4] ), .S(
        \u_div/SumTmp[4][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_3  ( .A(n61), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[5][3] ), .CO(\u_div/CryTmp[5][4] ), .S(
        \u_div/SumTmp[5][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_3  ( .A(n59), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[6][3] ), .CO(\u_div/CryTmp[6][4] ), .S(
        \u_div/SumTmp[6][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_3  ( .A(n57), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[7][3] ), .CO(\u_div/CryTmp[7][4] ), .S(
        \u_div/SumTmp[7][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_25_2  ( .A(n96), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[25][2] ), .CO(\u_div/CryTmp[25][3] ), .S(
        \u_div/SumTmp[25][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_24_2  ( .A(n217), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[24][2] ), .CO(\u_div/CryTmp[24][3] ), .S(
        \u_div/SumTmp[24][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_26_2  ( .A(n98), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[26][2] ), .CO(\u_div/CryTmp[26][3] ), .S(
        \u_div/SumTmp[26][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_23_2  ( .A(n94), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[23][2] ), .CO(\u_div/CryTmp[23][3] ), .S(
        \u_div/SumTmp[23][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_22_2  ( .A(n215), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[22][2] ), .CO(\u_div/CryTmp[22][3] ), .S(
        \u_div/SumTmp[22][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_27_2  ( .A(n100), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[27][2] ), .CO(\u_div/CryTmp[27][3] ), .S(
        \u_div/SumTmp[27][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_2  ( .A(n90), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[21][2] ), .CO(\u_div/CryTmp[21][3] ), .S(
        \u_div/SumTmp[21][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_2  ( .A(n92), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[20][2] ), .CO(\u_div/CryTmp[20][3] ), .S(
        \u_div/SumTmp[20][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_28_2  ( .A(n102), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[28][2] ), .CO(\u_div/CryTmp[28][3] ), .S(
        \u_div/SumTmp[28][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_2  ( .A(n53), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[19][2] ), .CO(\u_div/CryTmp[19][3] ), .S(
        \u_div/SumTmp[19][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_2  ( .A(n82), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[18][2] ), .CO(\u_div/CryTmp[18][3] ), .S(
        \u_div/SumTmp[18][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_2  ( .A(n80), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[17][2] ), .CO(\u_div/CryTmp[17][3] ), .S(
        \u_div/SumTmp[17][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/BInv [2]), .CI(\u_div/CryTmp[1][2] ), .CO(\u_div/CryTmp[1][3] ), 
        .S(\u_div/SumTmp[1][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_2  ( .A(n78), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[16][2] ), .CO(\u_div/CryTmp[16][3] ), .S(
        \u_div/SumTmp[16][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_2  ( .A(n76), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[15][2] ), .CO(\u_div/CryTmp[15][3] ), .S(
        \u_div/SumTmp[15][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_2  ( .A(n74), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[14][2] ), .CO(\u_div/CryTmp[14][3] ), .S(
        \u_div/SumTmp[14][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_2  ( .A(n87), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[2][2] ), .CO(\u_div/CryTmp[2][3] ), .S(
        \u_div/SumTmp[2][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_2  ( .A(n71), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[13][2] ), .CO(\u_div/CryTmp[13][3] ), .S(
        \u_div/SumTmp[13][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_2  ( .A(n68), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[12][2] ), .CO(\u_div/CryTmp[12][3] ), .S(
        \u_div/SumTmp[12][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_2  ( .A(n67), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[3][2] ), .CO(\u_div/CryTmp[3][3] ), .S(
        \u_div/SumTmp[3][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_2  ( .A(n66), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[11][2] ), .CO(\u_div/CryTmp[11][3] ), .S(
        \u_div/SumTmp[11][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_2  ( .A(n65), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[10][2] ), .CO(\u_div/CryTmp[10][3] ), .S(
        \u_div/SumTmp[10][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_2  ( .A(n63), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[9][2] ), .CO(\u_div/CryTmp[9][3] ), .S(
        \u_div/SumTmp[9][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_2  ( .A(n62), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[4][2] ), .CO(\u_div/CryTmp[4][3] ), .S(
        \u_div/SumTmp[4][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_2  ( .A(n60), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[5][2] ), .CO(\u_div/CryTmp[5][3] ), .S(
        \u_div/SumTmp[5][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_2  ( .A(n58), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[6][2] ), .CO(\u_div/CryTmp[6][3] ), .S(
        \u_div/SumTmp[6][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_2  ( .A(n56), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[7][2] ), .CO(\u_div/CryTmp[7][3] ), .S(
        \u_div/SumTmp[7][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_2  ( .A(n55), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[8][2] ), .CO(\u_div/CryTmp[8][3] ), .S(
        \u_div/SumTmp[8][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_26_1  ( .A(n46), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[26][1] ), .CO(\u_div/CryTmp[26][2] ), .S(
        \u_div/SumTmp[26][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_25_1  ( .A(n23), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[25][1] ), .CO(\u_div/CryTmp[25][2] ), .S(
        \u_div/SumTmp[25][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_27_1  ( .A(n47), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[27][1] ), .CO(\u_div/CryTmp[27][2] ), .S(
        \u_div/SumTmp[27][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_24_1  ( .A(n45), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[24][1] ), .CO(\u_div/CryTmp[24][2] ), .S(
        \u_div/SumTmp[24][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_23_1  ( .A(n44), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[23][2] ), .S(
        \u_div/SumTmp[23][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_28_1  ( .A(n48), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[28][1] ), .CO(\u_div/CryTmp[28][2] ), .S(
        \u_div/SumTmp[28][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_22_1  ( .A(n43), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[22][2] ), .S(
        \u_div/SumTmp[22][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_1  ( .A(n41), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[21][1] ), .CO(\u_div/CryTmp[21][2] ), .S(
        \u_div/SumTmp[21][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_29_1  ( .A(n49), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[29][1] ), .CO(\u_div/CryTmp[29][2] ), .S(
        \u_div/SumTmp[29][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_1  ( .A(n42), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[20][1] ), .CO(\u_div/CryTmp[20][2] ), .S(
        \u_div/SumTmp[20][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_1  ( .A(n40), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[19][1] ), .CO(\u_div/CryTmp[19][2] ), .S(
        \u_div/SumTmp[19][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_1  ( .A(n39), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[18][1] ), .CO(\u_div/CryTmp[18][2] ), .S(
        \u_div/SumTmp[18][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_1  ( .A(n38), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[17][1] ), .CO(\u_div/CryTmp[17][2] ), .S(
        \u_div/SumTmp[17][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_1  ( .A(n37), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[16][1] ), .CO(\u_div/CryTmp[16][2] ), .S(
        \u_div/SumTmp[16][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_1  ( .A(n36), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[15][1] ), .CO(\u_div/CryTmp[15][2] ), .S(
        \u_div/SumTmp[15][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_1  ( .A(n35), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[14][1] ), .CO(\u_div/CryTmp[14][2] ), .S(
        \u_div/SumTmp[14][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_1  ( .A(n34), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[13][1] ), .CO(\u_div/CryTmp[13][2] ), .S(
        \u_div/SumTmp[13][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_1  ( .A(n33), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[4][1] ), .CO(\u_div/CryTmp[4][2] ), .S(
        \u_div/SumTmp[4][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_1  ( .A(n32), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[12][1] ), .CO(\u_div/CryTmp[12][2] ), .S(
        \u_div/SumTmp[12][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_1  ( .A(n31), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[11][2] ), .S(
        \u_div/SumTmp[11][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_1  ( .A(n30), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[10][1] ), .CO(\u_div/CryTmp[10][2] ), .S(
        \u_div/SumTmp[10][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_1  ( .A(n29), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[5][1] ), .CO(\u_div/CryTmp[5][2] ), .S(
        \u_div/SumTmp[5][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_1  ( .A(n28), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[6][1] ), .CO(\u_div/CryTmp[6][2] ), .S(
        \u_div/SumTmp[6][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_1  ( .A(n27), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[7][1] ), .CO(\u_div/CryTmp[7][2] ), .S(
        \u_div/SumTmp[7][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_1  ( .A(n26), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[8][1] ), .CO(\u_div/CryTmp[8][2] ), .S(
        \u_div/SumTmp[8][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_1  ( .A(n25), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[9][1] ), .CO(\u_div/CryTmp[9][2] ), .S(
        \u_div/SumTmp[9][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_28_3  ( .A(n103), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[28][3] ), .CO(\u_div/CryTmp[28][4] ), .S(
        \u_div/SumTmp[28][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_23_8  ( .A(n214), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[23][8] ), .CO(\u_div/CryTmp[23][9] ), .S(
        \u_div/SumTmp[23][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_30_1  ( .A(n22), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[30][1] ), .CO(\u_div/CryTmp[30][2] ), .S(
        \u_div/SumTmp[30][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_26_5  ( .A(n172), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[26][5] ), .CO(\u_div/CryTmp[26][6] ), .S(
        \u_div/SumTmp[26][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_27_4  ( .A(n173), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[27][4] ), .CO(\u_div/CryTmp[27][5] ), .S(
        \u_div/SumTmp[27][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_29_2  ( .A(n104), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[29][2] ), .CO(\u_div/CryTmp[29][3] ), .S(
        \u_div/SumTmp[29][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_24_7  ( .A(n228), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[24][7] ), .CO(\u_div/CryTmp[24][8] ), .S(
        \u_div/SumTmp[24][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_25_6  ( .A(n170), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[25][6] ), .CO(\u_div/CryTmp[25][7] ), .S(
        \u_div/SumTmp[25][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_9  ( .A(\u_div/PartRem[1][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[0][9] ), .CO(\u_div/CryTmp[0][10] ) );
  ADDFXL \u_div/u_fa_PartRem_0_0_1  ( .A(n50), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[0][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/BInv [2]), .CI(\u_div/CryTmp[0][2] ), .CO(\u_div/CryTmp[0][3] )
         );
  ADDFXL \u_div/u_fa_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        \u_div/BInv [1]), .CI(\u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[1][2] ), 
        .S(\u_div/SumTmp[1][1] ) );
  ADDFXL \u_div/u_fa_PartRem_0_2_1  ( .A(n219), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[2][2] ), .S(
        \u_div/SumTmp[2][1] ) );
  ADDFXL \u_div/u_fa_PartRem_0_3_1  ( .A(n24), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[3][2] ), .S(
        \u_div/SumTmp[3][1] ) );
  ADDFX4 \u_div/u_fa_PartRem_0_22_9  ( .A(\u_div/PartRem[23][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[22][9] ), .CO(quotient[22]), .S(
        \u_div/SumTmp[22][9] ) );
  CLKINVX3 U1 ( .A(n304), .Y(quotient[23]) );
  CLKINVX3 U2 ( .A(n303), .Y(quotient[24]) );
  CLKINVX3 U3 ( .A(n301), .Y(quotient[25]) );
  MX2X1 U4 ( .A(n249), .B(n274), .S0(quotient[1]), .Y(n1) );
  MX2X1 U5 ( .A(n247), .B(n258), .S0(quotient[2]), .Y(n2) );
  MX2X1 U6 ( .A(n262), .B(n265), .S0(quotient[20]), .Y(n3) );
  MX2X1 U7 ( .A(n264), .B(n276), .S0(quotient[19]), .Y(n4) );
  MX2X1 U8 ( .A(n275), .B(n278), .S0(quotient[18]), .Y(n5) );
  MX2X1 U9 ( .A(n277), .B(n280), .S0(quotient[17]), .Y(n6) );
  MX2X1 U10 ( .A(n279), .B(n282), .S0(quotient[16]), .Y(n7) );
  MX2X1 U11 ( .A(n281), .B(n284), .S0(quotient[15]), .Y(n8) );
  MX2X1 U12 ( .A(n283), .B(n286), .S0(quotient[14]), .Y(n9) );
  MX2X1 U13 ( .A(n285), .B(n288), .S0(quotient[13]), .Y(n10) );
  MX2X1 U14 ( .A(n287), .B(n290), .S0(quotient[12]), .Y(n11) );
  MX2X1 U15 ( .A(n289), .B(n292), .S0(quotient[11]), .Y(n12) );
  MX2X1 U16 ( .A(n291), .B(n293), .S0(quotient[10]), .Y(n13) );
  MX2X1 U17 ( .A(n235), .B(n236), .S0(quotient[9]), .Y(n14) );
  MX2X1 U18 ( .A(n234), .B(n238), .S0(quotient[8]), .Y(n15) );
  MX2X1 U19 ( .A(n237), .B(n240), .S0(quotient[7]), .Y(n16) );
  MX2X1 U20 ( .A(n239), .B(n242), .S0(quotient[6]), .Y(n17) );
  MX2X1 U21 ( .A(n241), .B(n244), .S0(quotient[5]), .Y(n18) );
  MX2X1 U22 ( .A(n243), .B(n246), .S0(quotient[4]), .Y(n19) );
  MX2X1 U23 ( .A(n245), .B(n248), .S0(quotient[3]), .Y(n20) );
  MX2X1 U24 ( .A(n260), .B(n263), .S0(quotient[21]), .Y(n21) );
  MX2X1 U25 ( .A(a[31]), .B(\u_div/SumTmp[31][0] ), .S0(quotient[31]), .Y(n22)
         );
  MX2X1 U26 ( .A(a[30]), .B(\u_div/SumTmp[26][0] ), .S0(quotient[26]), .Y(n23)
         );
  MX2X1 U27 ( .A(a[4]), .B(\u_div/SumTmp[4][0] ), .S0(quotient[4]), .Y(n24) );
  MX2X1 U28 ( .A(a[10]), .B(\u_div/SumTmp[10][0] ), .S0(quotient[10]), .Y(n25)
         );
  MX2X1 U29 ( .A(a[9]), .B(\u_div/SumTmp[9][0] ), .S0(quotient[9]), .Y(n26) );
  MX2X1 U30 ( .A(a[8]), .B(\u_div/SumTmp[8][0] ), .S0(quotient[8]), .Y(n27) );
  MX2X1 U31 ( .A(a[7]), .B(\u_div/SumTmp[7][0] ), .S0(quotient[7]), .Y(n28) );
  MX2X1 U32 ( .A(a[6]), .B(\u_div/SumTmp[6][0] ), .S0(quotient[6]), .Y(n29) );
  MX2X1 U33 ( .A(a[11]), .B(\u_div/SumTmp[11][0] ), .S0(quotient[11]), .Y(n30)
         );
  MX2X1 U34 ( .A(a[12]), .B(\u_div/SumTmp[12][0] ), .S0(quotient[12]), .Y(n31)
         );
  MX2X1 U35 ( .A(a[13]), .B(\u_div/SumTmp[13][0] ), .S0(quotient[13]), .Y(n32)
         );
  MX2X1 U36 ( .A(a[5]), .B(\u_div/SumTmp[5][0] ), .S0(quotient[5]), .Y(n33) );
  MX2X1 U37 ( .A(a[14]), .B(\u_div/SumTmp[14][0] ), .S0(quotient[14]), .Y(n34)
         );
  MX2X1 U38 ( .A(a[15]), .B(\u_div/SumTmp[15][0] ), .S0(quotient[15]), .Y(n35)
         );
  MX2X1 U39 ( .A(a[16]), .B(\u_div/SumTmp[16][0] ), .S0(quotient[16]), .Y(n36)
         );
  MX2X1 U40 ( .A(a[17]), .B(\u_div/SumTmp[17][0] ), .S0(quotient[17]), .Y(n37)
         );
  MX2X1 U41 ( .A(a[18]), .B(\u_div/SumTmp[18][0] ), .S0(quotient[18]), .Y(n38)
         );
  MX2X1 U42 ( .A(a[19]), .B(\u_div/SumTmp[19][0] ), .S0(quotient[19]), .Y(n39)
         );
  MX2X1 U43 ( .A(a[20]), .B(\u_div/SumTmp[20][0] ), .S0(quotient[20]), .Y(n40)
         );
  MX2X1 U44 ( .A(a[30]), .B(\u_div/SumTmp[22][0] ), .S0(quotient[22]), .Y(n41)
         );
  MX2X1 U45 ( .A(a[21]), .B(\u_div/SumTmp[21][0] ), .S0(quotient[21]), .Y(n42)
         );
  MX2X1 U46 ( .A(a[30]), .B(\u_div/SumTmp[23][0] ), .S0(quotient[23]), .Y(n43)
         );
  MX2X1 U47 ( .A(a[30]), .B(\u_div/SumTmp[24][0] ), .S0(quotient[24]), .Y(n44)
         );
  MX2X1 U48 ( .A(a[30]), .B(\u_div/SumTmp[25][0] ), .S0(quotient[25]), .Y(n45)
         );
  MX2X1 U49 ( .A(a[30]), .B(\u_div/SumTmp[27][0] ), .S0(quotient[27]), .Y(n46)
         );
  MX2X1 U50 ( .A(a[30]), .B(\u_div/SumTmp[28][0] ), .S0(quotient[28]), .Y(n47)
         );
  MX2X1 U51 ( .A(a[30]), .B(\u_div/SumTmp[29][0] ), .S0(quotient[29]), .Y(n48)
         );
  MX2X1 U52 ( .A(a[30]), .B(\u_div/SumTmp[30][0] ), .S0(quotient[30]), .Y(n49)
         );
  AND2X2 U53 ( .A(quotient[1]), .B(b[0]), .Y(n50) );
  MX2X1 U54 ( .A(n259), .B(n261), .S0(quotient[22]), .Y(n51) );
  INVX12 U55 ( .A(b[0]), .Y(\u_div/CryTmp[3][1] ) );
  NOR2BXL U56 ( .AN(quotient[3]), .B(\u_div/CryTmp[3][1] ), .Y(n219) );
  NOR2XL U57 ( .A(a[31]), .B(\u_div/CryTmp[3][1] ), .Y(n231) );
  AND2X2 U58 ( .A(\u_div/CryTmp[26][6] ), .B(n232), .Y(quotient[26]) );
  INVX1 U59 ( .A(\u_div/SumTmp[21][9] ), .Y(n263) );
  INVX1 U60 ( .A(\u_div/SumTmp[5][9] ), .Y(n244) );
  INVX1 U61 ( .A(\u_div/SumTmp[6][9] ), .Y(n242) );
  INVX1 U62 ( .A(\u_div/SumTmp[7][9] ), .Y(n240) );
  INVX1 U63 ( .A(\u_div/SumTmp[8][9] ), .Y(n238) );
  INVX1 U64 ( .A(\u_div/SumTmp[9][9] ), .Y(n236) );
  INVX1 U65 ( .A(\u_div/SumTmp[10][9] ), .Y(n293) );
  INVX1 U66 ( .A(\u_div/SumTmp[11][9] ), .Y(n292) );
  INVX1 U67 ( .A(\u_div/SumTmp[12][9] ), .Y(n290) );
  INVX1 U68 ( .A(\u_div/SumTmp[13][9] ), .Y(n288) );
  INVX1 U69 ( .A(\u_div/SumTmp[14][9] ), .Y(n286) );
  INVX1 U70 ( .A(\u_div/SumTmp[15][9] ), .Y(n284) );
  INVX1 U71 ( .A(\u_div/SumTmp[16][9] ), .Y(n282) );
  INVX1 U72 ( .A(\u_div/SumTmp[17][9] ), .Y(n280) );
  INVX1 U73 ( .A(\u_div/SumTmp[18][9] ), .Y(n278) );
  INVX1 U74 ( .A(\u_div/SumTmp[19][9] ), .Y(n276) );
  INVX1 U75 ( .A(\u_div/SumTmp[20][9] ), .Y(n265) );
  INVX1 U76 ( .A(\u_div/SumTmp[3][9] ), .Y(n248) );
  INVX1 U77 ( .A(\u_div/SumTmp[4][9] ), .Y(n246) );
  INVX1 U78 ( .A(\u_div/SumTmp[2][9] ), .Y(n258) );
  INVX1 U79 ( .A(\u_div/SumTmp[22][9] ), .Y(n261) );
  MXI2X1 U80 ( .A(n219), .B(\u_div/SumTmp[2][1] ), .S0(quotient[2]), .Y(n256)
         );
  MXI2X1 U81 ( .A(n88), .B(\u_div/SumTmp[2][3] ), .S0(quotient[2]), .Y(n254)
         );
  MXI2X1 U82 ( .A(n87), .B(\u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(n255)
         );
  MXI2X1 U83 ( .A(n256), .B(n272), .S0(quotient[1]), .Y(\u_div/PartRem[1][3] )
         );
  INVX1 U84 ( .A(\u_div/SumTmp[1][2] ), .Y(n272) );
  MX2X1 U85 ( .A(n42), .B(\u_div/SumTmp[20][1] ), .S0(quotient[20]), .Y(n53)
         );
  MX2X1 U86 ( .A(n92), .B(\u_div/SumTmp[20][2] ), .S0(quotient[20]), .Y(n54)
         );
  MX2X1 U87 ( .A(n25), .B(\u_div/SumTmp[9][1] ), .S0(quotient[9]), .Y(n55) );
  MX2X1 U88 ( .A(n26), .B(\u_div/SumTmp[8][1] ), .S0(quotient[8]), .Y(n56) );
  MX2X1 U89 ( .A(n55), .B(\u_div/SumTmp[8][2] ), .S0(quotient[8]), .Y(n57) );
  MX2X1 U90 ( .A(n27), .B(\u_div/SumTmp[7][1] ), .S0(quotient[7]), .Y(n58) );
  MX2X1 U91 ( .A(n56), .B(\u_div/SumTmp[7][2] ), .S0(quotient[7]), .Y(n59) );
  MX2X1 U92 ( .A(n28), .B(\u_div/SumTmp[6][1] ), .S0(quotient[6]), .Y(n60) );
  MX2X1 U93 ( .A(n58), .B(\u_div/SumTmp[6][2] ), .S0(quotient[6]), .Y(n61) );
  MX2X1 U94 ( .A(n29), .B(\u_div/SumTmp[5][1] ), .S0(quotient[5]), .Y(n62) );
  MX2X1 U95 ( .A(n30), .B(\u_div/SumTmp[10][1] ), .S0(quotient[10]), .Y(n63)
         );
  MX2X1 U96 ( .A(n60), .B(\u_div/SumTmp[5][2] ), .S0(quotient[5]), .Y(n64) );
  MX2X1 U97 ( .A(n31), .B(\u_div/SumTmp[11][1] ), .S0(quotient[11]), .Y(n65)
         );
  MX2X1 U98 ( .A(n32), .B(\u_div/SumTmp[12][1] ), .S0(quotient[12]), .Y(n66)
         );
  MX2X1 U99 ( .A(n33), .B(\u_div/SumTmp[4][1] ), .S0(quotient[4]), .Y(n67) );
  MX2X1 U100 ( .A(n34), .B(\u_div/SumTmp[13][1] ), .S0(quotient[13]), .Y(n68)
         );
  MX2X1 U101 ( .A(n62), .B(\u_div/SumTmp[4][2] ), .S0(quotient[4]), .Y(n69) );
  MX2X1 U102 ( .A(n63), .B(\u_div/SumTmp[9][2] ), .S0(quotient[9]), .Y(n70) );
  MX2X1 U103 ( .A(n35), .B(\u_div/SumTmp[14][1] ), .S0(quotient[14]), .Y(n71)
         );
  MX2X1 U104 ( .A(n65), .B(\u_div/SumTmp[10][2] ), .S0(quotient[10]), .Y(n72)
         );
  MX2X1 U105 ( .A(n66), .B(\u_div/SumTmp[11][2] ), .S0(quotient[11]), .Y(n73)
         );
  MX2X1 U106 ( .A(n36), .B(\u_div/SumTmp[15][1] ), .S0(quotient[15]), .Y(n74)
         );
  MX2X1 U107 ( .A(n68), .B(\u_div/SumTmp[12][2] ), .S0(quotient[12]), .Y(n75)
         );
  MX2X1 U108 ( .A(n37), .B(\u_div/SumTmp[16][1] ), .S0(quotient[16]), .Y(n76)
         );
  MX2X1 U109 ( .A(n71), .B(\u_div/SumTmp[13][2] ), .S0(quotient[13]), .Y(n77)
         );
  MX2X1 U110 ( .A(n38), .B(\u_div/SumTmp[17][1] ), .S0(quotient[17]), .Y(n78)
         );
  MX2X1 U111 ( .A(n74), .B(\u_div/SumTmp[14][2] ), .S0(quotient[14]), .Y(n79)
         );
  MX2X1 U112 ( .A(n39), .B(\u_div/SumTmp[18][1] ), .S0(quotient[18]), .Y(n80)
         );
  MX2X1 U113 ( .A(n76), .B(\u_div/SumTmp[15][2] ), .S0(quotient[15]), .Y(n81)
         );
  MX2X1 U114 ( .A(n40), .B(\u_div/SumTmp[19][1] ), .S0(quotient[19]), .Y(n82)
         );
  MX2X1 U115 ( .A(n78), .B(\u_div/SumTmp[16][2] ), .S0(quotient[16]), .Y(n83)
         );
  MX2X1 U116 ( .A(n80), .B(\u_div/SumTmp[17][2] ), .S0(quotient[17]), .Y(n84)
         );
  MX2X1 U117 ( .A(n82), .B(\u_div/SumTmp[18][2] ), .S0(quotient[18]), .Y(n85)
         );
  MX2X1 U118 ( .A(n53), .B(\u_div/SumTmp[19][2] ), .S0(quotient[19]), .Y(n86)
         );
  MX2X1 U119 ( .A(n24), .B(\u_div/SumTmp[3][1] ), .S0(quotient[3]), .Y(n87) );
  MX2X1 U120 ( .A(n67), .B(\u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(n88) );
  MX2X1 U121 ( .A(n69), .B(\u_div/SumTmp[3][3] ), .S0(quotient[3]), .Y(n89) );
  MX2X1 U122 ( .A(n43), .B(\u_div/SumTmp[22][1] ), .S0(quotient[22]), .Y(n90)
         );
  MX2X1 U123 ( .A(n215), .B(\u_div/SumTmp[22][2] ), .S0(quotient[22]), .Y(n91)
         );
  MX2X1 U124 ( .A(n41), .B(\u_div/SumTmp[21][1] ), .S0(quotient[21]), .Y(n92)
         );
  MX2X1 U125 ( .A(n90), .B(\u_div/SumTmp[21][2] ), .S0(quotient[21]), .Y(n93)
         );
  MX2X1 U126 ( .A(n45), .B(\u_div/SumTmp[24][1] ), .S0(quotient[24]), .Y(n94)
         );
  MX2X1 U127 ( .A(n217), .B(\u_div/SumTmp[24][2] ), .S0(quotient[24]), .Y(n95)
         );
  MX2X1 U128 ( .A(n46), .B(\u_div/SumTmp[26][1] ), .S0(quotient[26]), .Y(n96)
         );
  MX2X1 U129 ( .A(n98), .B(\u_div/SumTmp[26][2] ), .S0(quotient[26]), .Y(n97)
         );
  MX2X1 U130 ( .A(n47), .B(\u_div/SumTmp[27][1] ), .S0(quotient[27]), .Y(n98)
         );
  MX2X1 U131 ( .A(n100), .B(\u_div/SumTmp[27][2] ), .S0(quotient[27]), .Y(n99)
         );
  MX2X1 U132 ( .A(n48), .B(\u_div/SumTmp[28][1] ), .S0(quotient[28]), .Y(n100)
         );
  MX2X1 U133 ( .A(n102), .B(\u_div/SumTmp[28][2] ), .S0(quotient[28]), .Y(n101) );
  MX2X1 U134 ( .A(n49), .B(\u_div/SumTmp[29][1] ), .S0(quotient[29]), .Y(n102)
         );
  MX2X1 U135 ( .A(n104), .B(\u_div/SumTmp[29][2] ), .S0(quotient[29]), .Y(n103) );
  MX2X1 U136 ( .A(n22), .B(\u_div/SumTmp[30][1] ), .S0(quotient[30]), .Y(n104)
         );
  MXI2X1 U137 ( .A(n156), .B(\u_div/SumTmp[2][5] ), .S0(quotient[2]), .Y(n252)
         );
  MXI2X1 U138 ( .A(n89), .B(\u_div/SumTmp[2][4] ), .S0(quotient[2]), .Y(n253)
         );
  MXI2X1 U139 ( .A(n157), .B(\u_div/SumTmp[2][6] ), .S0(quotient[2]), .Y(n251)
         );
  MXI2X1 U140 ( .A(n254), .B(n270), .S0(quotient[1]), .Y(\u_div/PartRem[1][5] ) );
  INVX1 U141 ( .A(\u_div/SumTmp[1][4] ), .Y(n270) );
  MX2X1 U142 ( .A(n93), .B(\u_div/SumTmp[20][3] ), .S0(quotient[20]), .Y(n105)
         );
  MX2X1 U143 ( .A(n162), .B(\u_div/SumTmp[20][4] ), .S0(quotient[20]), .Y(n106) );
  MX2X1 U144 ( .A(n163), .B(\u_div/SumTmp[20][5] ), .S0(quotient[20]), .Y(n107) );
  MX2X1 U145 ( .A(n57), .B(\u_div/SumTmp[7][3] ), .S0(quotient[7]), .Y(n108)
         );
  MX2X1 U146 ( .A(n59), .B(\u_div/SumTmp[6][3] ), .S0(quotient[6]), .Y(n109)
         );
  MX2X1 U147 ( .A(n108), .B(\u_div/SumTmp[6][4] ), .S0(quotient[6]), .Y(n110)
         );
  MX2X1 U148 ( .A(n61), .B(\u_div/SumTmp[5][3] ), .S0(quotient[5]), .Y(n111)
         );
  MX2X1 U149 ( .A(n109), .B(\u_div/SumTmp[5][4] ), .S0(quotient[5]), .Y(n112)
         );
  MX2X1 U150 ( .A(n64), .B(\u_div/SumTmp[4][3] ), .S0(quotient[4]), .Y(n113)
         );
  MX2X1 U151 ( .A(n110), .B(\u_div/SumTmp[5][5] ), .S0(quotient[5]), .Y(n114)
         );
  MX2X1 U152 ( .A(n111), .B(\u_div/SumTmp[4][4] ), .S0(quotient[4]), .Y(n115)
         );
  MX2X1 U153 ( .A(n112), .B(\u_div/SumTmp[4][5] ), .S0(quotient[4]), .Y(n116)
         );
  MX2X1 U154 ( .A(n70), .B(\u_div/SumTmp[8][3] ), .S0(quotient[8]), .Y(n117)
         );
  MX2X1 U155 ( .A(n72), .B(\u_div/SumTmp[9][3] ), .S0(quotient[9]), .Y(n118)
         );
  MX2X1 U156 ( .A(n73), .B(\u_div/SumTmp[10][3] ), .S0(quotient[10]), .Y(n119)
         );
  MX2X1 U157 ( .A(n75), .B(\u_div/SumTmp[11][3] ), .S0(quotient[11]), .Y(n120)
         );
  MX2X1 U158 ( .A(n117), .B(\u_div/SumTmp[7][4] ), .S0(quotient[7]), .Y(n121)
         );
  MX2X1 U159 ( .A(n77), .B(\u_div/SumTmp[12][3] ), .S0(quotient[12]), .Y(n122)
         );
  MX2X1 U160 ( .A(n118), .B(\u_div/SumTmp[8][4] ), .S0(quotient[8]), .Y(n123)
         );
  MX2X1 U161 ( .A(n119), .B(\u_div/SumTmp[9][4] ), .S0(quotient[9]), .Y(n124)
         );
  MX2X1 U162 ( .A(n79), .B(\u_div/SumTmp[13][3] ), .S0(quotient[13]), .Y(n125)
         );
  MX2X1 U163 ( .A(n120), .B(\u_div/SumTmp[10][4] ), .S0(quotient[10]), .Y(n126) );
  MX2X1 U164 ( .A(n81), .B(\u_div/SumTmp[14][3] ), .S0(quotient[14]), .Y(n127)
         );
  MX2X1 U165 ( .A(n121), .B(\u_div/SumTmp[6][5] ), .S0(quotient[6]), .Y(n128)
         );
  MX2X1 U166 ( .A(n122), .B(\u_div/SumTmp[11][4] ), .S0(quotient[11]), .Y(n129) );
  MX2X1 U167 ( .A(n83), .B(\u_div/SumTmp[15][3] ), .S0(quotient[15]), .Y(n130)
         );
  MX2X1 U168 ( .A(n123), .B(\u_div/SumTmp[7][5] ), .S0(quotient[7]), .Y(n131)
         );
  MX2X1 U169 ( .A(n124), .B(\u_div/SumTmp[8][5] ), .S0(quotient[8]), .Y(n132)
         );
  MX2X1 U170 ( .A(n125), .B(\u_div/SumTmp[12][4] ), .S0(quotient[12]), .Y(n133) );
  MX2X1 U171 ( .A(n84), .B(\u_div/SumTmp[16][3] ), .S0(quotient[16]), .Y(n134)
         );
  MX2X1 U172 ( .A(n126), .B(\u_div/SumTmp[9][5] ), .S0(quotient[9]), .Y(n135)
         );
  MX2X1 U173 ( .A(n127), .B(\u_div/SumTmp[13][4] ), .S0(quotient[13]), .Y(n136) );
  MX2X1 U174 ( .A(n85), .B(\u_div/SumTmp[17][3] ), .S0(quotient[17]), .Y(n137)
         );
  MX2X1 U175 ( .A(n129), .B(\u_div/SumTmp[10][5] ), .S0(quotient[10]), .Y(n138) );
  MX2X1 U176 ( .A(n130), .B(\u_div/SumTmp[14][4] ), .S0(quotient[14]), .Y(n139) );
  MX2X1 U177 ( .A(n86), .B(\u_div/SumTmp[18][3] ), .S0(quotient[18]), .Y(n140)
         );
  MX2X1 U178 ( .A(n133), .B(\u_div/SumTmp[11][5] ), .S0(quotient[11]), .Y(n141) );
  MX2X1 U179 ( .A(n134), .B(\u_div/SumTmp[15][4] ), .S0(quotient[15]), .Y(n142) );
  MX2X1 U180 ( .A(n54), .B(\u_div/SumTmp[19][3] ), .S0(quotient[19]), .Y(n143)
         );
  MX2X1 U181 ( .A(n136), .B(\u_div/SumTmp[12][5] ), .S0(quotient[12]), .Y(n144) );
  MX2X1 U182 ( .A(n137), .B(\u_div/SumTmp[16][4] ), .S0(quotient[16]), .Y(n145) );
  MX2X1 U183 ( .A(n139), .B(\u_div/SumTmp[13][5] ), .S0(quotient[13]), .Y(n146) );
  MX2X1 U184 ( .A(n140), .B(\u_div/SumTmp[17][4] ), .S0(quotient[17]), .Y(n147) );
  MX2X1 U185 ( .A(n142), .B(\u_div/SumTmp[14][5] ), .S0(quotient[14]), .Y(n148) );
  MX2X1 U186 ( .A(n143), .B(\u_div/SumTmp[18][4] ), .S0(quotient[18]), .Y(n149) );
  MX2X1 U187 ( .A(n145), .B(\u_div/SumTmp[15][5] ), .S0(quotient[15]), .Y(n150) );
  MX2X1 U188 ( .A(n105), .B(\u_div/SumTmp[19][4] ), .S0(quotient[19]), .Y(n151) );
  MX2X1 U189 ( .A(n147), .B(\u_div/SumTmp[16][5] ), .S0(quotient[16]), .Y(n152) );
  MX2X1 U190 ( .A(n149), .B(\u_div/SumTmp[17][5] ), .S0(quotient[17]), .Y(n153) );
  MX2X1 U191 ( .A(n151), .B(\u_div/SumTmp[18][5] ), .S0(quotient[18]), .Y(n154) );
  MX2X1 U192 ( .A(n106), .B(\u_div/SumTmp[19][5] ), .S0(quotient[19]), .Y(n155) );
  MX2X1 U193 ( .A(n113), .B(\u_div/SumTmp[3][4] ), .S0(quotient[3]), .Y(n156)
         );
  MX2X1 U194 ( .A(n115), .B(\u_div/SumTmp[3][5] ), .S0(quotient[3]), .Y(n157)
         );
  MX2X1 U195 ( .A(n116), .B(\u_div/SumTmp[3][6] ), .S0(quotient[3]), .Y(n158)
         );
  MX2X1 U196 ( .A(n216), .B(\u_div/SumTmp[22][3] ), .S0(quotient[22]), .Y(n159) );
  MX2X1 U197 ( .A(n220), .B(\u_div/SumTmp[22][4] ), .S0(quotient[22]), .Y(n160) );
  MX2X1 U198 ( .A(n221), .B(\u_div/SumTmp[22][5] ), .S0(quotient[22]), .Y(n161) );
  MX2X1 U199 ( .A(n91), .B(\u_div/SumTmp[21][3] ), .S0(quotient[21]), .Y(n162)
         );
  MX2X1 U200 ( .A(n159), .B(\u_div/SumTmp[21][4] ), .S0(quotient[21]), .Y(n163) );
  MX2X1 U201 ( .A(n160), .B(\u_div/SumTmp[21][5] ), .S0(quotient[21]), .Y(n164) );
  MX2X1 U202 ( .A(n218), .B(\u_div/SumTmp[24][3] ), .S0(quotient[24]), .Y(n165) );
  MX2X1 U203 ( .A(n223), .B(\u_div/SumTmp[24][4] ), .S0(quotient[24]), .Y(n166) );
  MX2X1 U204 ( .A(n224), .B(\u_div/SumTmp[24][5] ), .S0(quotient[24]), .Y(n167) );
  MX2X1 U205 ( .A(n99), .B(\u_div/SumTmp[26][3] ), .S0(quotient[26]), .Y(n168)
         );
  MX2X1 U206 ( .A(n171), .B(\u_div/SumTmp[26][4] ), .S0(quotient[26]), .Y(n169) );
  MX2X1 U207 ( .A(n172), .B(\u_div/SumTmp[26][5] ), .S0(quotient[26]), .Y(n170) );
  MX2X1 U208 ( .A(n101), .B(\u_div/SumTmp[27][3] ), .S0(quotient[27]), .Y(n171) );
  MX2X1 U209 ( .A(n173), .B(\u_div/SumTmp[27][4] ), .S0(quotient[27]), .Y(n172) );
  MX2X1 U210 ( .A(n103), .B(\u_div/SumTmp[28][3] ), .S0(quotient[28]), .Y(n173) );
  MXI2X1 U211 ( .A(n212), .B(\u_div/SumTmp[20][8] ), .S0(quotient[20]), .Y(
        n264) );
  MXI2X1 U212 ( .A(n183), .B(\u_div/SumTmp[4][8] ), .S0(quotient[4]), .Y(n245)
         );
  MXI2X1 U213 ( .A(n184), .B(\u_div/SumTmp[5][8] ), .S0(quotient[5]), .Y(n243)
         );
  MXI2X1 U214 ( .A(n186), .B(\u_div/SumTmp[6][8] ), .S0(quotient[6]), .Y(n241)
         );
  MXI2X1 U215 ( .A(n188), .B(\u_div/SumTmp[7][8] ), .S0(quotient[7]), .Y(n239)
         );
  MXI2X1 U216 ( .A(n190), .B(\u_div/SumTmp[8][8] ), .S0(quotient[8]), .Y(n237)
         );
  MXI2X1 U217 ( .A(n192), .B(\u_div/SumTmp[9][8] ), .S0(quotient[9]), .Y(n234)
         );
  MXI2X1 U218 ( .A(n194), .B(\u_div/SumTmp[10][8] ), .S0(quotient[10]), .Y(
        n235) );
  MXI2X1 U219 ( .A(n196), .B(\u_div/SumTmp[11][8] ), .S0(quotient[11]), .Y(
        n291) );
  MXI2X1 U220 ( .A(n198), .B(\u_div/SumTmp[12][8] ), .S0(quotient[12]), .Y(
        n289) );
  MXI2X1 U221 ( .A(n200), .B(\u_div/SumTmp[13][8] ), .S0(quotient[13]), .Y(
        n287) );
  MXI2X1 U222 ( .A(n202), .B(\u_div/SumTmp[14][8] ), .S0(quotient[14]), .Y(
        n285) );
  MXI2X1 U223 ( .A(n204), .B(\u_div/SumTmp[15][8] ), .S0(quotient[15]), .Y(
        n283) );
  MXI2X1 U224 ( .A(n205), .B(\u_div/SumTmp[16][8] ), .S0(quotient[16]), .Y(
        n281) );
  MXI2X1 U225 ( .A(n206), .B(\u_div/SumTmp[17][8] ), .S0(quotient[17]), .Y(
        n279) );
  MXI2X1 U226 ( .A(n207), .B(\u_div/SumTmp[18][8] ), .S0(quotient[18]), .Y(
        n277) );
  MXI2X1 U227 ( .A(n175), .B(\u_div/SumTmp[19][8] ), .S0(quotient[19]), .Y(
        n275) );
  MXI2X1 U228 ( .A(n158), .B(\u_div/SumTmp[2][7] ), .S0(quotient[2]), .Y(n250)
         );
  MXI2X1 U229 ( .A(n208), .B(\u_div/SumTmp[2][8] ), .S0(quotient[2]), .Y(n249)
         );
  MXI2X1 U230 ( .A(n181), .B(\u_div/SumTmp[3][8] ), .S0(quotient[3]), .Y(n247)
         );
  MXI2X1 U231 ( .A(n227), .B(\u_div/SumTmp[22][8] ), .S0(quotient[22]), .Y(
        n260) );
  MXI2X1 U232 ( .A(n210), .B(\u_div/SumTmp[21][8] ), .S0(quotient[21]), .Y(
        n262) );
  MXI2X1 U233 ( .A(n252), .B(n268), .S0(quotient[1]), .Y(\u_div/PartRem[1][7] ) );
  INVX1 U234 ( .A(\u_div/SumTmp[1][6] ), .Y(n268) );
  MXI2X1 U235 ( .A(n250), .B(n266), .S0(quotient[1]), .Y(\u_div/PartRem[1][9] ) );
  INVX1 U236 ( .A(\u_div/SumTmp[1][8] ), .Y(n266) );
  MX2X1 U237 ( .A(n164), .B(\u_div/SumTmp[20][6] ), .S0(quotient[20]), .Y(n174) );
  MX2X1 U238 ( .A(n211), .B(\u_div/SumTmp[20][7] ), .S0(quotient[20]), .Y(n175) );
  MX2X1 U239 ( .A(n114), .B(\u_div/SumTmp[4][6] ), .S0(quotient[4]), .Y(n176)
         );
  MX2X1 U240 ( .A(n128), .B(\u_div/SumTmp[5][6] ), .S0(quotient[5]), .Y(n177)
         );
  MX2X1 U241 ( .A(n131), .B(\u_div/SumTmp[6][6] ), .S0(quotient[6]), .Y(n178)
         );
  MX2X1 U242 ( .A(n132), .B(\u_div/SumTmp[7][6] ), .S0(quotient[7]), .Y(n179)
         );
  MX2X1 U243 ( .A(n135), .B(\u_div/SumTmp[8][6] ), .S0(quotient[8]), .Y(n180)
         );
  MX2X1 U244 ( .A(n177), .B(\u_div/SumTmp[4][7] ), .S0(quotient[4]), .Y(n181)
         );
  MX2X1 U245 ( .A(n138), .B(\u_div/SumTmp[9][6] ), .S0(quotient[9]), .Y(n182)
         );
  MX2X1 U246 ( .A(n178), .B(\u_div/SumTmp[5][7] ), .S0(quotient[5]), .Y(n183)
         );
  MX2X1 U247 ( .A(n179), .B(\u_div/SumTmp[6][7] ), .S0(quotient[6]), .Y(n184)
         );
  MX2X1 U248 ( .A(n141), .B(\u_div/SumTmp[10][6] ), .S0(quotient[10]), .Y(n185) );
  MX2X1 U249 ( .A(n180), .B(\u_div/SumTmp[7][7] ), .S0(quotient[7]), .Y(n186)
         );
  MX2X1 U250 ( .A(n144), .B(\u_div/SumTmp[11][6] ), .S0(quotient[11]), .Y(n187) );
  MX2X1 U251 ( .A(n182), .B(\u_div/SumTmp[8][7] ), .S0(quotient[8]), .Y(n188)
         );
  MX2X1 U252 ( .A(n146), .B(\u_div/SumTmp[12][6] ), .S0(quotient[12]), .Y(n189) );
  MX2X1 U253 ( .A(n185), .B(\u_div/SumTmp[9][7] ), .S0(quotient[9]), .Y(n190)
         );
  MX2X1 U254 ( .A(n148), .B(\u_div/SumTmp[13][6] ), .S0(quotient[13]), .Y(n191) );
  MX2X1 U255 ( .A(n187), .B(\u_div/SumTmp[10][7] ), .S0(quotient[10]), .Y(n192) );
  MX2X1 U256 ( .A(n150), .B(\u_div/SumTmp[14][6] ), .S0(quotient[14]), .Y(n193) );
  MX2X1 U257 ( .A(n189), .B(\u_div/SumTmp[11][7] ), .S0(quotient[11]), .Y(n194) );
  MX2X1 U258 ( .A(n152), .B(\u_div/SumTmp[15][6] ), .S0(quotient[15]), .Y(n195) );
  MX2X1 U259 ( .A(n191), .B(\u_div/SumTmp[12][7] ), .S0(quotient[12]), .Y(n196) );
  MX2X1 U260 ( .A(n153), .B(\u_div/SumTmp[16][6] ), .S0(quotient[16]), .Y(n197) );
  MX2X1 U261 ( .A(n193), .B(\u_div/SumTmp[13][7] ), .S0(quotient[13]), .Y(n198) );
  MX2X1 U262 ( .A(n154), .B(\u_div/SumTmp[17][6] ), .S0(quotient[17]), .Y(n199) );
  MX2X1 U263 ( .A(n195), .B(\u_div/SumTmp[14][7] ), .S0(quotient[14]), .Y(n200) );
  MX2X1 U264 ( .A(n155), .B(\u_div/SumTmp[18][6] ), .S0(quotient[18]), .Y(n201) );
  MX2X1 U265 ( .A(n197), .B(\u_div/SumTmp[15][7] ), .S0(quotient[15]), .Y(n202) );
  MX2X1 U266 ( .A(n107), .B(\u_div/SumTmp[19][6] ), .S0(quotient[19]), .Y(n203) );
  MX2X1 U267 ( .A(n199), .B(\u_div/SumTmp[16][7] ), .S0(quotient[16]), .Y(n204) );
  MX2X1 U268 ( .A(n201), .B(\u_div/SumTmp[17][7] ), .S0(quotient[17]), .Y(n205) );
  MX2X1 U269 ( .A(n203), .B(\u_div/SumTmp[18][7] ), .S0(quotient[18]), .Y(n206) );
  MX2X1 U270 ( .A(n174), .B(\u_div/SumTmp[19][7] ), .S0(quotient[19]), .Y(n207) );
  MX2X1 U271 ( .A(n176), .B(\u_div/SumTmp[3][7] ), .S0(quotient[3]), .Y(n208)
         );
  MX2X1 U272 ( .A(n222), .B(\u_div/SumTmp[22][6] ), .S0(quotient[22]), .Y(n209) );
  MX2X1 U273 ( .A(n226), .B(\u_div/SumTmp[22][7] ), .S0(quotient[22]), .Y(n210) );
  MX2X1 U274 ( .A(n161), .B(\u_div/SumTmp[21][6] ), .S0(quotient[21]), .Y(n211) );
  MX2X1 U275 ( .A(n209), .B(\u_div/SumTmp[21][7] ), .S0(quotient[21]), .Y(n212) );
  MX2X1 U276 ( .A(n225), .B(\u_div/SumTmp[24][6] ), .S0(quotient[24]), .Y(n213) );
  MX2X1 U277 ( .A(n228), .B(\u_div/SumTmp[24][7] ), .S0(quotient[24]), .Y(n214) );
  INVX1 U278 ( .A(\u_div/SumTmp[1][9] ), .Y(n274) );
  INVX1 U279 ( .A(\u_div/SumTmp[1][1] ), .Y(n273) );
  INVX1 U280 ( .A(n259), .Y(\u_div/PartRem[23][9] ) );
  NAND2BX1 U281 ( .AN(n300), .B(\u_div/CryTmp[24][8] ), .Y(n303) );
  CLKINVX3 U282 ( .A(n299), .Y(quotient[27]) );
  NAND2BX1 U283 ( .AN(n297), .B(\u_div/CryTmp[27][5] ), .Y(n299) );
  NAND2X1 U284 ( .A(quotient[2]), .B(b[0]), .Y(n257) );
  CLKINVX3 U285 ( .A(n295), .Y(quotient[30]) );
  NAND3BX1 U286 ( .AN(n294), .B(\u_div/BInv [2]), .C(\u_div/CryTmp[30][2] ), 
        .Y(n295) );
  CLKINVX3 U287 ( .A(n298), .Y(quotient[28]) );
  NAND3BX1 U288 ( .AN(n297), .B(\u_div/BInv [4]), .C(\u_div/CryTmp[28][4] ), 
        .Y(n298) );
  XNOR2X1 U289 ( .A(\u_div/CryTmp[3][1] ), .B(a[20]), .Y(\u_div/SumTmp[20][0] ) );
  XNOR2X1 U290 ( .A(\u_div/CryTmp[3][1] ), .B(a[10]), .Y(\u_div/SumTmp[10][0] ) );
  XNOR2X1 U291 ( .A(\u_div/CryTmp[3][1] ), .B(a[9]), .Y(\u_div/SumTmp[9][0] )
         );
  XNOR2X1 U292 ( .A(\u_div/CryTmp[3][1] ), .B(a[8]), .Y(\u_div/SumTmp[8][0] )
         );
  XNOR2X1 U293 ( .A(\u_div/CryTmp[3][1] ), .B(a[7]), .Y(\u_div/SumTmp[7][0] )
         );
  XNOR2X1 U294 ( .A(\u_div/CryTmp[3][1] ), .B(a[6]), .Y(\u_div/SumTmp[6][0] )
         );
  XNOR2X1 U295 ( .A(\u_div/CryTmp[3][1] ), .B(a[11]), .Y(\u_div/SumTmp[11][0] ) );
  XNOR2X1 U296 ( .A(\u_div/CryTmp[3][1] ), .B(a[12]), .Y(\u_div/SumTmp[12][0] ) );
  XNOR2X1 U297 ( .A(\u_div/CryTmp[3][1] ), .B(a[13]), .Y(\u_div/SumTmp[13][0] ) );
  XNOR2X1 U298 ( .A(\u_div/CryTmp[3][1] ), .B(a[5]), .Y(\u_div/SumTmp[5][0] )
         );
  XNOR2X1 U299 ( .A(\u_div/CryTmp[3][1] ), .B(a[14]), .Y(\u_div/SumTmp[14][0] ) );
  XNOR2X1 U300 ( .A(\u_div/CryTmp[3][1] ), .B(a[15]), .Y(\u_div/SumTmp[15][0] ) );
  XNOR2X1 U301 ( .A(\u_div/CryTmp[3][1] ), .B(a[4]), .Y(\u_div/SumTmp[4][0] )
         );
  XNOR2X1 U302 ( .A(\u_div/CryTmp[3][1] ), .B(a[16]), .Y(\u_div/SumTmp[16][0] ) );
  XNOR2X1 U303 ( .A(\u_div/CryTmp[3][1] ), .B(a[17]), .Y(\u_div/SumTmp[17][0] ) );
  XNOR2X1 U304 ( .A(\u_div/CryTmp[3][1] ), .B(a[18]), .Y(\u_div/SumTmp[18][0] ) );
  XNOR2X1 U305 ( .A(\u_div/CryTmp[3][1] ), .B(a[19]), .Y(\u_div/SumTmp[19][0] ) );
  XNOR2X1 U306 ( .A(\u_div/CryTmp[3][1] ), .B(a[22]), .Y(\u_div/SumTmp[22][0] ) );
  XNOR2X1 U307 ( .A(\u_div/CryTmp[3][1] ), .B(a[21]), .Y(\u_div/SumTmp[21][0] ) );
  XNOR2X1 U308 ( .A(\u_div/CryTmp[3][1] ), .B(a[23]), .Y(\u_div/SumTmp[23][0] ) );
  MX2X1 U309 ( .A(n44), .B(\u_div/SumTmp[23][1] ), .S0(quotient[23]), .Y(n215)
         );
  MX2X1 U310 ( .A(n94), .B(\u_div/SumTmp[23][2] ), .S0(quotient[23]), .Y(n216)
         );
  XNOR2X1 U311 ( .A(\u_div/CryTmp[3][1] ), .B(a[24]), .Y(\u_div/SumTmp[24][0] ) );
  XNOR2X1 U312 ( .A(\u_div/CryTmp[3][1] ), .B(a[25]), .Y(\u_div/SumTmp[25][0] ) );
  MX2X1 U313 ( .A(n23), .B(\u_div/SumTmp[25][1] ), .S0(quotient[25]), .Y(n217)
         );
  MX2X1 U314 ( .A(n96), .B(\u_div/SumTmp[25][2] ), .S0(quotient[25]), .Y(n218)
         );
  XNOR2X1 U315 ( .A(\u_div/CryTmp[3][1] ), .B(a[26]), .Y(\u_div/SumTmp[26][0] ) );
  XNOR2X1 U316 ( .A(\u_div/CryTmp[3][1] ), .B(a[27]), .Y(\u_div/SumTmp[27][0] ) );
  XNOR2X1 U317 ( .A(\u_div/CryTmp[3][1] ), .B(a[31]), .Y(\u_div/SumTmp[31][0] ) );
  XNOR2X1 U318 ( .A(\u_div/CryTmp[3][1] ), .B(a[28]), .Y(\u_div/SumTmp[28][0] ) );
  XNOR2X1 U319 ( .A(\u_div/CryTmp[3][1] ), .B(a[29]), .Y(\u_div/SumTmp[29][0] ) );
  XNOR2X1 U320 ( .A(\u_div/CryTmp[3][1] ), .B(a[30]), .Y(\u_div/SumTmp[30][0] ) );
  INVX1 U321 ( .A(n257), .Y(\u_div/PartRem[2][1] ) );
  MXI2X1 U322 ( .A(n257), .B(n273), .S0(quotient[1]), .Y(\u_div/PartRem[1][2] ) );
  NAND2BX1 U323 ( .AN(\u_div/CryTmp[0][10] ), .B(n1), .Y(quotient[0]) );
  CLKINVX3 U324 ( .A(n296), .Y(quotient[29]) );
  NAND2BX1 U325 ( .AN(n294), .B(\u_div/CryTmp[29][3] ), .Y(n296) );
  OR2XL U326 ( .A(a[30]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[30][1] )
         );
  OR2XL U327 ( .A(a[9]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[9][1] ) );
  OR2XL U328 ( .A(a[8]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[8][1] ) );
  OR2XL U329 ( .A(a[7]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[7][1] ) );
  OR2XL U330 ( .A(a[6]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[6][1] ) );
  OR2XL U331 ( .A(a[5]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[5][1] ) );
  OR2XL U332 ( .A(a[10]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[10][1] )
         );
  OR2XL U333 ( .A(a[11]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[11][1] )
         );
  OR2XL U334 ( .A(a[12]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[12][1] )
         );
  OR2XL U335 ( .A(a[4]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[4][1] ) );
  OR2XL U336 ( .A(a[13]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[13][1] )
         );
  OR2XL U337 ( .A(a[14]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[14][1] )
         );
  OR2XL U338 ( .A(a[15]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[15][1] )
         );
  OR2XL U339 ( .A(a[16]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[16][1] )
         );
  OR2XL U340 ( .A(a[17]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[17][1] )
         );
  OR2XL U341 ( .A(a[18]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[18][1] )
         );
  OR2XL U342 ( .A(a[19]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[19][1] )
         );
  OR2XL U343 ( .A(a[20]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[20][1] )
         );
  OR2XL U344 ( .A(a[29]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[29][1] )
         );
  OR2XL U345 ( .A(a[21]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[21][1] )
         );
  OR2XL U346 ( .A(a[22]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[22][1] )
         );
  OR2XL U347 ( .A(a[28]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[28][1] )
         );
  OR2XL U348 ( .A(a[23]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[23][1] )
         );
  OR2XL U349 ( .A(a[24]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[24][1] )
         );
  OR2XL U350 ( .A(a[27]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[27][1] )
         );
  OR2XL U351 ( .A(a[25]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[25][1] )
         );
  OR2XL U352 ( .A(a[26]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[26][1] )
         );
  INVX1 U353 ( .A(n256), .Y(\u_div/PartRem[2][2] ) );
  INVX1 U354 ( .A(n255), .Y(\u_div/PartRem[2][3] ) );
  INVX1 U355 ( .A(n254), .Y(\u_div/PartRem[2][4] ) );
  MXI2X1 U356 ( .A(n255), .B(n271), .S0(quotient[1]), .Y(\u_div/PartRem[1][4] ) );
  INVX1 U357 ( .A(\u_div/SumTmp[1][3] ), .Y(n271) );
  INVX1 U358 ( .A(n253), .Y(\u_div/PartRem[2][5] ) );
  INVX1 U359 ( .A(n252), .Y(\u_div/PartRem[2][6] ) );
  MXI2X1 U360 ( .A(n253), .B(n269), .S0(quotient[1]), .Y(\u_div/PartRem[1][6] ) );
  INVX1 U361 ( .A(\u_div/SumTmp[1][5] ), .Y(n269) );
  INVX1 U362 ( .A(n251), .Y(\u_div/PartRem[2][7] ) );
  INVX1 U363 ( .A(n250), .Y(\u_div/PartRem[2][8] ) );
  MXI2X1 U364 ( .A(n251), .B(n267), .S0(quotient[1]), .Y(\u_div/PartRem[1][8] ) );
  INVX1 U365 ( .A(\u_div/SumTmp[1][7] ), .Y(n267) );
  INVX1 U366 ( .A(n249), .Y(\u_div/PartRem[2][9] ) );
  INVX1 U367 ( .A(n245), .Y(\u_div/PartRem[4][9] ) );
  INVX1 U368 ( .A(n243), .Y(\u_div/PartRem[5][9] ) );
  INVX1 U369 ( .A(n247), .Y(\u_div/PartRem[3][9] ) );
  INVX1 U370 ( .A(n241), .Y(\u_div/PartRem[6][9] ) );
  INVX1 U371 ( .A(n239), .Y(\u_div/PartRem[7][9] ) );
  INVX1 U372 ( .A(n237), .Y(\u_div/PartRem[8][9] ) );
  INVX1 U373 ( .A(n234), .Y(\u_div/PartRem[9][9] ) );
  INVX1 U374 ( .A(n235), .Y(\u_div/PartRem[10][9] ) );
  INVX1 U375 ( .A(n291), .Y(\u_div/PartRem[11][9] ) );
  INVX1 U376 ( .A(n289), .Y(\u_div/PartRem[12][9] ) );
  INVX1 U377 ( .A(n287), .Y(\u_div/PartRem[13][9] ) );
  INVX1 U378 ( .A(n285), .Y(\u_div/PartRem[14][9] ) );
  INVX1 U379 ( .A(n283), .Y(\u_div/PartRem[15][9] ) );
  INVX1 U380 ( .A(n281), .Y(\u_div/PartRem[16][9] ) );
  INVX1 U381 ( .A(n279), .Y(\u_div/PartRem[17][9] ) );
  INVX1 U382 ( .A(n277), .Y(\u_div/PartRem[18][9] ) );
  INVX1 U383 ( .A(n275), .Y(\u_div/PartRem[19][9] ) );
  INVX1 U384 ( .A(n264), .Y(\u_div/PartRem[20][9] ) );
  INVX1 U385 ( .A(n260), .Y(\u_div/PartRem[22][9] ) );
  INVX1 U386 ( .A(n262), .Y(\u_div/PartRem[21][9] ) );
  MX2X1 U387 ( .A(n95), .B(\u_div/SumTmp[23][3] ), .S0(quotient[23]), .Y(n220)
         );
  MX2X1 U388 ( .A(n165), .B(\u_div/SumTmp[23][4] ), .S0(quotient[23]), .Y(n221) );
  MX2X1 U389 ( .A(n166), .B(\u_div/SumTmp[23][5] ), .S0(quotient[23]), .Y(n222) );
  MX2X1 U390 ( .A(n97), .B(\u_div/SumTmp[25][3] ), .S0(quotient[25]), .Y(n223)
         );
  MX2X1 U391 ( .A(n168), .B(\u_div/SumTmp[25][4] ), .S0(quotient[25]), .Y(n224) );
  MX2X1 U392 ( .A(n169), .B(\u_div/SumTmp[25][5] ), .S0(quotient[25]), .Y(n225) );
  MXI2X1 U393 ( .A(n214), .B(\u_div/SumTmp[23][8] ), .S0(quotient[23]), .Y(
        n259) );
  MX2X1 U394 ( .A(n167), .B(\u_div/SumTmp[23][6] ), .S0(quotient[23]), .Y(n226) );
  MX2X1 U395 ( .A(n213), .B(\u_div/SumTmp[23][7] ), .S0(quotient[23]), .Y(n227) );
  MX2X1 U396 ( .A(n170), .B(\u_div/SumTmp[25][6] ), .S0(quotient[25]), .Y(n228) );
  NAND2BX1 U397 ( .AN(b[9]), .B(\u_div/CryTmp[23][9] ), .Y(n304) );
  OR3XL U398 ( .A(b[7]), .B(n300), .C(n302), .Y(n301) );
  INVX1 U399 ( .A(\u_div/CryTmp[25][7] ), .Y(n302) );
  NOR3X1 U400 ( .A(n294), .B(n230), .C(n231), .Y(quotient[31]) );
  OR2X2 U401 ( .A(b[2]), .B(b[1]), .Y(n230) );
  NAND2BX1 U402 ( .AN(b[5]), .B(n232), .Y(n297) );
  OR3X2 U403 ( .A(b[4]), .B(b[3]), .C(n297), .Y(n294) );
  OR2X2 U404 ( .A(b[9]), .B(b[8]), .Y(n300) );
  NOR2X1 U405 ( .A(n300), .B(n233), .Y(n232) );
  OR2X2 U406 ( .A(b[7]), .B(b[6]), .Y(n233) );
  NAND2BX4 U407 ( .AN(\u_div/CryTmp[21][10] ), .B(n51), .Y(quotient[21]) );
  NAND2BX4 U408 ( .AN(\u_div/CryTmp[20][10] ), .B(n21), .Y(quotient[20]) );
  NAND2BX4 U409 ( .AN(\u_div/CryTmp[19][10] ), .B(n3), .Y(quotient[19]) );
  NAND2BX4 U410 ( .AN(\u_div/CryTmp[18][10] ), .B(n4), .Y(quotient[18]) );
  NAND2BX4 U411 ( .AN(\u_div/CryTmp[17][10] ), .B(n5), .Y(quotient[17]) );
  NAND2BX4 U412 ( .AN(\u_div/CryTmp[16][10] ), .B(n6), .Y(quotient[16]) );
  NAND2BX4 U413 ( .AN(\u_div/CryTmp[15][10] ), .B(n7), .Y(quotient[15]) );
  NAND2BX4 U414 ( .AN(\u_div/CryTmp[14][10] ), .B(n8), .Y(quotient[14]) );
  NAND2BX4 U415 ( .AN(\u_div/CryTmp[13][10] ), .B(n9), .Y(quotient[13]) );
  NAND2BX4 U416 ( .AN(\u_div/CryTmp[12][10] ), .B(n10), .Y(quotient[12]) );
  NAND2BX4 U417 ( .AN(\u_div/CryTmp[11][10] ), .B(n11), .Y(quotient[11]) );
  NAND2BX4 U418 ( .AN(\u_div/CryTmp[10][10] ), .B(n12), .Y(quotient[10]) );
  NAND2BX4 U419 ( .AN(\u_div/CryTmp[9][10] ), .B(n13), .Y(quotient[9]) );
  NAND2BX4 U420 ( .AN(\u_div/CryTmp[8][10] ), .B(n14), .Y(quotient[8]) );
  NAND2BX4 U421 ( .AN(\u_div/CryTmp[7][10] ), .B(n15), .Y(quotient[7]) );
  NAND2BX4 U422 ( .AN(\u_div/CryTmp[6][10] ), .B(n16), .Y(quotient[6]) );
  NAND2BX4 U423 ( .AN(\u_div/CryTmp[5][10] ), .B(n17), .Y(quotient[5]) );
  NAND2BX4 U424 ( .AN(\u_div/CryTmp[4][10] ), .B(n18), .Y(quotient[4]) );
  NAND2BX4 U425 ( .AN(\u_div/CryTmp[3][10] ), .B(n19), .Y(quotient[3]) );
  NAND2BX4 U426 ( .AN(\u_div/CryTmp[2][10] ), .B(n20), .Y(quotient[2]) );
  NAND2BX4 U427 ( .AN(\u_div/CryTmp[1][10] ), .B(n2), .Y(quotient[1]) );
  CLKINVX8 U428 ( .A(b[9]), .Y(\u_div/BInv [9]) );
  CLKINVX8 U429 ( .A(b[8]), .Y(\u_div/BInv [8]) );
  CLKINVX8 U430 ( .A(b[7]), .Y(\u_div/BInv [7]) );
  CLKINVX8 U431 ( .A(b[6]), .Y(\u_div/BInv [6]) );
  CLKINVX8 U432 ( .A(b[5]), .Y(\u_div/BInv [5]) );
  CLKINVX8 U433 ( .A(b[3]), .Y(\u_div/BInv [3]) );
  CLKINVX8 U434 ( .A(b[1]), .Y(\u_div/BInv [1]) );
  CLKINVX8 U435 ( .A(b[2]), .Y(\u_div/BInv [2]) );
  CLKINVX8 U436 ( .A(b[4]), .Y(\u_div/BInv [4]) );
endmodule


module Equation_Implementation_DW_div_uns_19 ( a, b, quotient, remainder, 
        divide_by_0 );
  input [31:0] a;
  input [9:0] b;
  output [31:0] quotient;
  output [9:0] remainder;
  output divide_by_0;
  wire   n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, \u_div/SumTmp[2][4] , \u_div/SumTmp[2][5] ,
         \u_div/SumTmp[2][6] , \u_div/SumTmp[2][7] , \u_div/SumTmp[2][8] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[3][4] , \u_div/SumTmp[3][5] ,
         \u_div/SumTmp[3][6] , \u_div/SumTmp[3][7] , \u_div/SumTmp[3][8] ,
         \u_div/SumTmp[4][0] , \u_div/SumTmp[4][4] , \u_div/SumTmp[4][5] ,
         \u_div/SumTmp[4][6] , \u_div/SumTmp[4][7] , \u_div/SumTmp[4][8] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[5][4] , \u_div/SumTmp[5][5] ,
         \u_div/SumTmp[5][6] , \u_div/SumTmp[5][7] , \u_div/SumTmp[5][8] ,
         \u_div/SumTmp[6][0] , \u_div/SumTmp[6][4] , \u_div/SumTmp[6][5] ,
         \u_div/SumTmp[6][6] , \u_div/SumTmp[6][7] , \u_div/SumTmp[6][8] ,
         \u_div/SumTmp[7][0] , \u_div/SumTmp[7][4] , \u_div/SumTmp[7][5] ,
         \u_div/SumTmp[7][6] , \u_div/SumTmp[7][7] , \u_div/SumTmp[7][8] ,
         \u_div/SumTmp[8][0] , \u_div/SumTmp[8][4] , \u_div/SumTmp[8][5] ,
         \u_div/SumTmp[8][6] , \u_div/SumTmp[8][7] , \u_div/SumTmp[8][8] ,
         \u_div/SumTmp[9][0] , \u_div/SumTmp[9][4] , \u_div/SumTmp[9][5] ,
         \u_div/SumTmp[9][6] , \u_div/SumTmp[9][7] , \u_div/SumTmp[9][8] ,
         \u_div/SumTmp[10][0] , \u_div/SumTmp[10][4] , \u_div/SumTmp[10][5] ,
         \u_div/SumTmp[10][6] , \u_div/SumTmp[10][7] , \u_div/SumTmp[10][8] ,
         \u_div/SumTmp[11][0] , \u_div/SumTmp[11][4] , \u_div/SumTmp[11][5] ,
         \u_div/SumTmp[11][6] , \u_div/SumTmp[11][7] , \u_div/SumTmp[11][8] ,
         \u_div/SumTmp[12][0] , \u_div/SumTmp[12][4] , \u_div/SumTmp[12][5] ,
         \u_div/SumTmp[12][6] , \u_div/SumTmp[12][7] , \u_div/SumTmp[12][8] ,
         \u_div/SumTmp[13][0] , \u_div/SumTmp[13][4] , \u_div/SumTmp[13][5] ,
         \u_div/SumTmp[13][6] , \u_div/SumTmp[13][7] , \u_div/SumTmp[13][8] ,
         \u_div/SumTmp[14][0] , \u_div/SumTmp[14][4] , \u_div/SumTmp[14][5] ,
         \u_div/SumTmp[14][6] , \u_div/SumTmp[14][7] , \u_div/SumTmp[14][8] ,
         \u_div/SumTmp[15][0] , \u_div/SumTmp[15][4] , \u_div/SumTmp[15][5] ,
         \u_div/SumTmp[15][6] , \u_div/SumTmp[15][7] , \u_div/SumTmp[15][8] ,
         \u_div/SumTmp[16][0] , \u_div/SumTmp[16][4] , \u_div/SumTmp[16][5] ,
         \u_div/SumTmp[16][6] , \u_div/SumTmp[16][7] , \u_div/SumTmp[16][8] ,
         \u_div/SumTmp[17][0] , \u_div/SumTmp[17][4] , \u_div/SumTmp[17][5] ,
         \u_div/SumTmp[17][6] , \u_div/SumTmp[17][7] , \u_div/SumTmp[17][8] ,
         \u_div/SumTmp[18][0] , \u_div/SumTmp[18][4] , \u_div/SumTmp[18][5] ,
         \u_div/SumTmp[18][6] , \u_div/SumTmp[18][7] , \u_div/SumTmp[18][8] ,
         \u_div/SumTmp[19][0] , \u_div/SumTmp[19][4] , \u_div/SumTmp[19][5] ,
         \u_div/SumTmp[19][6] , \u_div/SumTmp[19][7] , \u_div/SumTmp[19][8] ,
         \u_div/SumTmp[20][0] , \u_div/SumTmp[20][4] , \u_div/SumTmp[20][5] ,
         \u_div/SumTmp[20][6] , \u_div/SumTmp[20][7] , \u_div/SumTmp[20][8] ,
         \u_div/SumTmp[21][0] , \u_div/SumTmp[21][4] , \u_div/SumTmp[21][5] ,
         \u_div/SumTmp[21][6] , \u_div/SumTmp[21][7] , \u_div/SumTmp[21][8] ,
         \u_div/SumTmp[22][0] , \u_div/SumTmp[22][4] , \u_div/SumTmp[22][5] ,
         \u_div/SumTmp[22][6] , \u_div/SumTmp[22][7] , \u_div/SumTmp[22][8] ,
         \u_div/CryTmp[0][4] , \u_div/CryTmp[0][5] , \u_div/CryTmp[1][4] ,
         \u_div/CryTmp[1][5] , \u_div/CryTmp[1][6] , \u_div/CryTmp[1][7] ,
         \u_div/CryTmp[1][8] , \u_div/CryTmp[1][9] , \u_div/CryTmp[1][10] ,
         \u_div/CryTmp[2][4] , \u_div/CryTmp[2][5] , \u_div/CryTmp[2][6] ,
         \u_div/CryTmp[2][7] , \u_div/CryTmp[2][8] , \u_div/CryTmp[2][9] ,
         \u_div/CryTmp[2][10] , \u_div/CryTmp[3][4] , \u_div/CryTmp[3][5] ,
         \u_div/CryTmp[3][6] , \u_div/CryTmp[3][7] , \u_div/CryTmp[3][8] ,
         \u_div/CryTmp[3][9] , \u_div/CryTmp[3][10] , \u_div/CryTmp[4][4] ,
         \u_div/CryTmp[4][5] , \u_div/CryTmp[4][6] , \u_div/CryTmp[4][7] ,
         \u_div/CryTmp[4][8] , \u_div/CryTmp[4][9] , \u_div/CryTmp[4][10] ,
         \u_div/CryTmp[5][4] , \u_div/CryTmp[5][5] , \u_div/CryTmp[5][6] ,
         \u_div/CryTmp[5][7] , \u_div/CryTmp[5][8] , \u_div/CryTmp[5][9] ,
         \u_div/CryTmp[5][10] , \u_div/CryTmp[6][4] , \u_div/CryTmp[6][5] ,
         \u_div/CryTmp[6][6] , \u_div/CryTmp[6][7] , \u_div/CryTmp[6][8] ,
         \u_div/CryTmp[6][9] , \u_div/CryTmp[6][10] , \u_div/CryTmp[7][4] ,
         \u_div/CryTmp[7][5] , \u_div/CryTmp[7][6] , \u_div/CryTmp[7][7] ,
         \u_div/CryTmp[7][8] , \u_div/CryTmp[7][9] , \u_div/CryTmp[7][10] ,
         \u_div/CryTmp[8][4] , \u_div/CryTmp[8][5] , \u_div/CryTmp[8][6] ,
         \u_div/CryTmp[8][7] , \u_div/CryTmp[8][8] , \u_div/CryTmp[8][9] ,
         \u_div/CryTmp[8][10] , \u_div/CryTmp[9][4] , \u_div/CryTmp[9][5] ,
         \u_div/CryTmp[9][6] , \u_div/CryTmp[9][7] , \u_div/CryTmp[9][8] ,
         \u_div/CryTmp[9][9] , \u_div/CryTmp[9][10] , \u_div/CryTmp[10][4] ,
         \u_div/CryTmp[10][5] , \u_div/CryTmp[10][6] , \u_div/CryTmp[10][7] ,
         \u_div/CryTmp[10][8] , \u_div/CryTmp[10][9] , \u_div/CryTmp[10][10] ,
         \u_div/CryTmp[11][4] , \u_div/CryTmp[11][5] , \u_div/CryTmp[11][6] ,
         \u_div/CryTmp[11][7] , \u_div/CryTmp[11][8] , \u_div/CryTmp[11][9] ,
         \u_div/CryTmp[11][10] , \u_div/CryTmp[12][4] , \u_div/CryTmp[12][5] ,
         \u_div/CryTmp[12][6] , \u_div/CryTmp[12][7] , \u_div/CryTmp[12][8] ,
         \u_div/CryTmp[12][9] , \u_div/CryTmp[12][10] , \u_div/CryTmp[13][4] ,
         \u_div/CryTmp[13][5] , \u_div/CryTmp[13][6] , \u_div/CryTmp[13][7] ,
         \u_div/CryTmp[13][8] , \u_div/CryTmp[13][9] , \u_div/CryTmp[13][10] ,
         \u_div/CryTmp[14][4] , \u_div/CryTmp[14][5] , \u_div/CryTmp[14][6] ,
         \u_div/CryTmp[14][7] , \u_div/CryTmp[14][8] , \u_div/CryTmp[14][9] ,
         \u_div/CryTmp[14][10] , \u_div/CryTmp[15][4] , \u_div/CryTmp[15][5] ,
         \u_div/CryTmp[15][6] , \u_div/CryTmp[15][7] , \u_div/CryTmp[15][8] ,
         \u_div/CryTmp[15][9] , \u_div/CryTmp[15][10] , \u_div/CryTmp[16][4] ,
         \u_div/CryTmp[16][5] , \u_div/CryTmp[16][6] , \u_div/CryTmp[16][7] ,
         \u_div/CryTmp[16][8] , \u_div/CryTmp[16][9] , \u_div/CryTmp[16][10] ,
         \u_div/CryTmp[17][4] , \u_div/CryTmp[17][5] , \u_div/CryTmp[17][6] ,
         \u_div/CryTmp[17][7] , \u_div/CryTmp[17][8] , \u_div/CryTmp[17][9] ,
         \u_div/CryTmp[17][10] , \u_div/CryTmp[18][4] , \u_div/CryTmp[18][5] ,
         \u_div/CryTmp[18][6] , \u_div/CryTmp[18][7] , \u_div/CryTmp[18][8] ,
         \u_div/CryTmp[18][9] , \u_div/CryTmp[18][10] , \u_div/CryTmp[19][4] ,
         \u_div/CryTmp[19][5] , \u_div/CryTmp[19][6] , \u_div/CryTmp[19][7] ,
         \u_div/CryTmp[19][8] , \u_div/CryTmp[19][9] , \u_div/CryTmp[19][10] ,
         \u_div/CryTmp[20][4] , \u_div/CryTmp[20][5] , \u_div/CryTmp[20][6] ,
         \u_div/CryTmp[20][7] , \u_div/CryTmp[20][8] , \u_div/CryTmp[20][9] ,
         \u_div/CryTmp[20][10] , \u_div/CryTmp[21][4] , \u_div/CryTmp[21][5] ,
         \u_div/CryTmp[21][6] , \u_div/CryTmp[21][7] , \u_div/CryTmp[21][8] ,
         \u_div/CryTmp[21][9] , \u_div/CryTmp[21][10] , \u_div/CryTmp[22][5] ,
         \u_div/CryTmp[22][6] , \u_div/CryTmp[22][7] , \u_div/CryTmp[22][8] ,
         \u_div/CryTmp[22][9] , \u_div/CryTmp[22][10] , \u_div/PartRem[1][5] ,
         \u_div/PartRem[1][6] , \u_div/PartRem[1][7] , \u_div/PartRem[1][8] ,
         \u_div/PartRem[1][9] , \u_div/PartRem[2][4] , \u_div/PartRem[2][5] ,
         \u_div/PartRem[2][6] , \u_div/PartRem[2][7] , \u_div/PartRem[2][8] ,
         \u_div/PartRem[2][9] , \u_div/PartRem[2][10] , \u_div/PartRem[3][9] ,
         \u_div/PartRem[3][10] , \u_div/PartRem[4][9] , \u_div/PartRem[4][10] ,
         \u_div/PartRem[5][9] , \u_div/PartRem[6][9] , \u_div/PartRem[6][10] ,
         \u_div/PartRem[7][9] , \u_div/PartRem[7][10] , \u_div/PartRem[8][9] ,
         \u_div/PartRem[8][10] , \u_div/PartRem[9][9] , \u_div/PartRem[9][10] ,
         \u_div/PartRem[10][9] , \u_div/PartRem[11][9] ,
         \u_div/PartRem[11][10] , \u_div/PartRem[12][9] ,
         \u_div/PartRem[12][10] , \u_div/PartRem[13][9] ,
         \u_div/PartRem[13][10] , \u_div/PartRem[14][9] ,
         \u_div/PartRem[14][10] , \u_div/PartRem[15][9] ,
         \u_div/PartRem[15][10] , \u_div/PartRem[16][9] ,
         \u_div/PartRem[16][10] , \u_div/PartRem[17][9] ,
         \u_div/PartRem[17][10] , \u_div/PartRem[18][9] ,
         \u_div/PartRem[18][10] , \u_div/PartRem[19][9] ,
         \u_div/PartRem[19][10] , \u_div/PartRem[20][9] ,
         \u_div/PartRem[20][10] , \u_div/PartRem[21][9] ,
         \u_div/PartRem[22][9] , \u_div/PartRem[28][1] ,
         \u_div/PartRem[29][1] , \u_div/PartRem[30][1] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228;
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[12][0]  = a[12];
  assign \u_div/SumTmp[13][0]  = a[13];
  assign \u_div/SumTmp[14][0]  = a[14];
  assign \u_div/SumTmp[15][0]  = a[15];
  assign \u_div/SumTmp[16][0]  = a[16];
  assign \u_div/SumTmp[17][0]  = a[17];
  assign \u_div/SumTmp[18][0]  = a[18];
  assign \u_div/SumTmp[19][0]  = a[19];
  assign \u_div/SumTmp[20][0]  = a[20];
  assign \u_div/SumTmp[21][0]  = a[21];
  assign \u_div/SumTmp[22][0]  = a[22];
  assign \u_div/PartRem[28][1]  = a[28];
  assign \u_div/PartRem[29][1]  = a[29];
  assign \u_div/PartRem[30][1]  = a[30];

  NAND2BX2 U1 ( .AN(\u_div/CryTmp[21][10] ), .B(n159), .Y(n229) );
  NAND2BX2 U2 ( .AN(\u_div/CryTmp[20][10] ), .B(n157), .Y(n230) );
  AND2X2 U3 ( .A(\u_div/CryTmp[19][9] ), .B(\u_div/PartRem[20][9] ), .Y(
        \u_div/CryTmp[19][10] ) );
  AND2X2 U4 ( .A(\u_div/CryTmp[18][9] ), .B(\u_div/PartRem[19][9] ), .Y(
        \u_div/CryTmp[18][10] ) );
  AND2X2 U5 ( .A(\u_div/CryTmp[17][9] ), .B(\u_div/PartRem[18][9] ), .Y(
        \u_div/CryTmp[17][10] ) );
  AND2X2 U6 ( .A(\u_div/CryTmp[16][9] ), .B(\u_div/PartRem[17][9] ), .Y(
        \u_div/CryTmp[16][10] ) );
  AND2X2 U7 ( .A(\u_div/CryTmp[15][9] ), .B(\u_div/PartRem[16][9] ), .Y(
        \u_div/CryTmp[15][10] ) );
  AND2X2 U8 ( .A(\u_div/CryTmp[14][9] ), .B(\u_div/PartRem[15][9] ), .Y(
        \u_div/CryTmp[14][10] ) );
  AND2X2 U9 ( .A(\u_div/CryTmp[13][9] ), .B(\u_div/PartRem[14][9] ), .Y(
        \u_div/CryTmp[13][10] ) );
  AND2X2 U10 ( .A(\u_div/CryTmp[12][9] ), .B(\u_div/PartRem[13][9] ), .Y(
        \u_div/CryTmp[12][10] ) );
  AND2X2 U11 ( .A(\u_div/CryTmp[11][9] ), .B(\u_div/PartRem[12][9] ), .Y(
        \u_div/CryTmp[11][10] ) );
  AND2X2 U12 ( .A(\u_div/CryTmp[10][9] ), .B(\u_div/PartRem[11][9] ), .Y(
        \u_div/CryTmp[10][10] ) );
  AND2X2 U13 ( .A(\u_div/CryTmp[2][9] ), .B(\u_div/PartRem[3][9] ), .Y(
        \u_div/CryTmp[2][10] ) );
  AND2X2 U14 ( .A(\u_div/CryTmp[1][9] ), .B(\u_div/PartRem[2][9] ), .Y(
        \u_div/CryTmp[1][10] ) );
  AND2X2 U15 ( .A(\u_div/CryTmp[3][9] ), .B(\u_div/PartRem[4][9] ), .Y(
        \u_div/CryTmp[3][10] ) );
  NAND2BX2 U16 ( .AN(\u_div/CryTmp[4][10] ), .B(n142), .Y(quotient[4]) );
  AND2X2 U17 ( .A(\u_div/CryTmp[5][9] ), .B(\u_div/PartRem[6][9] ), .Y(
        \u_div/CryTmp[5][10] ) );
  AND2X2 U18 ( .A(\u_div/CryTmp[6][9] ), .B(\u_div/PartRem[7][9] ), .Y(
        \u_div/CryTmp[6][10] ) );
  AND2X2 U19 ( .A(\u_div/CryTmp[7][9] ), .B(\u_div/PartRem[8][9] ), .Y(
        \u_div/CryTmp[7][10] ) );
  AND2X2 U20 ( .A(\u_div/CryTmp[8][9] ), .B(\u_div/PartRem[9][9] ), .Y(
        \u_div/CryTmp[8][10] ) );
  MX2X1 U21 ( .A(a[25]), .B(n210), .S0(\u_div/CryTmp[22][10] ), .Y(n1) );
  MX2X1 U22 ( .A(\u_div/CryTmp[3][4] ), .B(n203), .S0(quotient[3]), .Y(n2) );
  MX2X1 U23 ( .A(\u_div/CryTmp[19][4] ), .B(n216), .S0(n231), .Y(n3) );
  MX2X1 U24 ( .A(\u_div/CryTmp[8][4] ), .B(n195), .S0(quotient[8]), .Y(n4) );
  MX2X1 U25 ( .A(\u_div/CryTmp[20][4] ), .B(n214), .S0(n230), .Y(n5) );
  MX2X1 U26 ( .A(n194), .B(\u_div/CryTmp[1][4] ), .S0(quotient[1]), .Y(n6) );
  AND2X2 U27 ( .A(\u_div/PartRem[1][8] ), .B(n34), .Y(n7) );
  AND2X2 U28 ( .A(\u_div/PartRem[1][6] ), .B(n35), .Y(n8) );
  AND2X2 U29 ( .A(\u_div/PartRem[1][9] ), .B(n7), .Y(n9) );
  MX2X1 U30 ( .A(n98), .B(\u_div/SumTmp[10][7] ), .S0(n240), .Y(n10) );
  MX2X1 U31 ( .A(n93), .B(\u_div/SumTmp[9][7] ), .S0(quotient[9]), .Y(n11) );
  MX2X1 U32 ( .A(n95), .B(\u_div/SumTmp[15][7] ), .S0(n235), .Y(n12) );
  MX2X1 U33 ( .A(n91), .B(\u_div/SumTmp[14][7] ), .S0(n236), .Y(n13) );
  MX2X1 U34 ( .A(n96), .B(\u_div/SumTmp[13][7] ), .S0(n237), .Y(n14) );
  MX2X1 U35 ( .A(n92), .B(\u_div/SumTmp[12][7] ), .S0(n238), .Y(n15) );
  MX2X1 U36 ( .A(n97), .B(\u_div/SumTmp[11][7] ), .S0(n239), .Y(n16) );
  MX2X1 U37 ( .A(n94), .B(\u_div/SumTmp[8][7] ), .S0(quotient[8]), .Y(n17) );
  MX2X1 U38 ( .A(n100), .B(\u_div/SumTmp[7][7] ), .S0(quotient[7]), .Y(n18) );
  MX2X1 U39 ( .A(n101), .B(\u_div/SumTmp[6][7] ), .S0(quotient[6]), .Y(n19) );
  MX2X1 U40 ( .A(n102), .B(\u_div/SumTmp[5][7] ), .S0(quotient[5]), .Y(n20) );
  MX2X1 U41 ( .A(n103), .B(\u_div/SumTmp[4][7] ), .S0(quotient[4]), .Y(n21) );
  MX2X1 U42 ( .A(n105), .B(\u_div/SumTmp[17][7] ), .S0(n233), .Y(n22) );
  MX2X1 U43 ( .A(n99), .B(\u_div/SumTmp[16][7] ), .S0(n234), .Y(n23) );
  MX2X1 U44 ( .A(n104), .B(\u_div/SumTmp[3][7] ), .S0(quotient[3]), .Y(n24) );
  MX2X1 U45 ( .A(n107), .B(\u_div/SumTmp[18][7] ), .S0(n232), .Y(n25) );
  MX2X1 U46 ( .A(n108), .B(\u_div/SumTmp[19][7] ), .S0(n231), .Y(n26) );
  MX2X1 U47 ( .A(n109), .B(\u_div/SumTmp[20][7] ), .S0(n230), .Y(n27) );
  MX2X1 U48 ( .A(n110), .B(\u_div/SumTmp[21][7] ), .S0(n229), .Y(n28) );
  MX2X1 U49 ( .A(a[23]), .B(a[23]), .S0(\u_div/CryTmp[22][10] ), .Y(n29) );
  MX2X1 U50 ( .A(n176), .B(n176), .S0(quotient[5]), .Y(n30) );
  MX2X1 U51 ( .A(n165), .B(n165), .S0(n240), .Y(n31) );
  MX2X1 U52 ( .A(n177), .B(n177), .S0(n229), .Y(n32) );
  MX2X1 U53 ( .A(n133), .B(n133), .S0(quotient[3]), .Y(n33) );
  AND2X2 U54 ( .A(\u_div/PartRem[1][7] ), .B(n8), .Y(n34) );
  AND2X2 U55 ( .A(\u_div/PartRem[1][5] ), .B(\u_div/CryTmp[0][5] ), .Y(n35) );
  MX2X1 U56 ( .A(\u_div/CryTmp[17][4] ), .B(n220), .S0(n233), .Y(n36) );
  MX2X1 U57 ( .A(\u_div/CryTmp[15][4] ), .B(n221), .S0(n235), .Y(n37) );
  MX2X1 U58 ( .A(\u_div/CryTmp[13][4] ), .B(n223), .S0(n237), .Y(n38) );
  MX2X1 U59 ( .A(\u_div/CryTmp[10][4] ), .B(n226), .S0(n240), .Y(n39) );
  MX2X1 U60 ( .A(\u_div/CryTmp[9][4] ), .B(n227), .S0(quotient[9]), .Y(n40) );
  MX2X1 U61 ( .A(\u_div/CryTmp[18][4] ), .B(n218), .S0(n232), .Y(n41) );
  MX2X1 U62 ( .A(\u_div/CryTmp[16][4] ), .B(n228), .S0(n234), .Y(n42) );
  MX2X1 U63 ( .A(\u_div/CryTmp[14][4] ), .B(n222), .S0(n236), .Y(n43) );
  MX2X1 U64 ( .A(\u_div/CryTmp[12][4] ), .B(n224), .S0(n238), .Y(n44) );
  MX2X1 U65 ( .A(\u_div/CryTmp[11][4] ), .B(n225), .S0(n239), .Y(n45) );
  MX2X1 U66 ( .A(\u_div/CryTmp[7][4] ), .B(n205), .S0(quotient[7]), .Y(n46) );
  MX2X1 U67 ( .A(\u_div/CryTmp[6][4] ), .B(n200), .S0(quotient[6]), .Y(n47) );
  MX2X1 U68 ( .A(\u_div/CryTmp[5][4] ), .B(n201), .S0(quotient[5]), .Y(n48) );
  MX2X1 U69 ( .A(\u_div/CryTmp[4][4] ), .B(n202), .S0(quotient[4]), .Y(n49) );
  MX2X1 U70 ( .A(\u_div/CryTmp[21][4] ), .B(n212), .S0(n229), .Y(n50) );
  MX2X1 U71 ( .A(n45), .B(\u_div/SumTmp[10][4] ), .S0(n240), .Y(n51) );
  MX2X1 U72 ( .A(n39), .B(\u_div/SumTmp[9][4] ), .S0(quotient[9]), .Y(n52) );
  MX2X1 U73 ( .A(n3), .B(\u_div/SumTmp[18][4] ), .S0(n232), .Y(n53) );
  MX2X1 U74 ( .A(n41), .B(\u_div/SumTmp[17][4] ), .S0(n233), .Y(n54) );
  MX2X1 U75 ( .A(n36), .B(\u_div/SumTmp[16][4] ), .S0(n234), .Y(n55) );
  MX2X1 U76 ( .A(n42), .B(\u_div/SumTmp[15][4] ), .S0(n235), .Y(n56) );
  MX2X1 U77 ( .A(n37), .B(\u_div/SumTmp[14][4] ), .S0(n236), .Y(n57) );
  MX2X1 U78 ( .A(n43), .B(\u_div/SumTmp[13][4] ), .S0(n237), .Y(n58) );
  MX2X1 U79 ( .A(n38), .B(\u_div/SumTmp[12][4] ), .S0(n238), .Y(n59) );
  MX2X1 U80 ( .A(n44), .B(\u_div/SumTmp[11][4] ), .S0(n239), .Y(n60) );
  MX2X1 U81 ( .A(n40), .B(\u_div/SumTmp[8][4] ), .S0(quotient[8]), .Y(n61) );
  MX2X1 U82 ( .A(n4), .B(\u_div/SumTmp[7][4] ), .S0(quotient[7]), .Y(n62) );
  MX2X1 U83 ( .A(n46), .B(\u_div/SumTmp[6][4] ), .S0(quotient[6]), .Y(n63) );
  MX2X1 U84 ( .A(n47), .B(\u_div/SumTmp[5][4] ), .S0(quotient[5]), .Y(n64) );
  MX2X1 U85 ( .A(n48), .B(\u_div/SumTmp[4][4] ), .S0(quotient[4]), .Y(n65) );
  MX2X1 U86 ( .A(n50), .B(\u_div/SumTmp[20][4] ), .S0(n230), .Y(n66) );
  MX2X1 U87 ( .A(n5), .B(\u_div/SumTmp[19][4] ), .S0(n231), .Y(n67) );
  MX2X1 U88 ( .A(n49), .B(\u_div/SumTmp[3][4] ), .S0(quotient[3]), .Y(n68) );
  MX2X1 U89 ( .A(n1), .B(\u_div/SumTmp[21][4] ), .S0(n229), .Y(n69) );
  MX2X1 U90 ( .A(a[26]), .B(\u_div/SumTmp[22][4] ), .S0(\u_div/CryTmp[22][10] ), .Y(n70) );
  MX2X1 U91 ( .A(n55), .B(\u_div/SumTmp[15][5] ), .S0(n235), .Y(n71) );
  MX2X1 U92 ( .A(n56), .B(\u_div/SumTmp[14][5] ), .S0(n236), .Y(n72) );
  MX2X1 U93 ( .A(n57), .B(\u_div/SumTmp[13][5] ), .S0(n237), .Y(n73) );
  MX2X1 U94 ( .A(n58), .B(\u_div/SumTmp[12][5] ), .S0(n238), .Y(n74) );
  MX2X1 U95 ( .A(n60), .B(\u_div/SumTmp[10][5] ), .S0(n240), .Y(n75) );
  MX2X1 U96 ( .A(n51), .B(\u_div/SumTmp[9][5] ), .S0(quotient[9]), .Y(n76) );
  MX2X1 U97 ( .A(n59), .B(\u_div/SumTmp[11][5] ), .S0(n239), .Y(n77) );
  MX2X1 U98 ( .A(n53), .B(\u_div/SumTmp[17][5] ), .S0(n233), .Y(n78) );
  MX2X1 U99 ( .A(n54), .B(\u_div/SumTmp[16][5] ), .S0(n234), .Y(n79) );
  MX2X1 U100 ( .A(n52), .B(\u_div/SumTmp[8][5] ), .S0(quotient[8]), .Y(n80) );
  MX2X1 U101 ( .A(n61), .B(\u_div/SumTmp[7][5] ), .S0(quotient[7]), .Y(n81) );
  MX2X1 U102 ( .A(n62), .B(\u_div/SumTmp[6][5] ), .S0(quotient[6]), .Y(n82) );
  MX2X1 U103 ( .A(n63), .B(\u_div/SumTmp[5][5] ), .S0(quotient[5]), .Y(n83) );
  MX2X1 U104 ( .A(n64), .B(\u_div/SumTmp[4][5] ), .S0(quotient[4]), .Y(n84) );
  MX2X1 U105 ( .A(n66), .B(\u_div/SumTmp[19][5] ), .S0(n231), .Y(n85) );
  MX2X1 U106 ( .A(n67), .B(\u_div/SumTmp[18][5] ), .S0(n232), .Y(n86) );
  MX2X1 U107 ( .A(n65), .B(\u_div/SumTmp[3][5] ), .S0(quotient[3]), .Y(n87) );
  MX2X1 U108 ( .A(n70), .B(\u_div/SumTmp[21][5] ), .S0(n229), .Y(n88) );
  MX2X1 U109 ( .A(n69), .B(\u_div/SumTmp[20][5] ), .S0(n230), .Y(n89) );
  MX2X1 U110 ( .A(a[27]), .B(\u_div/SumTmp[22][5] ), .S0(
        \u_div/CryTmp[22][10] ), .Y(n90) );
  MX2X1 U111 ( .A(n79), .B(\u_div/SumTmp[15][6] ), .S0(n235), .Y(n91) );
  MX2X1 U112 ( .A(n72), .B(\u_div/SumTmp[13][6] ), .S0(n237), .Y(n92) );
  MX2X1 U113 ( .A(n77), .B(\u_div/SumTmp[10][6] ), .S0(n240), .Y(n93) );
  MX2X1 U114 ( .A(n75), .B(\u_div/SumTmp[9][6] ), .S0(quotient[9]), .Y(n94) );
  MX2X1 U115 ( .A(n78), .B(\u_div/SumTmp[16][6] ), .S0(n234), .Y(n95) );
  MX2X1 U116 ( .A(n71), .B(\u_div/SumTmp[14][6] ), .S0(n236), .Y(n96) );
  MX2X1 U117 ( .A(n73), .B(\u_div/SumTmp[12][6] ), .S0(n238), .Y(n97) );
  MX2X1 U118 ( .A(n74), .B(\u_div/SumTmp[11][6] ), .S0(n239), .Y(n98) );
  MX2X1 U119 ( .A(n86), .B(\u_div/SumTmp[17][6] ), .S0(n233), .Y(n99) );
  MX2X1 U120 ( .A(n76), .B(\u_div/SumTmp[8][6] ), .S0(quotient[8]), .Y(n100)
         );
  MX2X1 U121 ( .A(n80), .B(\u_div/SumTmp[7][6] ), .S0(quotient[7]), .Y(n101)
         );
  MX2X1 U122 ( .A(n81), .B(\u_div/SumTmp[6][6] ), .S0(quotient[6]), .Y(n102)
         );
  MX2X1 U123 ( .A(n82), .B(\u_div/SumTmp[5][6] ), .S0(quotient[5]), .Y(n103)
         );
  MX2X1 U124 ( .A(n83), .B(\u_div/SumTmp[4][6] ), .S0(quotient[4]), .Y(n104)
         );
  MX2X1 U125 ( .A(n85), .B(\u_div/SumTmp[18][6] ), .S0(n232), .Y(n105) );
  MX2X1 U126 ( .A(n84), .B(\u_div/SumTmp[3][6] ), .S0(quotient[3]), .Y(n106)
         );
  MX2X1 U127 ( .A(n89), .B(\u_div/SumTmp[19][6] ), .S0(n231), .Y(n107) );
  MX2X1 U128 ( .A(n88), .B(\u_div/SumTmp[20][6] ), .S0(n230), .Y(n108) );
  MX2X1 U129 ( .A(n90), .B(\u_div/SumTmp[21][6] ), .S0(n229), .Y(n109) );
  MX2X1 U130 ( .A(\u_div/PartRem[28][1] ), .B(\u_div/SumTmp[22][6] ), .S0(
        \u_div/CryTmp[22][10] ), .Y(n110) );
  MX2X1 U131 ( .A(\u_div/PartRem[29][1] ), .B(\u_div/SumTmp[22][7] ), .S0(
        \u_div/CryTmp[22][10] ), .Y(n111) );
  MX2X1 U132 ( .A(n188), .B(n152), .S0(quotient[1]), .Y(n112) );
  XOR2X1 U133 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/CryTmp[1][4] ), .Y(n113)
         );
  XNOR2X1 U134 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/CryTmp[1][5] ), .Y(n114)
         );
  MX2X1 U135 ( .A(n173), .B(n173), .S0(quotient[8]), .Y(n115) );
  MX2X1 U136 ( .A(n174), .B(n174), .S0(quotient[7]), .Y(n116) );
  MX2X1 U137 ( .A(n175), .B(n175), .S0(quotient[6]), .Y(n117) );
  MX2X1 U138 ( .A(n168), .B(n168), .S0(n231), .Y(n118) );
  MX2X1 U139 ( .A(n169), .B(n169), .S0(n232), .Y(n119) );
  MX2X1 U140 ( .A(n166), .B(n166), .S0(n233), .Y(n120) );
  MX2X1 U141 ( .A(n170), .B(n170), .S0(n234), .Y(n121) );
  MX2X1 U142 ( .A(n160), .B(n160), .S0(n235), .Y(n122) );
  MX2X1 U143 ( .A(n163), .B(n163), .S0(n236), .Y(n123) );
  MX2X1 U144 ( .A(n161), .B(n161), .S0(n237), .Y(n124) );
  MX2X1 U145 ( .A(n164), .B(n164), .S0(n238), .Y(n125) );
  MX2X1 U146 ( .A(n162), .B(n162), .S0(n239), .Y(n126) );
  MX2X1 U147 ( .A(n172), .B(n172), .S0(quotient[9]), .Y(n127) );
  MX2X1 U148 ( .A(n179), .B(n179), .S0(quotient[4]), .Y(n128) );
  MX2X1 U149 ( .A(n167), .B(n167), .S0(n230), .Y(n129) );
  XNOR2X1 U150 ( .A(\u_div/PartRem[2][8] ), .B(\u_div/CryTmp[1][8] ), .Y(n130)
         );
  XNOR2X1 U151 ( .A(\u_div/PartRem[2][7] ), .B(\u_div/CryTmp[1][7] ), .Y(n131)
         );
  XNOR2X1 U152 ( .A(\u_div/PartRem[2][6] ), .B(\u_div/CryTmp[1][6] ), .Y(n132)
         );
  MX2X1 U153 ( .A(\u_div/SumTmp[4][0] ), .B(\u_div/SumTmp[4][0] ), .S0(
        quotient[4]), .Y(n133) );
  AND2X2 U154 ( .A(\u_div/CryTmp[9][9] ), .B(\u_div/PartRem[10][9] ), .Y(
        \u_div/CryTmp[9][10] ) );
  AND2X2 U155 ( .A(\u_div/CryTmp[4][9] ), .B(\u_div/PartRem[5][9] ), .Y(
        \u_div/CryTmp[4][10] ) );
  AND2X2 U156 ( .A(\u_div/CryTmp[20][9] ), .B(\u_div/PartRem[21][9] ), .Y(
        \u_div/CryTmp[20][10] ) );
  AND2X2 U157 ( .A(\u_div/CryTmp[21][9] ), .B(\u_div/PartRem[22][9] ), .Y(
        \u_div/CryTmp[21][10] ) );
  OR2X2 U158 ( .A(\u_div/CryTmp[8][10] ), .B(\u_div/PartRem[9][10] ), .Y(
        quotient[8]) );
  MXI2X1 U159 ( .A(n181), .B(n141), .S0(quotient[9]), .Y(
        \u_div/PartRem[9][10] ) );
  OR2X2 U160 ( .A(\u_div/CryTmp[12][10] ), .B(\u_div/PartRem[13][10] ), .Y(
        n238) );
  MXI2X1 U161 ( .A(n213), .B(n137), .S0(n237), .Y(\u_div/PartRem[13][10] ) );
  OR2X2 U162 ( .A(\u_div/CryTmp[10][10] ), .B(\u_div/PartRem[11][10] ), .Y(
        n240) );
  MXI2X1 U163 ( .A(n217), .B(n139), .S0(n239), .Y(\u_div/PartRem[11][10] ) );
  OR2X2 U164 ( .A(\u_div/CryTmp[11][10] ), .B(\u_div/PartRem[12][10] ), .Y(
        n239) );
  MXI2X1 U165 ( .A(n215), .B(n138), .S0(n238), .Y(\u_div/PartRem[12][10] ) );
  MX2X1 U166 ( .A(n219), .B(n140), .S0(n240), .Y(n134) );
  INVX1 U167 ( .A(n180), .Y(\u_div/PartRem[9][9] ) );
  INVX1 U168 ( .A(n182), .Y(\u_div/PartRem[8][9] ) );
  INVX1 U169 ( .A(n213), .Y(\u_div/PartRem[14][9] ) );
  INVX1 U170 ( .A(n215), .Y(\u_div/PartRem[13][9] ) );
  INVX1 U171 ( .A(n217), .Y(\u_div/PartRem[12][9] ) );
  INVX1 U172 ( .A(n219), .Y(\u_div/PartRem[11][9] ) );
  INVX1 U173 ( .A(n181), .Y(\u_div/PartRem[10][9] ) );
  XNOR2X1 U174 ( .A(\u_div/PartRem[9][9] ), .B(\u_div/CryTmp[8][9] ), .Y(n135)
         );
  XNOR2X1 U175 ( .A(\u_div/PartRem[15][9] ), .B(\u_div/CryTmp[14][9] ), .Y(
        n136) );
  XNOR2X1 U176 ( .A(\u_div/PartRem[14][9] ), .B(\u_div/CryTmp[13][9] ), .Y(
        n137) );
  XNOR2X1 U177 ( .A(\u_div/PartRem[13][9] ), .B(\u_div/CryTmp[12][9] ), .Y(
        n138) );
  XNOR2X1 U178 ( .A(\u_div/PartRem[12][9] ), .B(\u_div/CryTmp[11][9] ), .Y(
        n139) );
  XNOR2X1 U179 ( .A(\u_div/PartRem[11][9] ), .B(\u_div/CryTmp[10][9] ), .Y(
        n140) );
  XNOR2X1 U180 ( .A(\u_div/PartRem[10][9] ), .B(\u_div/CryTmp[9][9] ), .Y(n141) );
  OR2X2 U181 ( .A(\u_div/CryTmp[7][10] ), .B(\u_div/PartRem[8][10] ), .Y(
        quotient[7]) );
  MXI2X1 U182 ( .A(n180), .B(n135), .S0(quotient[8]), .Y(
        \u_div/PartRem[8][10] ) );
  OR2X2 U183 ( .A(\u_div/CryTmp[6][10] ), .B(\u_div/PartRem[7][10] ), .Y(
        quotient[6]) );
  MXI2X1 U184 ( .A(n182), .B(n143), .S0(quotient[7]), .Y(
        \u_div/PartRem[7][10] ) );
  OR2X2 U185 ( .A(\u_div/CryTmp[5][10] ), .B(\u_div/PartRem[6][10] ), .Y(
        quotient[5]) );
  MXI2X1 U186 ( .A(n183), .B(n144), .S0(quotient[6]), .Y(
        \u_div/PartRem[6][10] ) );
  MX2X1 U187 ( .A(n184), .B(n145), .S0(quotient[5]), .Y(n142) );
  OR2X2 U188 ( .A(\u_div/CryTmp[14][10] ), .B(\u_div/PartRem[15][10] ), .Y(
        n236) );
  MXI2X1 U189 ( .A(n209), .B(n149), .S0(n235), .Y(\u_div/PartRem[15][10] ) );
  OR2X2 U190 ( .A(\u_div/CryTmp[13][10] ), .B(\u_div/PartRem[14][10] ), .Y(
        n237) );
  MXI2X1 U191 ( .A(n211), .B(n136), .S0(n236), .Y(\u_div/PartRem[14][10] ) );
  AND2X2 U192 ( .A(\u_div/CryTmp[14][8] ), .B(n12), .Y(\u_div/CryTmp[14][9] )
         );
  AND2X2 U193 ( .A(\u_div/CryTmp[13][8] ), .B(n13), .Y(\u_div/CryTmp[13][9] )
         );
  AND2X2 U194 ( .A(\u_div/CryTmp[12][8] ), .B(n14), .Y(\u_div/CryTmp[12][9] )
         );
  AND2X2 U195 ( .A(\u_div/CryTmp[11][8] ), .B(n15), .Y(\u_div/CryTmp[11][9] )
         );
  AND2X2 U196 ( .A(\u_div/CryTmp[10][8] ), .B(n16), .Y(\u_div/CryTmp[10][9] )
         );
  AND2X2 U197 ( .A(\u_div/CryTmp[9][8] ), .B(n10), .Y(\u_div/CryTmp[9][9] ) );
  AND2X2 U198 ( .A(\u_div/CryTmp[8][8] ), .B(n11), .Y(\u_div/CryTmp[8][9] ) );
  OR2X2 U199 ( .A(\u_div/CryTmp[3][10] ), .B(\u_div/PartRem[4][10] ), .Y(
        quotient[3]) );
  MXI2X1 U200 ( .A(n185), .B(n146), .S0(quotient[4]), .Y(
        \u_div/PartRem[4][10] ) );
  MXI2X1 U201 ( .A(n10), .B(\u_div/SumTmp[9][8] ), .S0(quotient[9]), .Y(n180)
         );
  XOR2X1 U202 ( .A(n10), .B(\u_div/CryTmp[9][8] ), .Y(\u_div/SumTmp[9][8] ) );
  MXI2X1 U203 ( .A(n11), .B(\u_div/SumTmp[8][8] ), .S0(quotient[8]), .Y(n182)
         );
  XOR2X1 U204 ( .A(n11), .B(\u_div/CryTmp[8][8] ), .Y(\u_div/SumTmp[8][8] ) );
  MXI2X1 U205 ( .A(n12), .B(\u_div/SumTmp[14][8] ), .S0(n236), .Y(n213) );
  XOR2X1 U206 ( .A(n12), .B(\u_div/CryTmp[14][8] ), .Y(\u_div/SumTmp[14][8] )
         );
  MXI2X1 U207 ( .A(n13), .B(\u_div/SumTmp[13][8] ), .S0(n237), .Y(n215) );
  XOR2X1 U208 ( .A(n13), .B(\u_div/CryTmp[13][8] ), .Y(\u_div/SumTmp[13][8] )
         );
  MXI2X1 U209 ( .A(n14), .B(\u_div/SumTmp[12][8] ), .S0(n238), .Y(n217) );
  XOR2X1 U210 ( .A(n14), .B(\u_div/CryTmp[12][8] ), .Y(\u_div/SumTmp[12][8] )
         );
  MXI2X1 U211 ( .A(n15), .B(\u_div/SumTmp[11][8] ), .S0(n239), .Y(n219) );
  XOR2X1 U212 ( .A(n15), .B(\u_div/CryTmp[11][8] ), .Y(\u_div/SumTmp[11][8] )
         );
  MXI2X1 U213 ( .A(n16), .B(\u_div/SumTmp[10][8] ), .S0(n240), .Y(n181) );
  XOR2X1 U214 ( .A(n16), .B(\u_div/CryTmp[10][8] ), .Y(\u_div/SumTmp[10][8] )
         );
  INVX1 U215 ( .A(n183), .Y(\u_div/PartRem[7][9] ) );
  INVX1 U216 ( .A(n184), .Y(\u_div/PartRem[6][9] ) );
  INVX1 U217 ( .A(n185), .Y(\u_div/PartRem[5][9] ) );
  INVX1 U218 ( .A(n186), .Y(\u_div/PartRem[4][9] ) );
  INVX1 U219 ( .A(n187), .Y(\u_div/PartRem[3][9] ) );
  INVX1 U220 ( .A(n209), .Y(\u_div/PartRem[16][9] ) );
  INVX1 U221 ( .A(n211), .Y(\u_div/PartRem[15][9] ) );
  XNOR2X1 U222 ( .A(\u_div/PartRem[8][9] ), .B(\u_div/CryTmp[7][9] ), .Y(n143)
         );
  XNOR2X1 U223 ( .A(\u_div/PartRem[7][9] ), .B(\u_div/CryTmp[6][9] ), .Y(n144)
         );
  XNOR2X1 U224 ( .A(\u_div/PartRem[6][9] ), .B(\u_div/CryTmp[5][9] ), .Y(n145)
         );
  XNOR2X1 U225 ( .A(\u_div/PartRem[5][9] ), .B(\u_div/CryTmp[4][9] ), .Y(n146)
         );
  XNOR2X1 U226 ( .A(\u_div/PartRem[4][9] ), .B(\u_div/CryTmp[3][9] ), .Y(n147)
         );
  XNOR2X1 U227 ( .A(\u_div/PartRem[17][9] ), .B(\u_div/CryTmp[16][9] ), .Y(
        n148) );
  XNOR2X1 U228 ( .A(\u_div/PartRem[16][9] ), .B(\u_div/CryTmp[15][9] ), .Y(
        n149) );
  OR2X2 U229 ( .A(\u_div/CryTmp[2][10] ), .B(\u_div/PartRem[3][10] ), .Y(
        quotient[2]) );
  MXI2X1 U230 ( .A(n186), .B(n147), .S0(quotient[3]), .Y(
        \u_div/PartRem[3][10] ) );
  OR2X2 U231 ( .A(\u_div/CryTmp[16][10] ), .B(\u_div/PartRem[17][10] ), .Y(
        n234) );
  MXI2X1 U232 ( .A(n207), .B(n151), .S0(n233), .Y(\u_div/PartRem[17][10] ) );
  OR2X2 U233 ( .A(\u_div/CryTmp[15][10] ), .B(\u_div/PartRem[16][10] ), .Y(
        n235) );
  MXI2X1 U234 ( .A(n208), .B(n148), .S0(n234), .Y(\u_div/PartRem[16][10] ) );
  OR2X2 U235 ( .A(\u_div/CryTmp[1][10] ), .B(\u_div/PartRem[2][10] ), .Y(
        quotient[1]) );
  MXI2X1 U236 ( .A(n187), .B(n150), .S0(quotient[2]), .Y(
        \u_div/PartRem[2][10] ) );
  AND2X2 U237 ( .A(\u_div/CryTmp[16][8] ), .B(n22), .Y(\u_div/CryTmp[16][9] )
         );
  AND2X2 U238 ( .A(\u_div/CryTmp[15][7] ), .B(n95), .Y(\u_div/CryTmp[15][8] )
         );
  AND2X2 U239 ( .A(\u_div/CryTmp[15][8] ), .B(n23), .Y(\u_div/CryTmp[15][9] )
         );
  AND2X2 U240 ( .A(\u_div/CryTmp[14][7] ), .B(n91), .Y(\u_div/CryTmp[14][8] )
         );
  AND2X2 U241 ( .A(\u_div/CryTmp[13][7] ), .B(n96), .Y(\u_div/CryTmp[13][8] )
         );
  AND2X2 U242 ( .A(\u_div/CryTmp[12][7] ), .B(n92), .Y(\u_div/CryTmp[12][8] )
         );
  AND2X2 U243 ( .A(\u_div/CryTmp[11][7] ), .B(n97), .Y(\u_div/CryTmp[11][8] )
         );
  AND2X2 U244 ( .A(\u_div/CryTmp[10][7] ), .B(n98), .Y(\u_div/CryTmp[10][8] )
         );
  AND2X2 U245 ( .A(\u_div/CryTmp[9][7] ), .B(n93), .Y(\u_div/CryTmp[9][8] ) );
  AND2X2 U246 ( .A(\u_div/CryTmp[8][7] ), .B(n94), .Y(\u_div/CryTmp[8][8] ) );
  AND2X2 U247 ( .A(\u_div/CryTmp[7][8] ), .B(n17), .Y(\u_div/CryTmp[7][9] ) );
  AND2X2 U248 ( .A(\u_div/CryTmp[6][8] ), .B(n18), .Y(\u_div/CryTmp[6][9] ) );
  AND2X2 U249 ( .A(\u_div/CryTmp[5][8] ), .B(n19), .Y(\u_div/CryTmp[5][9] ) );
  AND2X2 U250 ( .A(\u_div/CryTmp[4][8] ), .B(n20), .Y(\u_div/CryTmp[4][9] ) );
  AND2X2 U251 ( .A(\u_div/CryTmp[3][8] ), .B(n21), .Y(\u_div/CryTmp[3][9] ) );
  NAND2BX1 U252 ( .AN(n9), .B(n112), .Y(quotient[0]) );
  MXI2X1 U253 ( .A(n17), .B(\u_div/SumTmp[7][8] ), .S0(quotient[7]), .Y(n183)
         );
  XOR2X1 U254 ( .A(n17), .B(\u_div/CryTmp[7][8] ), .Y(\u_div/SumTmp[7][8] ) );
  MXI2X1 U255 ( .A(n18), .B(\u_div/SumTmp[6][8] ), .S0(quotient[6]), .Y(n184)
         );
  XOR2X1 U256 ( .A(n18), .B(\u_div/CryTmp[6][8] ), .Y(\u_div/SumTmp[6][8] ) );
  MXI2X1 U257 ( .A(n19), .B(\u_div/SumTmp[5][8] ), .S0(quotient[5]), .Y(n185)
         );
  XOR2X1 U258 ( .A(n19), .B(\u_div/CryTmp[5][8] ), .Y(\u_div/SumTmp[5][8] ) );
  MXI2X1 U259 ( .A(n20), .B(\u_div/SumTmp[4][8] ), .S0(quotient[4]), .Y(n186)
         );
  XOR2X1 U260 ( .A(n20), .B(\u_div/CryTmp[4][8] ), .Y(\u_div/SumTmp[4][8] ) );
  MXI2X1 U261 ( .A(n21), .B(\u_div/SumTmp[3][8] ), .S0(quotient[3]), .Y(n187)
         );
  XOR2X1 U262 ( .A(n21), .B(\u_div/CryTmp[3][8] ), .Y(\u_div/SumTmp[3][8] ) );
  MXI2X1 U263 ( .A(n22), .B(\u_div/SumTmp[16][8] ), .S0(n234), .Y(n209) );
  XOR2X1 U264 ( .A(n22), .B(\u_div/CryTmp[16][8] ), .Y(\u_div/SumTmp[16][8] )
         );
  MXI2X1 U265 ( .A(n23), .B(\u_div/SumTmp[15][8] ), .S0(n235), .Y(n211) );
  XOR2X1 U266 ( .A(n23), .B(\u_div/CryTmp[15][8] ), .Y(\u_div/SumTmp[15][8] )
         );
  XOR2X1 U267 ( .A(n91), .B(\u_div/CryTmp[14][7] ), .Y(\u_div/SumTmp[14][7] )
         );
  XOR2X1 U268 ( .A(n92), .B(\u_div/CryTmp[12][7] ), .Y(\u_div/SumTmp[12][7] )
         );
  XOR2X1 U269 ( .A(n93), .B(\u_div/CryTmp[9][7] ), .Y(\u_div/SumTmp[9][7] ) );
  XOR2X1 U270 ( .A(n94), .B(\u_div/CryTmp[8][7] ), .Y(\u_div/SumTmp[8][7] ) );
  XOR2X1 U271 ( .A(n95), .B(\u_div/CryTmp[15][7] ), .Y(\u_div/SumTmp[15][7] )
         );
  XOR2X1 U272 ( .A(n96), .B(\u_div/CryTmp[13][7] ), .Y(\u_div/SumTmp[13][7] )
         );
  XOR2X1 U273 ( .A(n97), .B(\u_div/CryTmp[11][7] ), .Y(\u_div/SumTmp[11][7] )
         );
  XOR2X1 U274 ( .A(n98), .B(\u_div/CryTmp[10][7] ), .Y(\u_div/SumTmp[10][7] )
         );
  INVX1 U275 ( .A(n188), .Y(\u_div/PartRem[2][9] ) );
  INVX1 U276 ( .A(n208), .Y(\u_div/PartRem[17][9] ) );
  INVX1 U277 ( .A(n207), .Y(\u_div/PartRem[18][9] ) );
  XNOR2X1 U278 ( .A(\u_div/PartRem[3][9] ), .B(\u_div/CryTmp[2][9] ), .Y(n150)
         );
  XNOR2X1 U279 ( .A(\u_div/PartRem[18][9] ), .B(\u_div/CryTmp[17][9] ), .Y(
        n151) );
  XNOR2X1 U280 ( .A(\u_div/PartRem[2][9] ), .B(\u_div/CryTmp[1][9] ), .Y(n152)
         );
  XNOR2X1 U281 ( .A(\u_div/PartRem[19][9] ), .B(\u_div/CryTmp[18][9] ), .Y(
        n153) );
  OR2X2 U282 ( .A(\u_div/CryTmp[17][10] ), .B(\u_div/PartRem[18][10] ), .Y(
        n233) );
  MXI2X1 U283 ( .A(n206), .B(n153), .S0(n232), .Y(\u_div/PartRem[18][10] ) );
  AND2X2 U284 ( .A(\u_div/CryTmp[17][7] ), .B(n105), .Y(\u_div/CryTmp[17][8] )
         );
  AND2X2 U285 ( .A(\u_div/CryTmp[17][8] ), .B(n25), .Y(\u_div/CryTmp[17][9] )
         );
  AND2X2 U286 ( .A(\u_div/CryTmp[16][6] ), .B(n78), .Y(\u_div/CryTmp[16][7] )
         );
  AND2X2 U287 ( .A(\u_div/CryTmp[16][7] ), .B(n99), .Y(\u_div/CryTmp[16][8] )
         );
  AND2X2 U288 ( .A(\u_div/CryTmp[15][6] ), .B(n79), .Y(\u_div/CryTmp[15][7] )
         );
  AND2X2 U289 ( .A(\u_div/CryTmp[14][6] ), .B(n71), .Y(\u_div/CryTmp[14][7] )
         );
  AND2X2 U290 ( .A(\u_div/CryTmp[13][6] ), .B(n72), .Y(\u_div/CryTmp[13][7] )
         );
  AND2X2 U291 ( .A(\u_div/CryTmp[12][6] ), .B(n73), .Y(\u_div/CryTmp[12][7] )
         );
  AND2X2 U292 ( .A(\u_div/CryTmp[11][6] ), .B(n74), .Y(\u_div/CryTmp[11][7] )
         );
  AND2X2 U293 ( .A(\u_div/CryTmp[10][6] ), .B(n77), .Y(\u_div/CryTmp[10][7] )
         );
  AND2X2 U294 ( .A(\u_div/CryTmp[9][6] ), .B(n75), .Y(\u_div/CryTmp[9][7] ) );
  AND2X2 U295 ( .A(\u_div/CryTmp[8][6] ), .B(n76), .Y(\u_div/CryTmp[8][7] ) );
  AND2X2 U296 ( .A(\u_div/CryTmp[7][7] ), .B(n100), .Y(\u_div/CryTmp[7][8] )
         );
  AND2X2 U297 ( .A(\u_div/CryTmp[6][7] ), .B(n101), .Y(\u_div/CryTmp[6][8] )
         );
  AND2X2 U298 ( .A(\u_div/CryTmp[5][7] ), .B(n102), .Y(\u_div/CryTmp[5][8] )
         );
  AND2X2 U299 ( .A(\u_div/CryTmp[4][7] ), .B(n103), .Y(\u_div/CryTmp[4][8] )
         );
  AND2X2 U300 ( .A(\u_div/CryTmp[3][7] ), .B(n104), .Y(\u_div/CryTmp[3][8] )
         );
  AND2X2 U301 ( .A(\u_div/CryTmp[2][8] ), .B(n24), .Y(\u_div/CryTmp[2][9] ) );
  AND2X2 U302 ( .A(\u_div/CryTmp[1][8] ), .B(\u_div/PartRem[2][8] ), .Y(
        \u_div/CryTmp[1][9] ) );
  XOR2X1 U303 ( .A(n71), .B(\u_div/CryTmp[14][6] ), .Y(\u_div/SumTmp[14][6] )
         );
  XOR2X1 U304 ( .A(n72), .B(\u_div/CryTmp[13][6] ), .Y(\u_div/SumTmp[13][6] )
         );
  XOR2X1 U305 ( .A(n73), .B(\u_div/CryTmp[12][6] ), .Y(\u_div/SumTmp[12][6] )
         );
  XOR2X1 U306 ( .A(n74), .B(\u_div/CryTmp[11][6] ), .Y(\u_div/SumTmp[11][6] )
         );
  XOR2X1 U307 ( .A(n75), .B(\u_div/CryTmp[9][6] ), .Y(\u_div/SumTmp[9][6] ) );
  XOR2X1 U308 ( .A(n76), .B(\u_div/CryTmp[8][6] ), .Y(\u_div/SumTmp[8][6] ) );
  XOR2X1 U309 ( .A(n77), .B(\u_div/CryTmp[10][6] ), .Y(\u_div/SumTmp[10][6] )
         );
  AND2X2 U310 ( .A(\u_div/CryTmp[18][8] ), .B(n26), .Y(\u_div/CryTmp[18][9] )
         );
  MXI2X1 U311 ( .A(n189), .B(n130), .S0(quotient[1]), .Y(\u_div/PartRem[1][9] ) );
  MXI2X1 U312 ( .A(n24), .B(\u_div/SumTmp[2][8] ), .S0(quotient[2]), .Y(n188)
         );
  XOR2X1 U313 ( .A(n24), .B(\u_div/CryTmp[2][8] ), .Y(\u_div/SumTmp[2][8] ) );
  MXI2X1 U314 ( .A(n25), .B(\u_div/SumTmp[17][8] ), .S0(n233), .Y(n208) );
  XOR2X1 U315 ( .A(n25), .B(\u_div/CryTmp[17][8] ), .Y(\u_div/SumTmp[17][8] )
         );
  XOR2X1 U316 ( .A(n78), .B(\u_div/CryTmp[16][6] ), .Y(\u_div/SumTmp[16][6] )
         );
  XOR2X1 U317 ( .A(n99), .B(\u_div/CryTmp[16][7] ), .Y(\u_div/SumTmp[16][7] )
         );
  XOR2X1 U318 ( .A(n79), .B(\u_div/CryTmp[15][6] ), .Y(\u_div/SumTmp[15][6] )
         );
  XOR2X1 U319 ( .A(n100), .B(\u_div/CryTmp[7][7] ), .Y(\u_div/SumTmp[7][7] )
         );
  XOR2X1 U320 ( .A(n101), .B(\u_div/CryTmp[6][7] ), .Y(\u_div/SumTmp[6][7] )
         );
  XOR2X1 U321 ( .A(n102), .B(\u_div/CryTmp[5][7] ), .Y(\u_div/SumTmp[5][7] )
         );
  XOR2X1 U322 ( .A(n103), .B(\u_div/CryTmp[4][7] ), .Y(\u_div/SumTmp[4][7] )
         );
  XOR2X1 U323 ( .A(n104), .B(\u_div/CryTmp[3][7] ), .Y(\u_div/SumTmp[3][7] )
         );
  XOR2X1 U324 ( .A(n105), .B(\u_div/CryTmp[17][7] ), .Y(\u_div/SumTmp[17][7] )
         );
  INVX1 U325 ( .A(n189), .Y(\u_div/PartRem[2][8] ) );
  MXI2X1 U326 ( .A(n26), .B(\u_div/SumTmp[18][8] ), .S0(n232), .Y(n207) );
  XOR2X1 U327 ( .A(n26), .B(\u_div/CryTmp[18][8] ), .Y(\u_div/SumTmp[18][8] )
         );
  INVX1 U328 ( .A(n206), .Y(\u_div/PartRem[19][9] ) );
  XNOR2X1 U329 ( .A(\u_div/PartRem[20][9] ), .B(\u_div/CryTmp[19][9] ), .Y(
        n154) );
  AND2X2 U330 ( .A(\u_div/CryTmp[17][5] ), .B(n53), .Y(\u_div/CryTmp[17][6] )
         );
  AND2X2 U331 ( .A(\u_div/CryTmp[17][6] ), .B(n86), .Y(\u_div/CryTmp[17][7] )
         );
  AND2X2 U332 ( .A(\u_div/CryTmp[16][5] ), .B(n54), .Y(\u_div/CryTmp[16][6] )
         );
  AND2X2 U333 ( .A(\u_div/CryTmp[15][5] ), .B(n55), .Y(\u_div/CryTmp[15][6] )
         );
  AND2X2 U334 ( .A(\u_div/CryTmp[14][5] ), .B(n56), .Y(\u_div/CryTmp[14][6] )
         );
  AND2X2 U335 ( .A(\u_div/CryTmp[13][5] ), .B(n57), .Y(\u_div/CryTmp[13][6] )
         );
  AND2X2 U336 ( .A(\u_div/CryTmp[12][5] ), .B(n58), .Y(\u_div/CryTmp[12][6] )
         );
  AND2X2 U337 ( .A(\u_div/CryTmp[11][5] ), .B(n59), .Y(\u_div/CryTmp[11][6] )
         );
  AND2X2 U338 ( .A(\u_div/CryTmp[10][5] ), .B(n60), .Y(\u_div/CryTmp[10][6] )
         );
  AND2X2 U339 ( .A(\u_div/CryTmp[9][5] ), .B(n51), .Y(\u_div/CryTmp[9][6] ) );
  AND2X2 U340 ( .A(\u_div/CryTmp[8][5] ), .B(n52), .Y(\u_div/CryTmp[8][6] ) );
  AND2X2 U341 ( .A(\u_div/CryTmp[7][6] ), .B(n80), .Y(\u_div/CryTmp[7][7] ) );
  AND2X2 U342 ( .A(\u_div/CryTmp[6][6] ), .B(n81), .Y(\u_div/CryTmp[6][7] ) );
  AND2X2 U343 ( .A(\u_div/CryTmp[5][6] ), .B(n82), .Y(\u_div/CryTmp[5][7] ) );
  AND2X2 U344 ( .A(\u_div/CryTmp[4][6] ), .B(n83), .Y(\u_div/CryTmp[4][7] ) );
  AND2X2 U345 ( .A(\u_div/CryTmp[3][6] ), .B(n84), .Y(\u_div/CryTmp[3][7] ) );
  AND2X2 U346 ( .A(\u_div/CryTmp[2][7] ), .B(n106), .Y(\u_div/CryTmp[2][8] )
         );
  AND2X2 U347 ( .A(\u_div/CryTmp[1][7] ), .B(\u_div/PartRem[2][7] ), .Y(
        \u_div/CryTmp[1][8] ) );
  OR2X2 U348 ( .A(\u_div/CryTmp[18][10] ), .B(\u_div/PartRem[19][10] ), .Y(
        n232) );
  MXI2X1 U349 ( .A(n199), .B(n154), .S0(n231), .Y(\u_div/PartRem[19][10] ) );
  XOR2X1 U350 ( .A(n51), .B(\u_div/CryTmp[9][5] ), .Y(\u_div/SumTmp[9][5] ) );
  XOR2X1 U351 ( .A(n52), .B(\u_div/CryTmp[8][5] ), .Y(\u_div/SumTmp[8][5] ) );
  XOR2X1 U352 ( .A(n80), .B(\u_div/CryTmp[7][6] ), .Y(\u_div/SumTmp[7][6] ) );
  XOR2X1 U353 ( .A(n81), .B(\u_div/CryTmp[6][6] ), .Y(\u_div/SumTmp[6][6] ) );
  XOR2X1 U354 ( .A(n82), .B(\u_div/CryTmp[5][6] ), .Y(\u_div/SumTmp[5][6] ) );
  XOR2X1 U355 ( .A(n83), .B(\u_div/CryTmp[4][6] ), .Y(\u_div/SumTmp[4][6] ) );
  XOR2X1 U356 ( .A(n84), .B(\u_div/CryTmp[3][6] ), .Y(\u_div/SumTmp[3][6] ) );
  XOR2X1 U357 ( .A(n53), .B(\u_div/CryTmp[17][5] ), .Y(\u_div/SumTmp[17][5] )
         );
  XOR2X1 U358 ( .A(n54), .B(\u_div/CryTmp[16][5] ), .Y(\u_div/SumTmp[16][5] )
         );
  XOR2X1 U359 ( .A(n55), .B(\u_div/CryTmp[15][5] ), .Y(\u_div/SumTmp[15][5] )
         );
  XOR2X1 U360 ( .A(n56), .B(\u_div/CryTmp[14][5] ), .Y(\u_div/SumTmp[14][5] )
         );
  XOR2X1 U361 ( .A(n57), .B(\u_div/CryTmp[13][5] ), .Y(\u_div/SumTmp[13][5] )
         );
  XOR2X1 U362 ( .A(n58), .B(\u_div/CryTmp[12][5] ), .Y(\u_div/SumTmp[12][5] )
         );
  XOR2X1 U363 ( .A(n59), .B(\u_div/CryTmp[11][5] ), .Y(\u_div/SumTmp[11][5] )
         );
  XOR2X1 U364 ( .A(n60), .B(\u_div/CryTmp[10][5] ), .Y(\u_div/SumTmp[10][5] )
         );
  INVX1 U365 ( .A(n190), .Y(\u_div/PartRem[2][7] ) );
  AND2X2 U366 ( .A(\u_div/CryTmp[19][7] ), .B(n108), .Y(\u_div/CryTmp[19][8] )
         );
  AND2X2 U367 ( .A(\u_div/CryTmp[19][8] ), .B(n27), .Y(\u_div/CryTmp[19][9] )
         );
  AND2X2 U368 ( .A(\u_div/CryTmp[18][6] ), .B(n85), .Y(\u_div/CryTmp[18][7] )
         );
  AND2X2 U369 ( .A(\u_div/CryTmp[18][7] ), .B(n107), .Y(\u_div/CryTmp[18][8] )
         );
  MXI2X1 U370 ( .A(n190), .B(n131), .S0(quotient[1]), .Y(\u_div/PartRem[1][8] ) );
  MXI2X1 U371 ( .A(n106), .B(\u_div/SumTmp[2][7] ), .S0(quotient[2]), .Y(n189)
         );
  XOR2X1 U372 ( .A(n106), .B(\u_div/CryTmp[2][7] ), .Y(\u_div/SumTmp[2][7] )
         );
  XOR2X1 U373 ( .A(n85), .B(\u_div/CryTmp[18][6] ), .Y(\u_div/SumTmp[18][6] )
         );
  XOR2X1 U374 ( .A(n107), .B(\u_div/CryTmp[18][7] ), .Y(\u_div/SumTmp[18][7] )
         );
  XOR2X1 U375 ( .A(n86), .B(\u_div/CryTmp[17][6] ), .Y(\u_div/SumTmp[17][6] )
         );
  XOR2X1 U376 ( .A(n108), .B(\u_div/CryTmp[19][7] ), .Y(\u_div/SumTmp[19][7] )
         );
  MXI2X1 U377 ( .A(n27), .B(\u_div/SumTmp[19][8] ), .S0(n231), .Y(n206) );
  XOR2X1 U378 ( .A(n27), .B(\u_div/CryTmp[19][8] ), .Y(\u_div/SumTmp[19][8] )
         );
  INVX1 U379 ( .A(n199), .Y(\u_div/PartRem[20][9] ) );
  XNOR2X1 U380 ( .A(\u_div/PartRem[21][9] ), .B(\u_div/CryTmp[20][9] ), .Y(
        n155) );
  XNOR2X1 U381 ( .A(\u_div/PartRem[22][9] ), .B(\u_div/CryTmp[21][9] ), .Y(
        n156) );
  AND2X2 U382 ( .A(\u_div/CryTmp[7][5] ), .B(n61), .Y(\u_div/CryTmp[7][6] ) );
  AND2X2 U383 ( .A(\u_div/CryTmp[6][5] ), .B(n62), .Y(\u_div/CryTmp[6][6] ) );
  AND2X2 U384 ( .A(\u_div/CryTmp[5][5] ), .B(n63), .Y(\u_div/CryTmp[5][6] ) );
  AND2X2 U385 ( .A(\u_div/CryTmp[4][5] ), .B(n64), .Y(\u_div/CryTmp[4][6] ) );
  AND2X2 U386 ( .A(\u_div/CryTmp[3][5] ), .B(n65), .Y(\u_div/CryTmp[3][6] ) );
  AND2X2 U387 ( .A(\u_div/CryTmp[2][6] ), .B(n87), .Y(\u_div/CryTmp[2][7] ) );
  OR2X2 U388 ( .A(\u_div/CryTmp[17][4] ), .B(n41), .Y(\u_div/CryTmp[17][5] )
         );
  OR2X2 U389 ( .A(\u_div/CryTmp[16][4] ), .B(n36), .Y(\u_div/CryTmp[16][5] )
         );
  OR2X2 U390 ( .A(\u_div/CryTmp[15][4] ), .B(n42), .Y(\u_div/CryTmp[15][5] )
         );
  OR2X2 U391 ( .A(\u_div/CryTmp[14][4] ), .B(n37), .Y(\u_div/CryTmp[14][5] )
         );
  OR2X2 U392 ( .A(\u_div/CryTmp[13][4] ), .B(n43), .Y(\u_div/CryTmp[13][5] )
         );
  OR2X2 U393 ( .A(\u_div/CryTmp[12][4] ), .B(n38), .Y(\u_div/CryTmp[12][5] )
         );
  OR2X2 U394 ( .A(\u_div/CryTmp[11][4] ), .B(n44), .Y(\u_div/CryTmp[11][5] )
         );
  OR2X2 U395 ( .A(\u_div/CryTmp[10][4] ), .B(n45), .Y(\u_div/CryTmp[10][5] )
         );
  OR2X2 U396 ( .A(\u_div/CryTmp[9][4] ), .B(n39), .Y(\u_div/CryTmp[9][5] ) );
  OR2X2 U397 ( .A(\u_div/CryTmp[8][4] ), .B(n40), .Y(\u_div/CryTmp[8][5] ) );
  AND2X2 U398 ( .A(\u_div/CryTmp[1][6] ), .B(\u_div/PartRem[2][6] ), .Y(
        \u_div/CryTmp[1][7] ) );
  OR2X2 U399 ( .A(\u_div/CryTmp[19][10] ), .B(\u_div/PartRem[20][10] ), .Y(
        n231) );
  MXI2X1 U400 ( .A(n198), .B(n155), .S0(n230), .Y(\u_div/PartRem[20][10] ) );
  MXI2X1 U401 ( .A(n87), .B(\u_div/SumTmp[2][6] ), .S0(quotient[2]), .Y(n190)
         );
  XOR2X1 U402 ( .A(n87), .B(\u_div/CryTmp[2][6] ), .Y(\u_div/SumTmp[2][6] ) );
  XNOR2X1 U403 ( .A(n3), .B(\u_div/CryTmp[18][4] ), .Y(\u_div/SumTmp[18][4] )
         );
  XNOR2X1 U404 ( .A(n36), .B(\u_div/CryTmp[16][4] ), .Y(\u_div/SumTmp[16][4] )
         );
  XNOR2X1 U405 ( .A(n37), .B(\u_div/CryTmp[14][4] ), .Y(\u_div/SumTmp[14][4] )
         );
  XNOR2X1 U406 ( .A(n38), .B(\u_div/CryTmp[12][4] ), .Y(\u_div/SumTmp[12][4] )
         );
  XNOR2X1 U407 ( .A(n39), .B(\u_div/CryTmp[9][4] ), .Y(\u_div/SumTmp[9][4] )
         );
  XNOR2X1 U408 ( .A(n40), .B(\u_div/CryTmp[8][4] ), .Y(\u_div/SumTmp[8][4] )
         );
  XOR2X1 U409 ( .A(n61), .B(\u_div/CryTmp[7][5] ), .Y(\u_div/SumTmp[7][5] ) );
  XOR2X1 U410 ( .A(n62), .B(\u_div/CryTmp[6][5] ), .Y(\u_div/SumTmp[6][5] ) );
  XOR2X1 U411 ( .A(n63), .B(\u_div/CryTmp[5][5] ), .Y(\u_div/SumTmp[5][5] ) );
  XOR2X1 U412 ( .A(n64), .B(\u_div/CryTmp[4][5] ), .Y(\u_div/SumTmp[4][5] ) );
  XOR2X1 U413 ( .A(n65), .B(\u_div/CryTmp[3][5] ), .Y(\u_div/SumTmp[3][5] ) );
  XOR2X1 U414 ( .A(n66), .B(\u_div/CryTmp[19][5] ), .Y(\u_div/SumTmp[19][5] )
         );
  XOR2X1 U415 ( .A(n67), .B(\u_div/CryTmp[18][5] ), .Y(\u_div/SumTmp[18][5] )
         );
  XNOR2X1 U416 ( .A(n41), .B(\u_div/CryTmp[17][4] ), .Y(\u_div/SumTmp[17][4] )
         );
  XNOR2X1 U417 ( .A(n42), .B(\u_div/CryTmp[15][4] ), .Y(\u_div/SumTmp[15][4] )
         );
  XNOR2X1 U418 ( .A(n43), .B(\u_div/CryTmp[13][4] ), .Y(\u_div/SumTmp[13][4] )
         );
  XNOR2X1 U419 ( .A(n44), .B(\u_div/CryTmp[11][4] ), .Y(\u_div/SumTmp[11][4] )
         );
  XNOR2X1 U420 ( .A(n45), .B(\u_div/CryTmp[10][4] ), .Y(\u_div/SumTmp[10][4] )
         );
  INVX1 U421 ( .A(n191), .Y(\u_div/PartRem[2][6] ) );
  AND2X2 U422 ( .A(\u_div/CryTmp[21][6] ), .B(n90), .Y(\u_div/CryTmp[21][7] )
         );
  AND2X2 U423 ( .A(\u_div/CryTmp[21][7] ), .B(n110), .Y(\u_div/CryTmp[21][8] )
         );
  AND2X2 U424 ( .A(\u_div/CryTmp[21][8] ), .B(n111), .Y(\u_div/CryTmp[21][9] )
         );
  AND2X2 U425 ( .A(\u_div/CryTmp[20][6] ), .B(n88), .Y(\u_div/CryTmp[20][7] )
         );
  AND2X2 U426 ( .A(\u_div/CryTmp[20][7] ), .B(n109), .Y(\u_div/CryTmp[20][8] )
         );
  AND2X2 U427 ( .A(\u_div/CryTmp[20][8] ), .B(n28), .Y(\u_div/CryTmp[20][9] )
         );
  AND2X2 U428 ( .A(\u_div/CryTmp[19][5] ), .B(n66), .Y(\u_div/CryTmp[19][6] )
         );
  AND2X2 U429 ( .A(\u_div/CryTmp[19][6] ), .B(n89), .Y(\u_div/CryTmp[19][7] )
         );
  AND2X2 U430 ( .A(\u_div/CryTmp[18][5] ), .B(n67), .Y(\u_div/CryTmp[18][6] )
         );
  OR2X2 U431 ( .A(\u_div/CryTmp[18][4] ), .B(n3), .Y(\u_div/CryTmp[18][5] ) );
  MXI2X1 U432 ( .A(n191), .B(n132), .S0(quotient[1]), .Y(\u_div/PartRem[1][7] ) );
  XOR2X1 U433 ( .A(n88), .B(\u_div/CryTmp[20][6] ), .Y(\u_div/SumTmp[20][6] )
         );
  XOR2X1 U434 ( .A(n89), .B(\u_div/CryTmp[19][6] ), .Y(\u_div/SumTmp[19][6] )
         );
  XOR2X1 U435 ( .A(n109), .B(\u_div/CryTmp[20][7] ), .Y(\u_div/SumTmp[20][7] )
         );
  MXI2X1 U436 ( .A(n28), .B(\u_div/SumTmp[20][8] ), .S0(n230), .Y(n199) );
  XOR2X1 U437 ( .A(n28), .B(\u_div/CryTmp[20][8] ), .Y(\u_div/SumTmp[20][8] )
         );
  INVX1 U438 ( .A(n198), .Y(\u_div/PartRem[21][9] ) );
  INVX1 U439 ( .A(n196), .Y(\u_div/PartRem[22][9] ) );
  INVX1 U440 ( .A(n195), .Y(\u_div/CryTmp[8][4] ) );
  MXI2X1 U441 ( .A(n31), .B(n31), .S0(quotient[9]), .Y(n195) );
  INVX1 U442 ( .A(n220), .Y(\u_div/CryTmp[17][4] ) );
  MXI2X1 U443 ( .A(n118), .B(n118), .S0(n232), .Y(n220) );
  INVX1 U444 ( .A(n228), .Y(\u_div/CryTmp[16][4] ) );
  MXI2X1 U445 ( .A(n119), .B(n119), .S0(n233), .Y(n228) );
  INVX1 U446 ( .A(n221), .Y(\u_div/CryTmp[15][4] ) );
  MXI2X1 U447 ( .A(n120), .B(n120), .S0(n234), .Y(n221) );
  INVX1 U448 ( .A(n222), .Y(\u_div/CryTmp[14][4] ) );
  MXI2X1 U449 ( .A(n121), .B(n121), .S0(n235), .Y(n222) );
  INVX1 U450 ( .A(n223), .Y(\u_div/CryTmp[13][4] ) );
  MXI2X1 U451 ( .A(n122), .B(n122), .S0(n236), .Y(n223) );
  INVX1 U452 ( .A(n224), .Y(\u_div/CryTmp[12][4] ) );
  MXI2X1 U453 ( .A(n123), .B(n123), .S0(n237), .Y(n224) );
  INVX1 U454 ( .A(n225), .Y(\u_div/CryTmp[11][4] ) );
  MXI2X1 U455 ( .A(n124), .B(n124), .S0(n238), .Y(n225) );
  INVX1 U456 ( .A(n226), .Y(\u_div/CryTmp[10][4] ) );
  MXI2X1 U457 ( .A(n125), .B(n125), .S0(n239), .Y(n226) );
  INVX1 U458 ( .A(n227), .Y(\u_div/CryTmp[9][4] ) );
  MXI2X1 U459 ( .A(n126), .B(n126), .S0(n240), .Y(n227) );
  INVX1 U460 ( .A(n193), .Y(\u_div/PartRem[2][4] ) );
  AND2X2 U461 ( .A(\u_div/CryTmp[2][5] ), .B(n68), .Y(\u_div/CryTmp[2][6] ) );
  OR2X2 U462 ( .A(\u_div/CryTmp[7][4] ), .B(n4), .Y(\u_div/CryTmp[7][5] ) );
  OR2X2 U463 ( .A(\u_div/CryTmp[6][4] ), .B(n46), .Y(\u_div/CryTmp[6][5] ) );
  OR2X2 U464 ( .A(\u_div/CryTmp[5][4] ), .B(n47), .Y(\u_div/CryTmp[5][5] ) );
  OR2X2 U465 ( .A(\u_div/CryTmp[4][4] ), .B(n48), .Y(\u_div/CryTmp[4][5] ) );
  OR2X2 U466 ( .A(\u_div/CryTmp[3][4] ), .B(n49), .Y(\u_div/CryTmp[3][5] ) );
  AND2X2 U467 ( .A(\u_div/CryTmp[1][5] ), .B(\u_div/PartRem[2][5] ), .Y(
        \u_div/CryTmp[1][6] ) );
  AND2X2 U468 ( .A(\u_div/CryTmp[22][9] ), .B(a[31]), .Y(
        \u_div/CryTmp[22][10] ) );
  MXI2X1 U469 ( .A(n68), .B(\u_div/SumTmp[2][5] ), .S0(quotient[2]), .Y(n191)
         );
  XOR2X1 U470 ( .A(n68), .B(\u_div/CryTmp[2][5] ), .Y(\u_div/SumTmp[2][5] ) );
  INVX1 U471 ( .A(n218), .Y(\u_div/CryTmp[18][4] ) );
  MXI2X1 U472 ( .A(n129), .B(n129), .S0(n231), .Y(n218) );
  XNOR2X1 U473 ( .A(n4), .B(\u_div/CryTmp[7][4] ), .Y(\u_div/SumTmp[7][4] ) );
  XNOR2X1 U474 ( .A(n46), .B(\u_div/CryTmp[6][4] ), .Y(\u_div/SumTmp[6][4] )
         );
  XNOR2X1 U475 ( .A(n47), .B(\u_div/CryTmp[5][4] ), .Y(\u_div/SumTmp[5][4] )
         );
  XNOR2X1 U476 ( .A(n48), .B(\u_div/CryTmp[4][4] ), .Y(\u_div/SumTmp[4][4] )
         );
  XNOR2X1 U477 ( .A(n49), .B(\u_div/CryTmp[3][4] ), .Y(\u_div/SumTmp[3][4] )
         );
  XNOR2X1 U478 ( .A(n50), .B(\u_div/CryTmp[20][4] ), .Y(\u_div/SumTmp[20][4] )
         );
  XOR2X1 U479 ( .A(n69), .B(\u_div/CryTmp[20][5] ), .Y(\u_div/SumTmp[20][5] )
         );
  XNOR2X1 U480 ( .A(n5), .B(\u_div/CryTmp[19][4] ), .Y(\u_div/SumTmp[19][4] )
         );
  INVX1 U481 ( .A(n192), .Y(\u_div/PartRem[2][5] ) );
  AND2X2 U482 ( .A(\u_div/CryTmp[21][5] ), .B(n70), .Y(\u_div/CryTmp[21][6] )
         );
  AND2X2 U483 ( .A(\u_div/CryTmp[20][5] ), .B(n69), .Y(\u_div/CryTmp[20][6] )
         );
  OR2X2 U484 ( .A(\u_div/CryTmp[20][4] ), .B(n50), .Y(\u_div/CryTmp[20][5] )
         );
  OR2X2 U485 ( .A(\u_div/CryTmp[19][4] ), .B(n5), .Y(\u_div/CryTmp[19][5] ) );
  MXI2X1 U486 ( .A(n192), .B(n114), .S0(quotient[1]), .Y(\u_div/PartRem[1][6] ) );
  MX2X1 U487 ( .A(n196), .B(n156), .S0(n229), .Y(n157) );
  XOR2X1 U488 ( .A(n90), .B(\u_div/CryTmp[21][6] ), .Y(\u_div/SumTmp[21][6] )
         );
  XOR2X1 U489 ( .A(\u_div/PartRem[28][1] ), .B(\u_div/CryTmp[22][6] ), .Y(
        \u_div/SumTmp[22][6] ) );
  XOR2X1 U490 ( .A(n70), .B(\u_div/CryTmp[21][5] ), .Y(\u_div/SumTmp[21][5] )
         );
  XOR2X1 U491 ( .A(n110), .B(\u_div/CryTmp[21][7] ), .Y(\u_div/SumTmp[21][7] )
         );
  XOR2X1 U492 ( .A(a[27]), .B(\u_div/CryTmp[22][5] ), .Y(\u_div/SumTmp[22][5] ) );
  XOR2X1 U493 ( .A(\u_div/PartRem[29][1] ), .B(\u_div/CryTmp[22][7] ), .Y(
        \u_div/SumTmp[22][7] ) );
  AND2X2 U494 ( .A(\u_div/CryTmp[22][5] ), .B(a[27]), .Y(\u_div/CryTmp[22][6] ) );
  AND2X2 U495 ( .A(\u_div/CryTmp[22][6] ), .B(\u_div/PartRem[28][1] ), .Y(
        \u_div/CryTmp[22][7] ) );
  AND2X2 U496 ( .A(\u_div/CryTmp[22][7] ), .B(\u_div/PartRem[29][1] ), .Y(
        \u_div/CryTmp[22][8] ) );
  AND2X2 U497 ( .A(\u_div/CryTmp[22][8] ), .B(\u_div/PartRem[30][1] ), .Y(
        \u_div/CryTmp[22][9] ) );
  MXI2X1 U498 ( .A(n111), .B(\u_div/SumTmp[21][8] ), .S0(n229), .Y(n198) );
  XOR2X1 U499 ( .A(n111), .B(\u_div/CryTmp[21][8] ), .Y(\u_div/SumTmp[21][8] )
         );
  MXI2X1 U500 ( .A(\u_div/PartRem[30][1] ), .B(\u_div/SumTmp[22][8] ), .S0(
        \u_div/CryTmp[22][10] ), .Y(n196) );
  XOR2X1 U501 ( .A(\u_div/PartRem[30][1] ), .B(\u_div/CryTmp[22][8] ), .Y(
        \u_div/SumTmp[22][8] ) );
  XNOR2X1 U502 ( .A(a[31]), .B(\u_div/CryTmp[22][9] ), .Y(n158) );
  MXI2X1 U503 ( .A(\u_div/CryTmp[2][4] ), .B(n204), .S0(quotient[2]), .Y(n193)
         );
  INVX1 U504 ( .A(n205), .Y(\u_div/CryTmp[7][4] ) );
  MXI2X1 U505 ( .A(n127), .B(n127), .S0(quotient[8]), .Y(n205) );
  INVX1 U506 ( .A(n200), .Y(\u_div/CryTmp[6][4] ) );
  MXI2X1 U507 ( .A(n115), .B(n115), .S0(quotient[7]), .Y(n200) );
  INVX1 U508 ( .A(n201), .Y(\u_div/CryTmp[5][4] ) );
  MXI2X1 U509 ( .A(n116), .B(n116), .S0(quotient[6]), .Y(n201) );
  INVX1 U510 ( .A(n202), .Y(\u_div/CryTmp[4][4] ) );
  MXI2X1 U511 ( .A(n117), .B(n117), .S0(quotient[5]), .Y(n202) );
  INVX1 U512 ( .A(n203), .Y(\u_div/CryTmp[3][4] ) );
  MXI2X1 U513 ( .A(n30), .B(n30), .S0(quotient[4]), .Y(n203) );
  OR2X2 U514 ( .A(\u_div/CryTmp[2][4] ), .B(n2), .Y(\u_div/CryTmp[2][5] ) );
  OR2X2 U515 ( .A(\u_div/CryTmp[1][4] ), .B(\u_div/PartRem[2][4] ), .Y(
        \u_div/CryTmp[1][5] ) );
  MX2X1 U516 ( .A(n197), .B(n158), .S0(\u_div/CryTmp[22][10] ), .Y(n159) );
  MXI2X1 U517 ( .A(n2), .B(\u_div/SumTmp[2][4] ), .S0(quotient[2]), .Y(n192)
         );
  XNOR2X1 U518 ( .A(n2), .B(\u_div/CryTmp[2][4] ), .Y(\u_div/SumTmp[2][4] ) );
  INVX1 U519 ( .A(n214), .Y(\u_div/CryTmp[20][4] ) );
  MXI2X1 U520 ( .A(n29), .B(n29), .S0(n229), .Y(n214) );
  INVX1 U521 ( .A(n216), .Y(\u_div/CryTmp[19][4] ) );
  MXI2X1 U522 ( .A(n32), .B(n32), .S0(n230), .Y(n216) );
  XNOR2X1 U523 ( .A(n1), .B(\u_div/CryTmp[21][4] ), .Y(\u_div/SumTmp[21][4] )
         );
  XNOR2X1 U524 ( .A(a[26]), .B(a[25]), .Y(\u_div/SumTmp[22][4] ) );
  OR2X2 U525 ( .A(\u_div/CryTmp[21][4] ), .B(n1), .Y(\u_div/CryTmp[21][5] ) );
  MXI2X1 U526 ( .A(n193), .B(n113), .S0(quotient[1]), .Y(\u_div/PartRem[1][5] ) );
  NAND2BX1 U527 ( .AN(\u_div/CryTmp[0][4] ), .B(n6), .Y(\u_div/CryTmp[0][5] )
         );
  OR2X2 U528 ( .A(a[25]), .B(a[26]), .Y(\u_div/CryTmp[22][5] ) );
  MX2X1 U529 ( .A(\u_div/SumTmp[16][0] ), .B(\u_div/SumTmp[16][0] ), .S0(n234), 
        .Y(n160) );
  MX2X1 U530 ( .A(\u_div/SumTmp[14][0] ), .B(\u_div/SumTmp[14][0] ), .S0(n236), 
        .Y(n161) );
  MX2X1 U531 ( .A(\u_div/SumTmp[12][0] ), .B(\u_div/SumTmp[12][0] ), .S0(n238), 
        .Y(n162) );
  MX2X1 U532 ( .A(\u_div/SumTmp[15][0] ), .B(\u_div/SumTmp[15][0] ), .S0(n235), 
        .Y(n163) );
  MX2X1 U533 ( .A(\u_div/SumTmp[13][0] ), .B(\u_div/SumTmp[13][0] ), .S0(n237), 
        .Y(n164) );
  MX2X1 U534 ( .A(\u_div/SumTmp[11][0] ), .B(\u_div/SumTmp[11][0] ), .S0(n239), 
        .Y(n165) );
  MX2X1 U535 ( .A(\u_div/SumTmp[18][0] ), .B(\u_div/SumTmp[18][0] ), .S0(n232), 
        .Y(n166) );
  MX2X1 U536 ( .A(\u_div/SumTmp[21][0] ), .B(\u_div/SumTmp[21][0] ), .S0(n229), 
        .Y(n167) );
  MX2X1 U537 ( .A(\u_div/SumTmp[20][0] ), .B(\u_div/SumTmp[20][0] ), .S0(n230), 
        .Y(n168) );
  MX2X1 U538 ( .A(\u_div/SumTmp[19][0] ), .B(\u_div/SumTmp[19][0] ), .S0(n231), 
        .Y(n169) );
  MX2X1 U539 ( .A(\u_div/SumTmp[17][0] ), .B(\u_div/SumTmp[17][0] ), .S0(n233), 
        .Y(n170) );
  INVX1 U540 ( .A(n204), .Y(\u_div/CryTmp[2][4] ) );
  MXI2X1 U541 ( .A(n128), .B(n128), .S0(quotient[3]), .Y(n204) );
  INVX1 U542 ( .A(n194), .Y(\u_div/CryTmp[1][4] ) );
  INVX1 U543 ( .A(n212), .Y(\u_div/CryTmp[21][4] ) );
  MXI2X1 U544 ( .A(a[24]), .B(a[24]), .S0(\u_div/CryTmp[22][10] ), .Y(n212) );
  MX2X1 U545 ( .A(n171), .B(n171), .S0(quotient[1]), .Y(\u_div/CryTmp[0][4] )
         );
  MX2X1 U546 ( .A(n178), .B(n178), .S0(quotient[2]), .Y(n171) );
  MX2X1 U547 ( .A(\u_div/SumTmp[10][0] ), .B(\u_div/SumTmp[10][0] ), .S0(n240), 
        .Y(n172) );
  MX2X1 U548 ( .A(\u_div/SumTmp[9][0] ), .B(\u_div/SumTmp[9][0] ), .S0(
        quotient[9]), .Y(n173) );
  MX2X1 U549 ( .A(\u_div/SumTmp[8][0] ), .B(\u_div/SumTmp[8][0] ), .S0(
        quotient[8]), .Y(n174) );
  MX2X1 U550 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[7][0] ), .S0(
        quotient[7]), .Y(n175) );
  MX2X1 U551 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[6][0] ), .S0(
        quotient[6]), .Y(n176) );
  MX2X1 U552 ( .A(\u_div/SumTmp[22][0] ), .B(\u_div/SumTmp[22][0] ), .S0(
        \u_div/CryTmp[22][10] ), .Y(n177) );
  MXI2X1 U553 ( .A(n33), .B(n33), .S0(quotient[2]), .Y(n194) );
  INVX1 U554 ( .A(a[25]), .Y(n210) );
  MX2X1 U555 ( .A(\u_div/SumTmp[3][0] ), .B(\u_div/SumTmp[3][0] ), .S0(
        quotient[3]), .Y(n178) );
  MX2X1 U556 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[5][0] ), .S0(
        quotient[5]), .Y(n179) );
  INVX1 U557 ( .A(a[31]), .Y(n197) );
  NAND2BX4 U558 ( .AN(\u_div/CryTmp[9][10] ), .B(n134), .Y(quotient[9]) );
endmodule


module Equation_Implementation_DW_div_uns_24 ( a, b, quotient, remainder, 
        divide_by_0 );
  input [31:0] a;
  input [16:0] b;
  output [31:0] quotient;
  output [16:0] remainder;
  output divide_by_0;
  wire   n272, n273, n274, n275, n276, \u_div/SumTmp[2][6] ,
         \u_div/SumTmp[2][7] , \u_div/SumTmp[2][8] , \u_div/SumTmp[2][9] ,
         \u_div/SumTmp[2][10] , \u_div/SumTmp[2][11] , \u_div/SumTmp[2][12] ,
         \u_div/SumTmp[2][13] , \u_div/SumTmp[2][14] , \u_div/SumTmp[2][15] ,
         \u_div/SumTmp[3][6] , \u_div/SumTmp[3][7] , \u_div/SumTmp[3][8] ,
         \u_div/SumTmp[3][9] , \u_div/SumTmp[3][10] , \u_div/SumTmp[3][11] ,
         \u_div/SumTmp[3][12] , \u_div/SumTmp[3][13] , \u_div/SumTmp[3][14] ,
         \u_div/SumTmp[3][15] , \u_div/SumTmp[4][6] , \u_div/SumTmp[4][7] ,
         \u_div/SumTmp[4][8] , \u_div/SumTmp[4][9] , \u_div/SumTmp[4][10] ,
         \u_div/SumTmp[4][11] , \u_div/SumTmp[4][12] , \u_div/SumTmp[4][13] ,
         \u_div/SumTmp[4][14] , \u_div/SumTmp[4][15] , \u_div/SumTmp[5][0] ,
         \u_div/SumTmp[5][6] , \u_div/SumTmp[5][7] , \u_div/SumTmp[5][8] ,
         \u_div/SumTmp[5][9] , \u_div/SumTmp[5][10] , \u_div/SumTmp[5][11] ,
         \u_div/SumTmp[5][12] , \u_div/SumTmp[5][13] , \u_div/SumTmp[5][14] ,
         \u_div/SumTmp[5][15] , \u_div/SumTmp[6][0] , \u_div/SumTmp[6][6] ,
         \u_div/SumTmp[6][7] , \u_div/SumTmp[6][8] , \u_div/SumTmp[6][9] ,
         \u_div/SumTmp[6][10] , \u_div/SumTmp[6][11] , \u_div/SumTmp[6][12] ,
         \u_div/SumTmp[6][13] , \u_div/SumTmp[6][14] , \u_div/SumTmp[6][15] ,
         \u_div/SumTmp[7][0] , \u_div/SumTmp[7][6] , \u_div/SumTmp[7][7] ,
         \u_div/SumTmp[7][8] , \u_div/SumTmp[7][9] , \u_div/SumTmp[7][10] ,
         \u_div/SumTmp[7][11] , \u_div/SumTmp[7][12] , \u_div/SumTmp[7][13] ,
         \u_div/SumTmp[7][14] , \u_div/SumTmp[7][15] , \u_div/SumTmp[8][0] ,
         \u_div/SumTmp[8][6] , \u_div/SumTmp[8][7] , \u_div/SumTmp[8][8] ,
         \u_div/SumTmp[8][9] , \u_div/SumTmp[8][10] , \u_div/SumTmp[8][11] ,
         \u_div/SumTmp[8][12] , \u_div/SumTmp[8][13] , \u_div/SumTmp[8][14] ,
         \u_div/SumTmp[8][15] , \u_div/SumTmp[9][0] , \u_div/SumTmp[9][6] ,
         \u_div/SumTmp[9][7] , \u_div/SumTmp[9][8] , \u_div/SumTmp[9][9] ,
         \u_div/SumTmp[9][10] , \u_div/SumTmp[9][11] , \u_div/SumTmp[9][12] ,
         \u_div/SumTmp[9][13] , \u_div/SumTmp[9][14] , \u_div/SumTmp[9][15] ,
         \u_div/SumTmp[10][0] , \u_div/SumTmp[10][6] , \u_div/SumTmp[10][7] ,
         \u_div/SumTmp[10][8] , \u_div/SumTmp[10][9] , \u_div/SumTmp[10][10] ,
         \u_div/SumTmp[10][11] , \u_div/SumTmp[10][12] ,
         \u_div/SumTmp[10][13] , \u_div/SumTmp[10][14] ,
         \u_div/SumTmp[10][15] , \u_div/SumTmp[11][0] , \u_div/SumTmp[11][6] ,
         \u_div/SumTmp[11][7] , \u_div/SumTmp[11][8] , \u_div/SumTmp[11][9] ,
         \u_div/SumTmp[11][10] , \u_div/SumTmp[11][11] ,
         \u_div/SumTmp[11][12] , \u_div/SumTmp[11][13] ,
         \u_div/SumTmp[11][14] , \u_div/SumTmp[11][15] , \u_div/SumTmp[12][0] ,
         \u_div/SumTmp[12][6] , \u_div/SumTmp[12][7] , \u_div/SumTmp[12][8] ,
         \u_div/SumTmp[12][9] , \u_div/SumTmp[12][10] , \u_div/SumTmp[12][11] ,
         \u_div/SumTmp[12][12] , \u_div/SumTmp[12][13] ,
         \u_div/SumTmp[12][14] , \u_div/SumTmp[12][15] , \u_div/SumTmp[13][0] ,
         \u_div/SumTmp[13][6] , \u_div/SumTmp[13][7] , \u_div/SumTmp[13][8] ,
         \u_div/SumTmp[13][9] , \u_div/SumTmp[13][10] , \u_div/SumTmp[13][11] ,
         \u_div/SumTmp[13][12] , \u_div/SumTmp[13][13] ,
         \u_div/SumTmp[13][14] , \u_div/SumTmp[13][15] , \u_div/SumTmp[14][0] ,
         \u_div/SumTmp[14][6] , \u_div/SumTmp[14][7] , \u_div/SumTmp[14][8] ,
         \u_div/SumTmp[14][9] , \u_div/SumTmp[14][10] , \u_div/SumTmp[14][11] ,
         \u_div/SumTmp[14][12] , \u_div/SumTmp[14][13] ,
         \u_div/SumTmp[14][14] , \u_div/SumTmp[14][15] , \u_div/SumTmp[15][0] ,
         \u_div/SumTmp[15][6] , \u_div/SumTmp[15][7] , \u_div/SumTmp[15][8] ,
         \u_div/SumTmp[15][9] , \u_div/SumTmp[15][10] , \u_div/SumTmp[15][11] ,
         \u_div/SumTmp[15][12] , \u_div/SumTmp[15][13] ,
         \u_div/SumTmp[15][14] , \u_div/SumTmp[15][15] , \u_div/CryTmp[0][6] ,
         \u_div/CryTmp[0][7] , \u_div/CryTmp[0][9] , \u_div/CryTmp[0][12] ,
         \u_div/CryTmp[0][13] , \u_div/CryTmp[0][14] , \u_div/CryTmp[0][15] ,
         \u_div/CryTmp[1][6] , \u_div/CryTmp[1][7] , \u_div/CryTmp[1][8] ,
         \u_div/CryTmp[1][9] , \u_div/CryTmp[1][10] , \u_div/CryTmp[1][11] ,
         \u_div/CryTmp[1][12] , \u_div/CryTmp[1][13] , \u_div/CryTmp[1][14] ,
         \u_div/CryTmp[1][15] , \u_div/CryTmp[1][16] , \u_div/CryTmp[1][17] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[2][7] , \u_div/CryTmp[2][8] ,
         \u_div/CryTmp[2][9] , \u_div/CryTmp[2][10] , \u_div/CryTmp[2][11] ,
         \u_div/CryTmp[2][12] , \u_div/CryTmp[2][13] , \u_div/CryTmp[2][14] ,
         \u_div/CryTmp[2][15] , \u_div/CryTmp[2][16] , \u_div/CryTmp[2][17] ,
         \u_div/CryTmp[3][6] , \u_div/CryTmp[3][7] , \u_div/CryTmp[3][8] ,
         \u_div/CryTmp[3][9] , \u_div/CryTmp[3][10] , \u_div/CryTmp[3][11] ,
         \u_div/CryTmp[3][12] , \u_div/CryTmp[3][13] , \u_div/CryTmp[3][14] ,
         \u_div/CryTmp[3][15] , \u_div/CryTmp[3][16] , \u_div/CryTmp[3][17] ,
         \u_div/CryTmp[4][6] , \u_div/CryTmp[4][7] , \u_div/CryTmp[4][8] ,
         \u_div/CryTmp[4][9] , \u_div/CryTmp[4][10] , \u_div/CryTmp[4][11] ,
         \u_div/CryTmp[4][12] , \u_div/CryTmp[4][13] , \u_div/CryTmp[4][14] ,
         \u_div/CryTmp[4][15] , \u_div/CryTmp[4][16] , \u_div/CryTmp[4][17] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[5][7] , \u_div/CryTmp[5][8] ,
         \u_div/CryTmp[5][9] , \u_div/CryTmp[5][10] , \u_div/CryTmp[5][11] ,
         \u_div/CryTmp[5][12] , \u_div/CryTmp[5][13] , \u_div/CryTmp[5][14] ,
         \u_div/CryTmp[5][15] , \u_div/CryTmp[5][16] , \u_div/CryTmp[5][17] ,
         \u_div/CryTmp[6][6] , \u_div/CryTmp[6][7] , \u_div/CryTmp[6][8] ,
         \u_div/CryTmp[6][9] , \u_div/CryTmp[6][10] , \u_div/CryTmp[6][11] ,
         \u_div/CryTmp[6][12] , \u_div/CryTmp[6][13] , \u_div/CryTmp[6][14] ,
         \u_div/CryTmp[6][15] , \u_div/CryTmp[6][16] , \u_div/CryTmp[6][17] ,
         \u_div/CryTmp[7][6] , \u_div/CryTmp[7][7] , \u_div/CryTmp[7][8] ,
         \u_div/CryTmp[7][9] , \u_div/CryTmp[7][10] , \u_div/CryTmp[7][11] ,
         \u_div/CryTmp[7][12] , \u_div/CryTmp[7][13] , \u_div/CryTmp[7][14] ,
         \u_div/CryTmp[7][15] , \u_div/CryTmp[7][16] , \u_div/CryTmp[7][17] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[8][7] , \u_div/CryTmp[8][8] ,
         \u_div/CryTmp[8][9] , \u_div/CryTmp[8][10] , \u_div/CryTmp[8][11] ,
         \u_div/CryTmp[8][12] , \u_div/CryTmp[8][13] , \u_div/CryTmp[8][14] ,
         \u_div/CryTmp[8][15] , \u_div/CryTmp[8][16] , \u_div/CryTmp[8][17] ,
         \u_div/CryTmp[9][6] , \u_div/CryTmp[9][7] , \u_div/CryTmp[9][8] ,
         \u_div/CryTmp[9][9] , \u_div/CryTmp[9][10] , \u_div/CryTmp[9][11] ,
         \u_div/CryTmp[9][12] , \u_div/CryTmp[9][13] , \u_div/CryTmp[9][14] ,
         \u_div/CryTmp[9][15] , \u_div/CryTmp[9][16] , \u_div/CryTmp[9][17] ,
         \u_div/CryTmp[10][6] , \u_div/CryTmp[10][7] , \u_div/CryTmp[10][8] ,
         \u_div/CryTmp[10][9] , \u_div/CryTmp[10][10] , \u_div/CryTmp[10][11] ,
         \u_div/CryTmp[10][12] , \u_div/CryTmp[10][13] ,
         \u_div/CryTmp[10][14] , \u_div/CryTmp[10][15] ,
         \u_div/CryTmp[10][16] , \u_div/CryTmp[10][17] , \u_div/CryTmp[11][6] ,
         \u_div/CryTmp[11][7] , \u_div/CryTmp[11][8] , \u_div/CryTmp[11][9] ,
         \u_div/CryTmp[11][10] , \u_div/CryTmp[11][11] ,
         \u_div/CryTmp[11][12] , \u_div/CryTmp[11][13] ,
         \u_div/CryTmp[11][14] , \u_div/CryTmp[11][15] ,
         \u_div/CryTmp[11][16] , \u_div/CryTmp[11][17] , \u_div/CryTmp[12][6] ,
         \u_div/CryTmp[12][7] , \u_div/CryTmp[12][8] , \u_div/CryTmp[12][9] ,
         \u_div/CryTmp[12][10] , \u_div/CryTmp[12][11] ,
         \u_div/CryTmp[12][12] , \u_div/CryTmp[12][13] ,
         \u_div/CryTmp[12][14] , \u_div/CryTmp[12][15] ,
         \u_div/CryTmp[12][16] , \u_div/CryTmp[12][17] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[13][7] , \u_div/CryTmp[13][8] , \u_div/CryTmp[13][9] ,
         \u_div/CryTmp[13][10] , \u_div/CryTmp[13][11] ,
         \u_div/CryTmp[13][12] , \u_div/CryTmp[13][13] ,
         \u_div/CryTmp[13][14] , \u_div/CryTmp[13][15] ,
         \u_div/CryTmp[13][16] , \u_div/CryTmp[13][17] , \u_div/CryTmp[14][6] ,
         \u_div/CryTmp[14][7] , \u_div/CryTmp[14][8] , \u_div/CryTmp[14][9] ,
         \u_div/CryTmp[14][10] , \u_div/CryTmp[14][11] ,
         \u_div/CryTmp[14][12] , \u_div/CryTmp[14][13] ,
         \u_div/CryTmp[14][14] , \u_div/CryTmp[14][15] ,
         \u_div/CryTmp[14][16] , \u_div/CryTmp[14][17] , \u_div/CryTmp[15][7] ,
         \u_div/CryTmp[15][8] , \u_div/CryTmp[15][9] , \u_div/CryTmp[15][10] ,
         \u_div/CryTmp[15][11] , \u_div/CryTmp[15][12] ,
         \u_div/CryTmp[15][13] , \u_div/CryTmp[15][14] ,
         \u_div/CryTmp[15][15] , \u_div/CryTmp[15][16] ,
         \u_div/CryTmp[15][17] , \u_div/PartRem[1][7] , \u_div/PartRem[1][9] ,
         \u_div/PartRem[1][10] , \u_div/PartRem[1][15] ,
         \u_div/PartRem[1][16] , \u_div/PartRem[2][6] , \u_div/PartRem[2][7] ,
         \u_div/PartRem[2][8] , \u_div/PartRem[2][9] , \u_div/PartRem[2][10] ,
         \u_div/PartRem[2][11] , \u_div/PartRem[2][12] ,
         \u_div/PartRem[2][13] , \u_div/PartRem[2][14] ,
         \u_div/PartRem[2][15] , \u_div/PartRem[2][16] ,
         \u_div/PartRem[2][17] , \u_div/PartRem[3][16] ,
         \u_div/PartRem[3][17] , \u_div/PartRem[4][16] ,
         \u_div/PartRem[4][17] , \u_div/PartRem[5][16] ,
         \u_div/PartRem[5][17] , \u_div/PartRem[6][16] ,
         \u_div/PartRem[6][17] , \u_div/PartRem[7][16] ,
         \u_div/PartRem[7][17] , \u_div/PartRem[8][16] ,
         \u_div/PartRem[8][17] , \u_div/PartRem[9][16] ,
         \u_div/PartRem[9][17] , \u_div/PartRem[10][16] ,
         \u_div/PartRem[10][17] , \u_div/PartRem[11][16] ,
         \u_div/PartRem[12][16] , \u_div/PartRem[13][16] ,
         \u_div/PartRem[14][16] , \u_div/PartRem[15][16] ,
         \u_div/PartRem[18][1] , \u_div/PartRem[19][1] ,
         \u_div/PartRem[20][1] , \u_div/PartRem[21][1] ,
         \u_div/PartRem[22][1] , \u_div/PartRem[23][1] ,
         \u_div/PartRem[24][1] , \u_div/PartRem[25][1] ,
         \u_div/PartRem[31][1] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271;
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[12][0]  = a[12];
  assign \u_div/SumTmp[13][0]  = a[13];
  assign \u_div/SumTmp[14][0]  = a[14];
  assign \u_div/SumTmp[15][0]  = a[15];
  assign \u_div/PartRem[18][1]  = a[18];
  assign \u_div/PartRem[19][1]  = a[19];
  assign \u_div/PartRem[20][1]  = a[20];
  assign \u_div/PartRem[21][1]  = a[21];
  assign \u_div/PartRem[22][1]  = a[22];
  assign \u_div/PartRem[23][1]  = a[23];
  assign \u_div/PartRem[24][1]  = a[24];
  assign \u_div/PartRem[25][1]  = a[25];
  assign \u_div/PartRem[31][1]  = a[31];

  AND2X2 U1 ( .A(\u_div/CryTmp[2][16] ), .B(\u_div/PartRem[3][16] ), .Y(
        \u_div/CryTmp[2][17] ) );
  AND2X2 U2 ( .A(\u_div/CryTmp[1][16] ), .B(\u_div/PartRem[2][16] ), .Y(
        \u_div/CryTmp[1][17] ) );
  AND2X2 U3 ( .A(\u_div/CryTmp[3][16] ), .B(\u_div/PartRem[4][16] ), .Y(
        \u_div/CryTmp[3][17] ) );
  AND2X2 U4 ( .A(\u_div/CryTmp[4][16] ), .B(\u_div/PartRem[5][16] ), .Y(
        \u_div/CryTmp[4][17] ) );
  AND2X2 U5 ( .A(\u_div/CryTmp[5][16] ), .B(\u_div/PartRem[6][16] ), .Y(
        \u_div/CryTmp[5][17] ) );
  AND2X2 U6 ( .A(\u_div/CryTmp[6][16] ), .B(\u_div/PartRem[7][16] ), .Y(
        \u_div/CryTmp[6][17] ) );
  AND2X2 U7 ( .A(\u_div/CryTmp[7][16] ), .B(\u_div/PartRem[8][16] ), .Y(
        \u_div/CryTmp[7][17] ) );
  AND2X2 U8 ( .A(\u_div/CryTmp[8][16] ), .B(\u_div/PartRem[9][16] ), .Y(
        \u_div/CryTmp[8][17] ) );
  AND2X2 U9 ( .A(\u_div/CryTmp[9][16] ), .B(\u_div/PartRem[10][16] ), .Y(
        \u_div/CryTmp[9][17] ) );
  MX2X1 U10 ( .A(\u_div/PartRem[20][1] ), .B(n261), .S0(\u_div/CryTmp[15][17] ), .Y(n1) );
  MX2X1 U11 ( .A(n61), .B(n61), .S0(n275), .Y(n2) );
  MX2X1 U12 ( .A(n62), .B(n62), .S0(n276), .Y(n3) );
  MX2X1 U13 ( .A(n63), .B(n63), .S0(n271), .Y(n4) );
  MX2X1 U14 ( .A(n64), .B(n64), .S0(n266), .Y(n5) );
  MX2X1 U15 ( .A(n65), .B(n65), .S0(n267), .Y(n6) );
  MX2X1 U16 ( .A(n66), .B(n66), .S0(n263), .Y(n7) );
  MX2X1 U17 ( .A(\u_div/CryTmp[11][6] ), .B(n258), .S0(n275), .Y(n8) );
  MX2X1 U18 ( .A(\u_div/CryTmp[9][6] ), .B(n260), .S0(n271), .Y(n9) );
  MX2X1 U19 ( .A(\u_div/CryTmp[7][6] ), .B(n247), .S0(n266), .Y(n10) );
  MX2X1 U20 ( .A(\u_div/CryTmp[6][6] ), .B(n248), .S0(n263), .Y(n11) );
  MX2X1 U21 ( .A(\u_div/CryTmp[8][6] ), .B(n246), .S0(n267), .Y(n12) );
  MX2X1 U22 ( .A(\u_div/CryTmp[13][6] ), .B(n256), .S0(n273), .Y(n13) );
  MX2X1 U23 ( .A(\u_div/CryTmp[4][6] ), .B(n243), .S0(n270), .Y(n14) );
  MX2X1 U24 ( .A(\u_div/CryTmp[5][6] ), .B(n249), .S0(n269), .Y(n15) );
  MX2X1 U25 ( .A(n235), .B(\u_div/CryTmp[1][6] ), .S0(n264), .Y(n16) );
  AND2X2 U26 ( .A(\u_div/PartRem[1][16] ), .B(n78), .Y(n17) );
  AND2X2 U27 ( .A(\u_div/PartRem[1][10] ), .B(n79), .Y(n18) );
  MX2X1 U28 ( .A(n90), .B(\u_div/SumTmp[3][7] ), .S0(n268), .Y(n19) );
  MX2X1 U29 ( .A(n89), .B(\u_div/SumTmp[11][7] ), .S0(n275), .Y(n20) );
  MX2X1 U30 ( .A(n91), .B(\u_div/SumTmp[4][7] ), .S0(n270), .Y(n21) );
  MX2X1 U31 ( .A(n92), .B(\u_div/SumTmp[13][7] ), .S0(n273), .Y(n22) );
  MX2X1 U32 ( .A(\u_div/PartRem[22][1] ), .B(\u_div/SumTmp[15][7] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n23) );
  MX2X1 U33 ( .A(n233), .B(n170), .S0(n264), .Y(n24) );
  MX2X1 U34 ( .A(n81), .B(\u_div/SumTmp[10][7] ), .S0(n276), .Y(n25) );
  MX2X1 U35 ( .A(n82), .B(\u_div/SumTmp[9][7] ), .S0(n271), .Y(n26) );
  MX2X1 U36 ( .A(n84), .B(\u_div/SumTmp[7][7] ), .S0(n266), .Y(n27) );
  MX2X1 U37 ( .A(n85), .B(\u_div/SumTmp[6][7] ), .S0(n263), .Y(n28) );
  MX2X1 U38 ( .A(n83), .B(\u_div/SumTmp[8][7] ), .S0(n267), .Y(n29) );
  MX2X1 U39 ( .A(n88), .B(\u_div/SumTmp[12][7] ), .S0(n274), .Y(n30) );
  MX2X1 U40 ( .A(n86), .B(\u_div/SumTmp[5][7] ), .S0(n269), .Y(n31) );
  MX2X1 U41 ( .A(n93), .B(\u_div/SumTmp[14][7] ), .S0(n272), .Y(n32) );
  MX2X1 U42 ( .A(n114), .B(\u_div/SumTmp[3][10] ), .S0(n268), .Y(n33) );
  MX2X1 U43 ( .A(n108), .B(\u_div/SumTmp[7][10] ), .S0(n266), .Y(n34) );
  MX2X1 U44 ( .A(n109), .B(\u_div/SumTmp[6][10] ), .S0(n263), .Y(n35) );
  MX2X1 U45 ( .A(n112), .B(\u_div/SumTmp[9][10] ), .S0(n271), .Y(n36) );
  MX2X1 U46 ( .A(n113), .B(\u_div/SumTmp[8][10] ), .S0(n267), .Y(n37) );
  MX2X1 U47 ( .A(n115), .B(\u_div/SumTmp[4][10] ), .S0(n270), .Y(n38) );
  MX2X1 U48 ( .A(n110), .B(\u_div/SumTmp[5][10] ), .S0(n269), .Y(n39) );
  MX2X1 U49 ( .A(n116), .B(\u_div/SumTmp[10][10] ), .S0(n276), .Y(n40) );
  MX2X1 U50 ( .A(n117), .B(\u_div/SumTmp[11][10] ), .S0(n275), .Y(n41) );
  MX2X1 U51 ( .A(n118), .B(\u_div/SumTmp[12][10] ), .S0(n274), .Y(n42) );
  MX2X1 U52 ( .A(n119), .B(\u_div/SumTmp[13][10] ), .S0(n273), .Y(n43) );
  MX2X1 U53 ( .A(n120), .B(\u_div/SumTmp[14][10] ), .S0(n272), .Y(n44) );
  MX2X1 U54 ( .A(n241), .B(n168), .S0(n264), .Y(n45) );
  MX2X1 U55 ( .A(n126), .B(\u_div/SumTmp[3][12] ), .S0(n268), .Y(n46) );
  MX2X1 U56 ( .A(n124), .B(\u_div/SumTmp[7][12] ), .S0(n266), .Y(n47) );
  MX2X1 U57 ( .A(n125), .B(\u_div/SumTmp[6][12] ), .S0(n263), .Y(n48) );
  MX2X1 U58 ( .A(n127), .B(\u_div/SumTmp[4][12] ), .S0(n270), .Y(n49) );
  MX2X1 U59 ( .A(n128), .B(\u_div/SumTmp[8][12] ), .S0(n267), .Y(n50) );
  MX2X1 U60 ( .A(n129), .B(\u_div/SumTmp[9][12] ), .S0(n271), .Y(n51) );
  MX2X1 U61 ( .A(n130), .B(\u_div/SumTmp[10][12] ), .S0(n276), .Y(n52) );
  MX2X1 U62 ( .A(n131), .B(\u_div/SumTmp[11][12] ), .S0(n275), .Y(n53) );
  MX2X1 U63 ( .A(n132), .B(\u_div/SumTmp[12][12] ), .S0(n274), .Y(n54) );
  MX2X1 U64 ( .A(n133), .B(\u_div/SumTmp[13][12] ), .S0(n273), .Y(n55) );
  MX2X1 U65 ( .A(n134), .B(\u_div/SumTmp[14][12] ), .S0(n272), .Y(n56) );
  MX2X1 U66 ( .A(n239), .B(n167), .S0(n264), .Y(n57) );
  MX2X1 U67 ( .A(n176), .B(n176), .S0(n273), .Y(n58) );
  MX2X1 U68 ( .A(\u_div/PartRem[18][1] ), .B(\u_div/PartRem[18][1] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n59) );
  MX2X1 U69 ( .A(n177), .B(n177), .S0(n268), .Y(n60) );
  MX2X1 U70 ( .A(n178), .B(n178), .S0(n274), .Y(n61) );
  MX2X1 U71 ( .A(n181), .B(n181), .S0(n275), .Y(n62) );
  MX2X1 U72 ( .A(n180), .B(n180), .S0(n276), .Y(n63) );
  MX2X1 U73 ( .A(n182), .B(n182), .S0(n267), .Y(n64) );
  MX2X1 U74 ( .A(n184), .B(n184), .S0(n271), .Y(n65) );
  MX2X1 U75 ( .A(n183), .B(n183), .S0(n266), .Y(n66) );
  MX2X1 U76 ( .A(n179), .B(n179), .S0(n273), .Y(n67) );
  MX2X1 U77 ( .A(a[17]), .B(a[17]), .S0(\u_div/CryTmp[15][17] ), .Y(n68) );
  MX2X1 U78 ( .A(n185), .B(n185), .S0(n269), .Y(n69) );
  MX2X1 U79 ( .A(n186), .B(n186), .S0(n263), .Y(n70) );
  MX2X1 U80 ( .A(n187), .B(n187), .S0(n268), .Y(n71) );
  MX2X1 U81 ( .A(a[16]), .B(a[16]), .S0(\u_div/CryTmp[15][17] ), .Y(n72) );
  MX2X1 U82 ( .A(n188), .B(n188), .S0(n269), .Y(n73) );
  MX2X1 U83 ( .A(\u_div/CryTmp[10][6] ), .B(n259), .S0(n276), .Y(n74) );
  MX2X1 U84 ( .A(\u_div/CryTmp[3][6] ), .B(n244), .S0(n268), .Y(n75) );
  MX2X1 U85 ( .A(\u_div/CryTmp[12][6] ), .B(n257), .S0(n274), .Y(n76) );
  MX2X1 U86 ( .A(\u_div/CryTmp[14][6] ), .B(n262), .S0(n272), .Y(n77) );
  AND2X2 U87 ( .A(\u_div/PartRem[1][15] ), .B(\u_div/CryTmp[0][15] ), .Y(n78)
         );
  AND2X2 U88 ( .A(\u_div/PartRem[1][9] ), .B(\u_div/CryTmp[0][9] ), .Y(n79) );
  AND2X2 U89 ( .A(\u_div/PartRem[1][7] ), .B(\u_div/CryTmp[0][7] ), .Y(n80) );
  MX2X1 U90 ( .A(n76), .B(\u_div/SumTmp[11][6] ), .S0(n275), .Y(n81) );
  MX2X1 U91 ( .A(n8), .B(\u_div/SumTmp[10][6] ), .S0(n276), .Y(n82) );
  MX2X1 U92 ( .A(n74), .B(\u_div/SumTmp[9][6] ), .S0(n271), .Y(n83) );
  MX2X1 U93 ( .A(n9), .B(\u_div/SumTmp[8][6] ), .S0(n267), .Y(n84) );
  MX2X1 U94 ( .A(n12), .B(\u_div/SumTmp[7][6] ), .S0(n266), .Y(n85) );
  MX2X1 U95 ( .A(n10), .B(\u_div/SumTmp[6][6] ), .S0(n263), .Y(n86) );
  MX2X1 U96 ( .A(n14), .B(\u_div/SumTmp[3][6] ), .S0(n268), .Y(n87) );
  MX2X1 U97 ( .A(n77), .B(\u_div/SumTmp[13][6] ), .S0(n273), .Y(n88) );
  MX2X1 U98 ( .A(n13), .B(\u_div/SumTmp[12][6] ), .S0(n274), .Y(n89) );
  MX2X1 U99 ( .A(n15), .B(\u_div/SumTmp[4][6] ), .S0(n270), .Y(n90) );
  MX2X1 U100 ( .A(n11), .B(\u_div/SumTmp[5][6] ), .S0(n269), .Y(n91) );
  MX2X1 U101 ( .A(n1), .B(\u_div/SumTmp[14][6] ), .S0(n272), .Y(n92) );
  MX2X1 U102 ( .A(\u_div/PartRem[21][1] ), .B(\u_div/SumTmp[15][6] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n93) );
  MX2X1 U103 ( .A(n25), .B(\u_div/SumTmp[9][8] ), .S0(n271), .Y(n94) );
  MX2X1 U104 ( .A(n29), .B(\u_div/SumTmp[7][8] ), .S0(n266), .Y(n95) );
  MX2X1 U105 ( .A(n27), .B(\u_div/SumTmp[6][8] ), .S0(n263), .Y(n96) );
  MX2X1 U106 ( .A(n26), .B(\u_div/SumTmp[8][8] ), .S0(n267), .Y(n97) );
  MX2X1 U107 ( .A(n21), .B(\u_div/SumTmp[3][8] ), .S0(n268), .Y(n98) );
  MX2X1 U108 ( .A(n30), .B(\u_div/SumTmp[11][8] ), .S0(n275), .Y(n99) );
  MX2X1 U109 ( .A(n20), .B(\u_div/SumTmp[10][8] ), .S0(n276), .Y(n100) );
  MX2X1 U110 ( .A(n31), .B(\u_div/SumTmp[4][8] ), .S0(n270), .Y(n101) );
  MX2X1 U111 ( .A(n28), .B(\u_div/SumTmp[5][8] ), .S0(n269), .Y(n102) );
  MX2X1 U112 ( .A(n22), .B(\u_div/SumTmp[12][8] ), .S0(n274), .Y(n103) );
  MX2X1 U113 ( .A(n32), .B(\u_div/SumTmp[13][8] ), .S0(n273), .Y(n104) );
  MX2X1 U114 ( .A(n23), .B(\u_div/SumTmp[14][8] ), .S0(n272), .Y(n105) );
  MX2X1 U115 ( .A(\u_div/PartRem[23][1] ), .B(\u_div/SumTmp[15][8] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n106) );
  MX2X1 U116 ( .A(\u_div/PartRem[25][1] ), .B(\u_div/SumTmp[15][10] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n107) );
  MX2X1 U117 ( .A(n94), .B(\u_div/SumTmp[8][9] ), .S0(n267), .Y(n108) );
  MX2X1 U118 ( .A(n97), .B(\u_div/SumTmp[7][9] ), .S0(n266), .Y(n109) );
  MX2X1 U119 ( .A(n95), .B(\u_div/SumTmp[6][9] ), .S0(n263), .Y(n110) );
  MX2X1 U120 ( .A(n101), .B(\u_div/SumTmp[3][9] ), .S0(n268), .Y(n111) );
  MX2X1 U121 ( .A(n99), .B(\u_div/SumTmp[10][9] ), .S0(n276), .Y(n112) );
  MX2X1 U122 ( .A(n100), .B(\u_div/SumTmp[9][9] ), .S0(n271), .Y(n113) );
  MX2X1 U123 ( .A(n102), .B(\u_div/SumTmp[4][9] ), .S0(n270), .Y(n114) );
  MX2X1 U124 ( .A(n96), .B(\u_div/SumTmp[5][9] ), .S0(n269), .Y(n115) );
  MX2X1 U125 ( .A(n103), .B(\u_div/SumTmp[11][9] ), .S0(n275), .Y(n116) );
  MX2X1 U126 ( .A(n104), .B(\u_div/SumTmp[12][9] ), .S0(n274), .Y(n117) );
  MX2X1 U127 ( .A(n105), .B(\u_div/SumTmp[13][9] ), .S0(n273), .Y(n118) );
  MX2X1 U128 ( .A(n106), .B(\u_div/SumTmp[14][9] ), .S0(n272), .Y(n119) );
  MX2X1 U129 ( .A(\u_div/PartRem[24][1] ), .B(\u_div/SumTmp[15][9] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n120) );
  MX2X1 U130 ( .A(n34), .B(\u_div/SumTmp[6][11] ), .S0(n263), .Y(n121) );
  MX2X1 U131 ( .A(n121), .B(\u_div/SumTmp[5][12] ), .S0(n269), .Y(n122) );
  MX2X1 U132 ( .A(n38), .B(\u_div/SumTmp[3][11] ), .S0(n268), .Y(n123) );
  MX2X1 U133 ( .A(n36), .B(\u_div/SumTmp[8][11] ), .S0(n267), .Y(n124) );
  MX2X1 U134 ( .A(n37), .B(\u_div/SumTmp[7][11] ), .S0(n266), .Y(n125) );
  MX2X1 U135 ( .A(n39), .B(\u_div/SumTmp[4][11] ), .S0(n270), .Y(n126) );
  MX2X1 U136 ( .A(n35), .B(\u_div/SumTmp[5][11] ), .S0(n269), .Y(n127) );
  MX2X1 U137 ( .A(n40), .B(\u_div/SumTmp[9][11] ), .S0(n271), .Y(n128) );
  MX2X1 U138 ( .A(n41), .B(\u_div/SumTmp[10][11] ), .S0(n276), .Y(n129) );
  MX2X1 U139 ( .A(n42), .B(\u_div/SumTmp[11][11] ), .S0(n275), .Y(n130) );
  MX2X1 U140 ( .A(n43), .B(\u_div/SumTmp[12][11] ), .S0(n274), .Y(n131) );
  MX2X1 U141 ( .A(n44), .B(\u_div/SumTmp[13][11] ), .S0(n273), .Y(n132) );
  MX2X1 U142 ( .A(n107), .B(\u_div/SumTmp[14][11] ), .S0(n272), .Y(n133) );
  MX2X1 U143 ( .A(a[26]), .B(\u_div/SumTmp[15][11] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n134) );
  MX2X1 U144 ( .A(a[27]), .B(\u_div/SumTmp[15][12] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n135) );
  MX2X1 U145 ( .A(n242), .B(n198), .S0(n264), .Y(n136) );
  MX2X1 U146 ( .A(n49), .B(\u_div/SumTmp[3][13] ), .S0(n268), .Y(n137) );
  MX2X1 U147 ( .A(n47), .B(\u_div/SumTmp[6][13] ), .S0(n263), .Y(n138) );
  MX2X1 U148 ( .A(n122), .B(\u_div/SumTmp[4][13] ), .S0(n270), .Y(n139) );
  MX2X1 U149 ( .A(n48), .B(\u_div/SumTmp[5][13] ), .S0(n269), .Y(n140) );
  MX2X1 U150 ( .A(n50), .B(\u_div/SumTmp[7][13] ), .S0(n266), .Y(n141) );
  MX2X1 U151 ( .A(n51), .B(\u_div/SumTmp[8][13] ), .S0(n267), .Y(n142) );
  MX2X1 U152 ( .A(n52), .B(\u_div/SumTmp[9][13] ), .S0(n271), .Y(n143) );
  MX2X1 U153 ( .A(n53), .B(\u_div/SumTmp[10][13] ), .S0(n276), .Y(n144) );
  MX2X1 U154 ( .A(n54), .B(\u_div/SumTmp[11][13] ), .S0(n275), .Y(n145) );
  MX2X1 U155 ( .A(n55), .B(\u_div/SumTmp[12][13] ), .S0(n274), .Y(n146) );
  MX2X1 U156 ( .A(n56), .B(\u_div/SumTmp[13][13] ), .S0(n273), .Y(n147) );
  MX2X1 U157 ( .A(n135), .B(\u_div/SumTmp[14][13] ), .S0(n272), .Y(n148) );
  MX2X1 U158 ( .A(a[28]), .B(\u_div/SumTmp[15][13] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n149) );
  MX2X1 U159 ( .A(n240), .B(n195), .S0(n264), .Y(n150) );
  MX2X1 U160 ( .A(n138), .B(\u_div/SumTmp[5][14] ), .S0(n269), .Y(n151) );
  MX2X1 U161 ( .A(n140), .B(\u_div/SumTmp[4][14] ), .S0(n270), .Y(n152) );
  MX2X1 U162 ( .A(n139), .B(\u_div/SumTmp[3][14] ), .S0(n268), .Y(n153) );
  MX2X1 U163 ( .A(n141), .B(\u_div/SumTmp[6][14] ), .S0(n263), .Y(n154) );
  MX2X1 U164 ( .A(n142), .B(\u_div/SumTmp[7][14] ), .S0(n266), .Y(n155) );
  MX2X1 U165 ( .A(n143), .B(\u_div/SumTmp[8][14] ), .S0(n267), .Y(n156) );
  MX2X1 U166 ( .A(n144), .B(\u_div/SumTmp[9][14] ), .S0(n271), .Y(n157) );
  MX2X1 U167 ( .A(n145), .B(\u_div/SumTmp[10][14] ), .S0(n276), .Y(n158) );
  MX2X1 U168 ( .A(n146), .B(\u_div/SumTmp[11][14] ), .S0(n275), .Y(n159) );
  MX2X1 U169 ( .A(n147), .B(\u_div/SumTmp[12][14] ), .S0(n274), .Y(n160) );
  MX2X1 U170 ( .A(n148), .B(\u_div/SumTmp[13][14] ), .S0(n273), .Y(n161) );
  MX2X1 U171 ( .A(n149), .B(\u_div/SumTmp[14][14] ), .S0(n272), .Y(n162) );
  MX2X1 U172 ( .A(a[29]), .B(\u_div/SumTmp[15][14] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n163) );
  MX2X1 U173 ( .A(n236), .B(n189), .S0(n264), .Y(n164) );
  MX2X1 U174 ( .A(n67), .B(n67), .S0(n274), .Y(n165) );
  MX2X1 U175 ( .A(n68), .B(n68), .S0(n272), .Y(n166) );
  XOR2X1 U176 ( .A(\u_div/PartRem[2][13] ), .B(\u_div/CryTmp[1][13] ), .Y(n167) );
  XOR2X1 U177 ( .A(\u_div/PartRem[2][11] ), .B(\u_div/CryTmp[1][11] ), .Y(n168) );
  XOR2X1 U178 ( .A(\u_div/PartRem[2][8] ), .B(\u_div/CryTmp[1][8] ), .Y(n169)
         );
  XNOR2X1 U179 ( .A(\u_div/PartRem[2][7] ), .B(\u_div/CryTmp[1][7] ), .Y(n170)
         );
  MX2X1 U180 ( .A(n69), .B(n69), .S0(n270), .Y(n171) );
  MX2X1 U181 ( .A(n70), .B(n70), .S0(n269), .Y(n172) );
  XOR2X1 U182 ( .A(\u_div/PartRem[2][14] ), .B(\u_div/CryTmp[1][14] ), .Y(n173) );
  XNOR2X1 U183 ( .A(\u_div/PartRem[2][15] ), .B(\u_div/CryTmp[1][15] ), .Y(
        n174) );
  XNOR2X1 U184 ( .A(\u_div/PartRem[2][9] ), .B(\u_div/CryTmp[1][9] ), .Y(n175)
         );
  MX2X1 U185 ( .A(n72), .B(n72), .S0(n272), .Y(n176) );
  MX2X1 U186 ( .A(n73), .B(n73), .S0(n270), .Y(n177) );
  MX2X1 U187 ( .A(n212), .B(n212), .S0(n273), .Y(n178) );
  MX2X1 U188 ( .A(n213), .B(n213), .S0(n272), .Y(n179) );
  MX2X1 U189 ( .A(n219), .B(n219), .S0(n275), .Y(n180) );
  MX2X1 U190 ( .A(n220), .B(n220), .S0(n274), .Y(n181) );
  MX2X1 U191 ( .A(n215), .B(n215), .S0(n271), .Y(n182) );
  MX2X1 U192 ( .A(n221), .B(n221), .S0(n267), .Y(n183) );
  MX2X1 U193 ( .A(n218), .B(n218), .S0(n276), .Y(n184) );
  MX2X1 U194 ( .A(n216), .B(n216), .S0(n263), .Y(n185) );
  MX2X1 U195 ( .A(n222), .B(n222), .S0(n266), .Y(n186) );
  MX2X1 U196 ( .A(n217), .B(n217), .S0(n270), .Y(n187) );
  MX2X1 U197 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[6][0] ), .S0(n263), 
        .Y(n188) );
  AND2X2 U198 ( .A(\u_div/CryTmp[10][16] ), .B(\u_div/PartRem[11][16] ), .Y(
        \u_div/CryTmp[10][17] ) );
  AND2X2 U199 ( .A(\u_div/CryTmp[11][16] ), .B(\u_div/PartRem[12][16] ), .Y(
        \u_div/CryTmp[11][17] ) );
  AND2X2 U200 ( .A(\u_div/CryTmp[12][16] ), .B(\u_div/PartRem[13][16] ), .Y(
        \u_div/CryTmp[12][17] ) );
  AND2X2 U201 ( .A(\u_div/CryTmp[13][16] ), .B(\u_div/PartRem[14][16] ), .Y(
        \u_div/CryTmp[13][17] ) );
  AND2X2 U202 ( .A(\u_div/CryTmp[14][16] ), .B(\u_div/PartRem[15][16] ), .Y(
        \u_div/CryTmp[14][17] ) );
  BUFX3 U203 ( .A(quotient[2]), .Y(n265) );
  BUFX3 U204 ( .A(quotient[1]), .Y(n264) );
  XNOR2X1 U205 ( .A(\u_div/PartRem[2][16] ), .B(\u_div/CryTmp[1][16] ), .Y(
        n189) );
  OR2X2 U206 ( .A(\u_div/CryTmp[1][17] ), .B(\u_div/PartRem[2][17] ), .Y(
        quotient[1]) );
  MXI2X1 U207 ( .A(n230), .B(n192), .S0(n265), .Y(\u_div/PartRem[2][17] ) );
  OR2X2 U208 ( .A(\u_div/CryTmp[2][17] ), .B(\u_div/PartRem[3][17] ), .Y(
        quotient[2]) );
  MXI2X1 U209 ( .A(n229), .B(n191), .S0(n268), .Y(\u_div/PartRem[3][17] ) );
  BUFX3 U210 ( .A(quotient[3]), .Y(n268) );
  AND2X2 U211 ( .A(\u_div/CryTmp[1][15] ), .B(\u_div/PartRem[2][15] ), .Y(
        \u_div/CryTmp[1][16] ) );
  INVX1 U212 ( .A(n229), .Y(\u_div/PartRem[4][16] ) );
  INVX1 U213 ( .A(n230), .Y(\u_div/PartRem[3][16] ) );
  INVX1 U214 ( .A(n236), .Y(\u_div/PartRem[2][16] ) );
  XNOR2X1 U215 ( .A(\u_div/PartRem[5][16] ), .B(\u_div/CryTmp[4][16] ), .Y(
        n190) );
  XNOR2X1 U216 ( .A(\u_div/PartRem[4][16] ), .B(\u_div/CryTmp[3][16] ), .Y(
        n191) );
  XNOR2X1 U217 ( .A(\u_div/PartRem[3][16] ), .B(\u_div/CryTmp[2][16] ), .Y(
        n192) );
  OR2X2 U218 ( .A(\u_div/CryTmp[3][17] ), .B(\u_div/PartRem[4][17] ), .Y(
        quotient[3]) );
  MXI2X1 U219 ( .A(n228), .B(n190), .S0(n270), .Y(\u_div/PartRem[4][17] ) );
  BUFX3 U220 ( .A(quotient[4]), .Y(n270) );
  AND2X2 U221 ( .A(\u_div/CryTmp[4][15] ), .B(n151), .Y(\u_div/CryTmp[4][16] )
         );
  AND2X2 U222 ( .A(\u_div/CryTmp[3][15] ), .B(n152), .Y(\u_div/CryTmp[3][16] )
         );
  AND2X2 U223 ( .A(\u_div/CryTmp[2][15] ), .B(n153), .Y(\u_div/CryTmp[2][16] )
         );
  OR2X2 U224 ( .A(\u_div/CryTmp[1][14] ), .B(\u_div/PartRem[2][14] ), .Y(
        \u_div/CryTmp[1][15] ) );
  MXI2X1 U225 ( .A(n151), .B(\u_div/SumTmp[4][15] ), .S0(n270), .Y(n229) );
  XOR2X1 U226 ( .A(n151), .B(\u_div/CryTmp[4][15] ), .Y(\u_div/SumTmp[4][15] )
         );
  MXI2X1 U227 ( .A(n152), .B(\u_div/SumTmp[3][15] ), .S0(n268), .Y(n230) );
  XOR2X1 U228 ( .A(n152), .B(\u_div/CryTmp[3][15] ), .Y(\u_div/SumTmp[3][15] )
         );
  MXI2X1 U229 ( .A(n153), .B(\u_div/SumTmp[2][15] ), .S0(n265), .Y(n236) );
  XOR2X1 U230 ( .A(n153), .B(\u_div/CryTmp[2][15] ), .Y(\u_div/SumTmp[2][15] )
         );
  INVX1 U231 ( .A(n228), .Y(\u_div/PartRem[5][16] ) );
  INVX1 U232 ( .A(n237), .Y(\u_div/PartRem[2][15] ) );
  XNOR2X1 U233 ( .A(\u_div/PartRem[6][16] ), .B(\u_div/CryTmp[5][16] ), .Y(
        n193) );
  OR2X2 U234 ( .A(\u_div/CryTmp[4][17] ), .B(\u_div/PartRem[5][17] ), .Y(
        quotient[4]) );
  MXI2X1 U235 ( .A(n227), .B(n193), .S0(n269), .Y(\u_div/PartRem[5][17] ) );
  BUFX4 U236 ( .A(quotient[5]), .Y(n269) );
  AND2X2 U237 ( .A(\u_div/CryTmp[5][15] ), .B(n154), .Y(\u_div/CryTmp[5][16] )
         );
  OR2X2 U238 ( .A(\u_div/CryTmp[1][13] ), .B(\u_div/PartRem[2][13] ), .Y(
        \u_div/CryTmp[1][14] ) );
  OR2X2 U239 ( .A(\u_div/CryTmp[5][14] ), .B(n138), .Y(\u_div/CryTmp[5][15] )
         );
  OR2X2 U240 ( .A(\u_div/CryTmp[4][14] ), .B(n140), .Y(\u_div/CryTmp[4][15] )
         );
  OR2X2 U241 ( .A(\u_div/CryTmp[3][14] ), .B(n139), .Y(\u_div/CryTmp[3][15] )
         );
  OR2X2 U242 ( .A(\u_div/CryTmp[2][14] ), .B(n137), .Y(\u_div/CryTmp[2][15] )
         );
  NAND2BX1 U243 ( .AN(n17), .B(n164), .Y(quotient[0]) );
  MXI2X1 U244 ( .A(n154), .B(\u_div/SumTmp[5][15] ), .S0(n269), .Y(n228) );
  XOR2X1 U245 ( .A(n154), .B(\u_div/CryTmp[5][15] ), .Y(\u_div/SumTmp[5][15] )
         );
  MXI2X1 U246 ( .A(n137), .B(\u_div/SumTmp[2][14] ), .S0(n265), .Y(n237) );
  XNOR2X1 U247 ( .A(n137), .B(\u_div/CryTmp[2][14] ), .Y(\u_div/SumTmp[2][14] ) );
  XNOR2X1 U248 ( .A(n138), .B(\u_div/CryTmp[5][14] ), .Y(\u_div/SumTmp[5][14] ) );
  XNOR2X1 U249 ( .A(n139), .B(\u_div/CryTmp[3][14] ), .Y(\u_div/SumTmp[3][14] ) );
  XNOR2X1 U250 ( .A(n140), .B(\u_div/CryTmp[4][14] ), .Y(\u_div/SumTmp[4][14] ) );
  INVX1 U251 ( .A(n227), .Y(\u_div/PartRem[6][16] ) );
  INVX1 U252 ( .A(n238), .Y(\u_div/PartRem[2][14] ) );
  XNOR2X1 U253 ( .A(\u_div/PartRem[7][16] ), .B(\u_div/CryTmp[6][16] ), .Y(
        n194) );
  BUFX4 U254 ( .A(quotient[6]), .Y(n263) );
  AND2X2 U255 ( .A(\u_div/CryTmp[6][15] ), .B(n155), .Y(\u_div/CryTmp[6][16] )
         );
  OR2X2 U256 ( .A(\u_div/CryTmp[6][13] ), .B(n47), .Y(\u_div/CryTmp[6][14] )
         );
  OR2X2 U257 ( .A(\u_div/CryTmp[5][12] ), .B(n121), .Y(\u_div/CryTmp[5][13] )
         );
  OR2X2 U258 ( .A(\u_div/CryTmp[5][13] ), .B(n48), .Y(\u_div/CryTmp[5][14] )
         );
  OR2X2 U259 ( .A(\u_div/CryTmp[4][13] ), .B(n122), .Y(\u_div/CryTmp[4][14] )
         );
  OR2X2 U260 ( .A(\u_div/CryTmp[3][13] ), .B(n49), .Y(\u_div/CryTmp[3][14] )
         );
  OR2X2 U261 ( .A(\u_div/CryTmp[2][13] ), .B(n46), .Y(\u_div/CryTmp[2][14] )
         );
  OR2X2 U262 ( .A(\u_div/CryTmp[1][12] ), .B(\u_div/PartRem[2][12] ), .Y(
        \u_div/CryTmp[1][13] ) );
  OR2X2 U263 ( .A(\u_div/CryTmp[6][14] ), .B(n141), .Y(\u_div/CryTmp[6][15] )
         );
  MXI2X1 U264 ( .A(n237), .B(n174), .S0(n264), .Y(\u_div/PartRem[1][16] ) );
  OR2X2 U265 ( .A(\u_div/CryTmp[5][17] ), .B(\u_div/PartRem[6][17] ), .Y(
        quotient[5]) );
  MXI2X1 U266 ( .A(n226), .B(n194), .S0(n263), .Y(\u_div/PartRem[6][17] ) );
  XNOR2X1 U267 ( .A(n121), .B(\u_div/CryTmp[5][12] ), .Y(\u_div/SumTmp[5][12] ) );
  INVX1 U268 ( .A(n239), .Y(\u_div/PartRem[2][13] ) );
  MXI2X1 U269 ( .A(n155), .B(\u_div/SumTmp[6][15] ), .S0(n263), .Y(n227) );
  XOR2X1 U270 ( .A(n155), .B(\u_div/CryTmp[6][15] ), .Y(\u_div/SumTmp[6][15] )
         );
  MXI2X1 U271 ( .A(n46), .B(\u_div/SumTmp[2][13] ), .S0(n265), .Y(n238) );
  XNOR2X1 U272 ( .A(n46), .B(\u_div/CryTmp[2][13] ), .Y(\u_div/SumTmp[2][13] )
         );
  XNOR2X1 U273 ( .A(n141), .B(\u_div/CryTmp[6][14] ), .Y(\u_div/SumTmp[6][14] ) );
  XNOR2X1 U274 ( .A(n47), .B(\u_div/CryTmp[6][13] ), .Y(\u_div/SumTmp[6][13] )
         );
  XNOR2X1 U275 ( .A(n48), .B(\u_div/CryTmp[5][13] ), .Y(\u_div/SumTmp[5][13] )
         );
  XNOR2X1 U276 ( .A(n49), .B(\u_div/CryTmp[3][13] ), .Y(\u_div/SumTmp[3][13] )
         );
  XNOR2X1 U277 ( .A(n122), .B(\u_div/CryTmp[4][13] ), .Y(\u_div/SumTmp[4][13] ) );
  INVX1 U278 ( .A(n226), .Y(\u_div/PartRem[7][16] ) );
  XOR2X1 U279 ( .A(\u_div/PartRem[2][12] ), .B(\u_div/CryTmp[1][12] ), .Y(n195) );
  XNOR2X1 U280 ( .A(\u_div/PartRem[8][16] ), .B(\u_div/CryTmp[7][16] ), .Y(
        n196) );
  OR2X2 U281 ( .A(\u_div/CryTmp[6][17] ), .B(\u_div/PartRem[7][17] ), .Y(
        quotient[6]) );
  MXI2X1 U282 ( .A(n225), .B(n196), .S0(n266), .Y(\u_div/PartRem[7][17] ) );
  BUFX4 U283 ( .A(quotient[7]), .Y(n266) );
  AND2X2 U284 ( .A(\u_div/CryTmp[7][15] ), .B(n156), .Y(\u_div/CryTmp[7][16] )
         );
  OR2X2 U285 ( .A(\u_div/CryTmp[7][12] ), .B(n124), .Y(\u_div/CryTmp[7][13] )
         );
  OR2X2 U286 ( .A(\u_div/CryTmp[7][13] ), .B(n50), .Y(\u_div/CryTmp[7][14] )
         );
  OR2X2 U287 ( .A(\u_div/CryTmp[6][11] ), .B(n34), .Y(\u_div/CryTmp[6][12] )
         );
  OR2X2 U288 ( .A(\u_div/CryTmp[6][12] ), .B(n125), .Y(\u_div/CryTmp[6][13] )
         );
  OR2X2 U289 ( .A(\u_div/CryTmp[5][11] ), .B(n35), .Y(\u_div/CryTmp[5][12] )
         );
  OR2X2 U290 ( .A(\u_div/CryTmp[4][12] ), .B(n127), .Y(\u_div/CryTmp[4][13] )
         );
  OR2X2 U291 ( .A(\u_div/CryTmp[3][12] ), .B(n126), .Y(\u_div/CryTmp[3][13] )
         );
  OR2X2 U292 ( .A(\u_div/CryTmp[2][12] ), .B(n123), .Y(\u_div/CryTmp[2][13] )
         );
  OR2X2 U293 ( .A(\u_div/CryTmp[1][11] ), .B(\u_div/PartRem[2][11] ), .Y(
        \u_div/CryTmp[1][12] ) );
  OR2X2 U294 ( .A(\u_div/CryTmp[7][14] ), .B(n142), .Y(\u_div/CryTmp[7][15] )
         );
  MXI2X1 U295 ( .A(n238), .B(n173), .S0(n264), .Y(\u_div/PartRem[1][15] ) );
  NAND2BX1 U296 ( .AN(\u_div/CryTmp[0][14] ), .B(n57), .Y(
        \u_div/CryTmp[0][15] ) );
  MXI2X1 U297 ( .A(n123), .B(\u_div/SumTmp[2][12] ), .S0(n265), .Y(n239) );
  XNOR2X1 U298 ( .A(n123), .B(\u_div/CryTmp[2][12] ), .Y(\u_div/SumTmp[2][12] ) );
  XNOR2X1 U299 ( .A(n124), .B(\u_div/CryTmp[7][12] ), .Y(\u_div/SumTmp[7][12] ) );
  XNOR2X1 U300 ( .A(n34), .B(\u_div/CryTmp[6][11] ), .Y(\u_div/SumTmp[6][11] )
         );
  XNOR2X1 U301 ( .A(n125), .B(\u_div/CryTmp[6][12] ), .Y(\u_div/SumTmp[6][12] ) );
  XNOR2X1 U302 ( .A(n35), .B(\u_div/CryTmp[5][11] ), .Y(\u_div/SumTmp[5][11] )
         );
  XNOR2X1 U303 ( .A(n126), .B(\u_div/CryTmp[3][12] ), .Y(\u_div/SumTmp[3][12] ) );
  XNOR2X1 U304 ( .A(n127), .B(\u_div/CryTmp[4][12] ), .Y(\u_div/SumTmp[4][12] ) );
  INVX1 U305 ( .A(n240), .Y(\u_div/PartRem[2][12] ) );
  MXI2X1 U306 ( .A(n156), .B(\u_div/SumTmp[7][15] ), .S0(n266), .Y(n226) );
  XOR2X1 U307 ( .A(n156), .B(\u_div/CryTmp[7][15] ), .Y(\u_div/SumTmp[7][15] )
         );
  XNOR2X1 U308 ( .A(n50), .B(\u_div/CryTmp[7][13] ), .Y(\u_div/SumTmp[7][13] )
         );
  XNOR2X1 U309 ( .A(n142), .B(\u_div/CryTmp[7][14] ), .Y(\u_div/SumTmp[7][14] ) );
  INVX1 U310 ( .A(n225), .Y(\u_div/PartRem[8][16] ) );
  XNOR2X1 U311 ( .A(\u_div/PartRem[9][16] ), .B(\u_div/CryTmp[8][16] ), .Y(
        n197) );
  OR2X2 U312 ( .A(\u_div/CryTmp[7][17] ), .B(\u_div/PartRem[8][17] ), .Y(
        quotient[7]) );
  MXI2X1 U313 ( .A(n224), .B(n197), .S0(n267), .Y(\u_div/PartRem[8][17] ) );
  BUFX4 U314 ( .A(quotient[8]), .Y(n267) );
  AND2X2 U315 ( .A(\u_div/CryTmp[7][10] ), .B(n108), .Y(\u_div/CryTmp[7][11] )
         );
  AND2X2 U316 ( .A(\u_div/CryTmp[6][10] ), .B(n109), .Y(\u_div/CryTmp[6][11] )
         );
  AND2X2 U317 ( .A(\u_div/CryTmp[5][10] ), .B(n110), .Y(\u_div/CryTmp[5][11] )
         );
  AND2X2 U318 ( .A(\u_div/CryTmp[1][10] ), .B(\u_div/PartRem[2][10] ), .Y(
        \u_div/CryTmp[1][11] ) );
  AND2X2 U319 ( .A(\u_div/CryTmp[8][15] ), .B(n157), .Y(\u_div/CryTmp[8][16] )
         );
  OR2X2 U320 ( .A(\u_div/CryTmp[8][11] ), .B(n36), .Y(\u_div/CryTmp[8][12] )
         );
  OR2X2 U321 ( .A(\u_div/CryTmp[8][12] ), .B(n128), .Y(\u_div/CryTmp[8][13] )
         );
  OR2X2 U322 ( .A(\u_div/CryTmp[8][13] ), .B(n51), .Y(\u_div/CryTmp[8][14] )
         );
  OR2X2 U323 ( .A(\u_div/CryTmp[7][11] ), .B(n37), .Y(\u_div/CryTmp[7][12] )
         );
  OR2X2 U324 ( .A(\u_div/CryTmp[4][11] ), .B(n39), .Y(\u_div/CryTmp[4][12] )
         );
  OR2X2 U325 ( .A(\u_div/CryTmp[3][11] ), .B(n38), .Y(\u_div/CryTmp[3][12] )
         );
  OR2X2 U326 ( .A(\u_div/CryTmp[2][11] ), .B(n33), .Y(\u_div/CryTmp[2][12] )
         );
  OR2X2 U327 ( .A(\u_div/CryTmp[8][14] ), .B(n143), .Y(\u_div/CryTmp[8][15] )
         );
  NAND2BX1 U328 ( .AN(\u_div/CryTmp[0][13] ), .B(n150), .Y(
        \u_div/CryTmp[0][14] ) );
  NAND2BX1 U329 ( .AN(\u_div/CryTmp[0][12] ), .B(n45), .Y(
        \u_div/CryTmp[0][13] ) );
  XOR2X1 U330 ( .A(n108), .B(\u_div/CryTmp[7][10] ), .Y(\u_div/SumTmp[7][10] )
         );
  XOR2X1 U331 ( .A(n109), .B(\u_div/CryTmp[6][10] ), .Y(\u_div/SumTmp[6][10] )
         );
  XOR2X1 U332 ( .A(n110), .B(\u_div/CryTmp[5][10] ), .Y(\u_div/SumTmp[5][10] )
         );
  INVX1 U333 ( .A(n241), .Y(\u_div/PartRem[2][11] ) );
  MXI2X1 U334 ( .A(n33), .B(\u_div/SumTmp[2][11] ), .S0(n265), .Y(n240) );
  XNOR2X1 U335 ( .A(n33), .B(\u_div/CryTmp[2][11] ), .Y(\u_div/SumTmp[2][11] )
         );
  XNOR2X1 U336 ( .A(n36), .B(\u_div/CryTmp[8][11] ), .Y(\u_div/SumTmp[8][11] )
         );
  XNOR2X1 U337 ( .A(n128), .B(\u_div/CryTmp[8][12] ), .Y(\u_div/SumTmp[8][12] ) );
  XNOR2X1 U338 ( .A(n37), .B(\u_div/CryTmp[7][11] ), .Y(\u_div/SumTmp[7][11] )
         );
  XNOR2X1 U339 ( .A(n38), .B(\u_div/CryTmp[3][11] ), .Y(\u_div/SumTmp[3][11] )
         );
  XNOR2X1 U340 ( .A(n39), .B(\u_div/CryTmp[4][11] ), .Y(\u_div/SumTmp[4][11] )
         );
  MXI2X1 U341 ( .A(n157), .B(\u_div/SumTmp[8][15] ), .S0(n267), .Y(n225) );
  XOR2X1 U342 ( .A(n157), .B(\u_div/CryTmp[8][15] ), .Y(\u_div/SumTmp[8][15] )
         );
  XNOR2X1 U343 ( .A(n143), .B(\u_div/CryTmp[8][14] ), .Y(\u_div/SumTmp[8][14] ) );
  XNOR2X1 U344 ( .A(n51), .B(\u_div/CryTmp[8][13] ), .Y(\u_div/SumTmp[8][13] )
         );
  INVX1 U345 ( .A(n224), .Y(\u_div/PartRem[9][16] ) );
  XNOR2X1 U346 ( .A(\u_div/PartRem[2][10] ), .B(\u_div/CryTmp[1][10] ), .Y(
        n198) );
  XNOR2X1 U347 ( .A(\u_div/PartRem[10][16] ), .B(\u_div/CryTmp[9][16] ), .Y(
        n199) );
  BUFX4 U348 ( .A(quotient[9]), .Y(n271) );
  AND2X2 U349 ( .A(\u_div/CryTmp[9][10] ), .B(n112), .Y(\u_div/CryTmp[9][11] )
         );
  AND2X2 U350 ( .A(\u_div/CryTmp[8][10] ), .B(n113), .Y(\u_div/CryTmp[8][11] )
         );
  AND2X2 U351 ( .A(\u_div/CryTmp[4][10] ), .B(n115), .Y(\u_div/CryTmp[4][11] )
         );
  AND2X2 U352 ( .A(\u_div/CryTmp[3][10] ), .B(n114), .Y(\u_div/CryTmp[3][11] )
         );
  AND2X2 U353 ( .A(\u_div/CryTmp[2][10] ), .B(n111), .Y(\u_div/CryTmp[2][11] )
         );
  AND2X2 U354 ( .A(\u_div/CryTmp[9][15] ), .B(n158), .Y(\u_div/CryTmp[9][16] )
         );
  AND2X2 U355 ( .A(\u_div/CryTmp[8][9] ), .B(n94), .Y(\u_div/CryTmp[8][10] )
         );
  AND2X2 U356 ( .A(\u_div/CryTmp[7][9] ), .B(n97), .Y(\u_div/CryTmp[7][10] )
         );
  AND2X2 U357 ( .A(\u_div/CryTmp[6][9] ), .B(n95), .Y(\u_div/CryTmp[6][10] )
         );
  AND2X2 U358 ( .A(\u_div/CryTmp[5][9] ), .B(n96), .Y(\u_div/CryTmp[5][10] )
         );
  OR2X2 U359 ( .A(\u_div/CryTmp[9][11] ), .B(n40), .Y(\u_div/CryTmp[9][12] )
         );
  OR2X2 U360 ( .A(\u_div/CryTmp[9][12] ), .B(n129), .Y(\u_div/CryTmp[9][13] )
         );
  OR2X2 U361 ( .A(\u_div/CryTmp[9][13] ), .B(n52), .Y(\u_div/CryTmp[9][14] )
         );
  AND2X2 U362 ( .A(\u_div/CryTmp[1][9] ), .B(\u_div/PartRem[2][9] ), .Y(
        \u_div/CryTmp[1][10] ) );
  OR2X2 U363 ( .A(\u_div/CryTmp[9][14] ), .B(n144), .Y(\u_div/CryTmp[9][15] )
         );
  NAND2BX1 U364 ( .AN(n18), .B(n136), .Y(\u_div/CryTmp[0][12] ) );
  OR2X2 U365 ( .A(\u_div/CryTmp[8][17] ), .B(\u_div/PartRem[9][17] ), .Y(
        quotient[8]) );
  MXI2X1 U366 ( .A(n223), .B(n199), .S0(n271), .Y(\u_div/PartRem[9][17] ) );
  MXI2X1 U367 ( .A(n111), .B(\u_div/SumTmp[2][10] ), .S0(n265), .Y(n241) );
  XOR2X1 U368 ( .A(n111), .B(\u_div/CryTmp[2][10] ), .Y(\u_div/SumTmp[2][10] )
         );
  XOR2X1 U369 ( .A(n94), .B(\u_div/CryTmp[8][9] ), .Y(\u_div/SumTmp[8][9] ) );
  XOR2X1 U370 ( .A(n95), .B(\u_div/CryTmp[6][9] ), .Y(\u_div/SumTmp[6][9] ) );
  XOR2X1 U371 ( .A(n96), .B(\u_div/CryTmp[5][9] ), .Y(\u_div/SumTmp[5][9] ) );
  XOR2X1 U372 ( .A(n112), .B(\u_div/CryTmp[9][10] ), .Y(\u_div/SumTmp[9][10] )
         );
  XOR2X1 U373 ( .A(n113), .B(\u_div/CryTmp[8][10] ), .Y(\u_div/SumTmp[8][10] )
         );
  XOR2X1 U374 ( .A(n114), .B(\u_div/CryTmp[3][10] ), .Y(\u_div/SumTmp[3][10] )
         );
  XOR2X1 U375 ( .A(n97), .B(\u_div/CryTmp[7][9] ), .Y(\u_div/SumTmp[7][9] ) );
  XOR2X1 U376 ( .A(n115), .B(\u_div/CryTmp[4][10] ), .Y(\u_div/SumTmp[4][10] )
         );
  INVX1 U377 ( .A(n242), .Y(\u_div/PartRem[2][10] ) );
  XNOR2X1 U378 ( .A(n40), .B(\u_div/CryTmp[9][11] ), .Y(\u_div/SumTmp[9][11] )
         );
  XNOR2X1 U379 ( .A(n129), .B(\u_div/CryTmp[9][12] ), .Y(\u_div/SumTmp[9][12] ) );
  MXI2X1 U380 ( .A(n158), .B(\u_div/SumTmp[9][15] ), .S0(n271), .Y(n224) );
  XOR2X1 U381 ( .A(n158), .B(\u_div/CryTmp[9][15] ), .Y(\u_div/SumTmp[9][15] )
         );
  XNOR2X1 U382 ( .A(n144), .B(\u_div/CryTmp[9][14] ), .Y(\u_div/SumTmp[9][14] ) );
  XNOR2X1 U383 ( .A(n52), .B(\u_div/CryTmp[9][13] ), .Y(\u_div/SumTmp[9][13] )
         );
  INVX1 U384 ( .A(n223), .Y(\u_div/PartRem[10][16] ) );
  XNOR2X1 U385 ( .A(\u_div/PartRem[11][16] ), .B(\u_div/CryTmp[10][16] ), .Y(
        n200) );
  OR2X2 U386 ( .A(\u_div/CryTmp[9][17] ), .B(\u_div/PartRem[10][17] ), .Y(
        quotient[9]) );
  MXI2X1 U387 ( .A(n255), .B(n200), .S0(n276), .Y(\u_div/PartRem[10][17] ) );
  AND2X2 U388 ( .A(\u_div/CryTmp[10][10] ), .B(n116), .Y(
        \u_div/CryTmp[10][11] ) );
  AND2X2 U389 ( .A(\u_div/CryTmp[1][7] ), .B(\u_div/PartRem[2][7] ), .Y(
        \u_div/CryTmp[1][8] ) );
  AND2X2 U390 ( .A(\u_div/CryTmp[10][9] ), .B(n99), .Y(\u_div/CryTmp[10][10] )
         );
  AND2X2 U391 ( .A(\u_div/CryTmp[9][9] ), .B(n100), .Y(\u_div/CryTmp[9][10] )
         );
  AND2X2 U392 ( .A(\u_div/CryTmp[10][15] ), .B(n159), .Y(
        \u_div/CryTmp[10][16] ) );
  AND2X2 U393 ( .A(\u_div/CryTmp[4][9] ), .B(n102), .Y(\u_div/CryTmp[4][10] )
         );
  AND2X2 U394 ( .A(\u_div/CryTmp[3][9] ), .B(n101), .Y(\u_div/CryTmp[3][10] )
         );
  AND2X2 U395 ( .A(\u_div/CryTmp[2][9] ), .B(n98), .Y(\u_div/CryTmp[2][10] )
         );
  OR2X2 U396 ( .A(\u_div/CryTmp[10][11] ), .B(n41), .Y(\u_div/CryTmp[10][12] )
         );
  OR2X2 U397 ( .A(\u_div/CryTmp[10][12] ), .B(n130), .Y(\u_div/CryTmp[10][13] ) );
  OR2X2 U398 ( .A(\u_div/CryTmp[10][13] ), .B(n53), .Y(\u_div/CryTmp[10][14] )
         );
  OR2X2 U399 ( .A(\u_div/CryTmp[9][8] ), .B(n25), .Y(\u_div/CryTmp[9][9] ) );
  OR2X2 U400 ( .A(\u_div/CryTmp[10][14] ), .B(n145), .Y(\u_div/CryTmp[10][15] ) );
  OR2X2 U401 ( .A(\u_div/CryTmp[8][8] ), .B(n26), .Y(\u_div/CryTmp[8][9] ) );
  OR2X2 U402 ( .A(\u_div/CryTmp[7][8] ), .B(n29), .Y(\u_div/CryTmp[7][9] ) );
  OR2X2 U403 ( .A(\u_div/CryTmp[6][8] ), .B(n27), .Y(\u_div/CryTmp[6][9] ) );
  OR2X2 U404 ( .A(\u_div/CryTmp[5][8] ), .B(n28), .Y(\u_div/CryTmp[5][9] ) );
  OR2X2 U405 ( .A(\u_div/CryTmp[1][8] ), .B(\u_div/PartRem[2][8] ), .Y(
        \u_div/CryTmp[1][9] ) );
  MXI2X1 U406 ( .A(n231), .B(n175), .S0(n264), .Y(\u_div/PartRem[1][10] ) );
  MXI2X1 U407 ( .A(n98), .B(\u_div/SumTmp[2][9] ), .S0(n265), .Y(n242) );
  XOR2X1 U408 ( .A(n98), .B(\u_div/CryTmp[2][9] ), .Y(\u_div/SumTmp[2][9] ) );
  XOR2X1 U409 ( .A(n99), .B(\u_div/CryTmp[10][9] ), .Y(\u_div/SumTmp[10][9] )
         );
  XOR2X1 U410 ( .A(n116), .B(\u_div/CryTmp[10][10] ), .Y(
        \u_div/SumTmp[10][10] ) );
  XNOR2X1 U411 ( .A(n25), .B(\u_div/CryTmp[9][8] ), .Y(\u_div/SumTmp[9][8] )
         );
  XOR2X1 U412 ( .A(n100), .B(\u_div/CryTmp[9][9] ), .Y(\u_div/SumTmp[9][9] )
         );
  XNOR2X1 U413 ( .A(n26), .B(\u_div/CryTmp[8][8] ), .Y(\u_div/SumTmp[8][8] )
         );
  XNOR2X1 U414 ( .A(n27), .B(\u_div/CryTmp[6][8] ), .Y(\u_div/SumTmp[6][8] )
         );
  XNOR2X1 U415 ( .A(n28), .B(\u_div/CryTmp[5][8] ), .Y(\u_div/SumTmp[5][8] )
         );
  XOR2X1 U416 ( .A(n101), .B(\u_div/CryTmp[3][9] ), .Y(\u_div/SumTmp[3][9] )
         );
  XOR2X1 U417 ( .A(n102), .B(\u_div/CryTmp[4][9] ), .Y(\u_div/SumTmp[4][9] )
         );
  XNOR2X1 U418 ( .A(n29), .B(\u_div/CryTmp[7][8] ), .Y(\u_div/SumTmp[7][8] )
         );
  INVX1 U419 ( .A(n231), .Y(\u_div/PartRem[2][9] ) );
  XNOR2X1 U420 ( .A(n41), .B(\u_div/CryTmp[10][11] ), .Y(
        \u_div/SumTmp[10][11] ) );
  XNOR2X1 U421 ( .A(n130), .B(\u_div/CryTmp[10][12] ), .Y(
        \u_div/SumTmp[10][12] ) );
  MXI2X1 U422 ( .A(n159), .B(\u_div/SumTmp[10][15] ), .S0(n276), .Y(n223) );
  XOR2X1 U423 ( .A(n159), .B(\u_div/CryTmp[10][15] ), .Y(
        \u_div/SumTmp[10][15] ) );
  XNOR2X1 U424 ( .A(n145), .B(\u_div/CryTmp[10][14] ), .Y(
        \u_div/SumTmp[10][14] ) );
  XNOR2X1 U425 ( .A(n53), .B(\u_div/CryTmp[10][13] ), .Y(
        \u_div/SumTmp[10][13] ) );
  INVX1 U426 ( .A(n255), .Y(\u_div/PartRem[11][16] ) );
  XNOR2X1 U427 ( .A(\u_div/PartRem[12][16] ), .B(\u_div/CryTmp[11][16] ), .Y(
        n201) );
  MX2X1 U428 ( .A(n254), .B(n201), .S0(n275), .Y(n202) );
  AND2X2 U429 ( .A(\u_div/CryTmp[11][10] ), .B(n117), .Y(
        \u_div/CryTmp[11][11] ) );
  AND2X2 U430 ( .A(\u_div/CryTmp[10][7] ), .B(n81), .Y(\u_div/CryTmp[10][8] )
         );
  AND2X2 U431 ( .A(\u_div/CryTmp[9][7] ), .B(n82), .Y(\u_div/CryTmp[9][8] ) );
  AND2X2 U432 ( .A(\u_div/CryTmp[8][7] ), .B(n83), .Y(\u_div/CryTmp[8][8] ) );
  AND2X2 U433 ( .A(\u_div/CryTmp[7][7] ), .B(n84), .Y(\u_div/CryTmp[7][8] ) );
  AND2X2 U434 ( .A(\u_div/CryTmp[6][7] ), .B(n85), .Y(\u_div/CryTmp[6][8] ) );
  AND2X2 U435 ( .A(\u_div/CryTmp[5][7] ), .B(n86), .Y(\u_div/CryTmp[5][8] ) );
  AND2X2 U436 ( .A(\u_div/CryTmp[11][9] ), .B(n103), .Y(\u_div/CryTmp[11][10] ) );
  AND2X2 U437 ( .A(\u_div/CryTmp[11][15] ), .B(n160), .Y(
        \u_div/CryTmp[11][16] ) );
  OR2X2 U438 ( .A(\u_div/CryTmp[11][11] ), .B(n42), .Y(\u_div/CryTmp[11][12] )
         );
  OR2X2 U439 ( .A(\u_div/CryTmp[11][12] ), .B(n131), .Y(\u_div/CryTmp[11][13] ) );
  OR2X2 U440 ( .A(\u_div/CryTmp[11][13] ), .B(n54), .Y(\u_div/CryTmp[11][14] )
         );
  OR2X2 U441 ( .A(\u_div/CryTmp[9][6] ), .B(n74), .Y(\u_div/CryTmp[9][7] ) );
  OR2X2 U442 ( .A(\u_div/CryTmp[11][8] ), .B(n30), .Y(\u_div/CryTmp[11][9] )
         );
  OR2X2 U443 ( .A(\u_div/CryTmp[10][8] ), .B(n20), .Y(\u_div/CryTmp[10][9] )
         );
  OR2X2 U444 ( .A(\u_div/CryTmp[11][14] ), .B(n146), .Y(\u_div/CryTmp[11][15] ) );
  OR2X2 U445 ( .A(\u_div/CryTmp[4][8] ), .B(n31), .Y(\u_div/CryTmp[4][9] ) );
  OR2X2 U446 ( .A(\u_div/CryTmp[3][8] ), .B(n21), .Y(\u_div/CryTmp[3][9] ) );
  OR2X2 U447 ( .A(\u_div/CryTmp[2][8] ), .B(n19), .Y(\u_div/CryTmp[2][9] ) );
  OR2X2 U448 ( .A(\u_div/CryTmp[1][6] ), .B(\u_div/PartRem[2][6] ), .Y(
        \u_div/CryTmp[1][7] ) );
  MXI2X1 U449 ( .A(n232), .B(n169), .S0(n264), .Y(\u_div/PartRem[1][9] ) );
  NAND2BX1 U450 ( .AN(n80), .B(n24), .Y(\u_div/CryTmp[0][9] ) );
  XOR2X1 U451 ( .A(n81), .B(\u_div/CryTmp[10][7] ), .Y(\u_div/SumTmp[10][7] )
         );
  XNOR2X1 U452 ( .A(n74), .B(\u_div/CryTmp[9][6] ), .Y(\u_div/SumTmp[9][6] )
         );
  XOR2X1 U453 ( .A(n82), .B(\u_div/CryTmp[9][7] ), .Y(\u_div/SumTmp[9][7] ) );
  XOR2X1 U454 ( .A(n83), .B(\u_div/CryTmp[8][7] ), .Y(\u_div/SumTmp[8][7] ) );
  XOR2X1 U455 ( .A(n84), .B(\u_div/CryTmp[7][7] ), .Y(\u_div/SumTmp[7][7] ) );
  XOR2X1 U456 ( .A(n85), .B(\u_div/CryTmp[6][7] ), .Y(\u_div/SumTmp[6][7] ) );
  XOR2X1 U457 ( .A(n86), .B(\u_div/CryTmp[5][7] ), .Y(\u_div/SumTmp[5][7] ) );
  INVX1 U458 ( .A(n234), .Y(\u_div/PartRem[2][6] ) );
  INVX1 U459 ( .A(n233), .Y(\u_div/PartRem[2][7] ) );
  INVX1 U460 ( .A(n232), .Y(\u_div/PartRem[2][8] ) );
  MXI2X1 U461 ( .A(n19), .B(\u_div/SumTmp[2][8] ), .S0(n265), .Y(n231) );
  XNOR2X1 U462 ( .A(n19), .B(\u_div/CryTmp[2][8] ), .Y(\u_div/SumTmp[2][8] )
         );
  XNOR2X1 U463 ( .A(n30), .B(\u_div/CryTmp[11][8] ), .Y(\u_div/SumTmp[11][8] )
         );
  XOR2X1 U464 ( .A(n103), .B(\u_div/CryTmp[11][9] ), .Y(\u_div/SumTmp[11][9] )
         );
  XNOR2X1 U465 ( .A(n20), .B(\u_div/CryTmp[10][8] ), .Y(\u_div/SumTmp[10][8] )
         );
  XOR2X1 U466 ( .A(n117), .B(\u_div/CryTmp[11][10] ), .Y(
        \u_div/SumTmp[11][10] ) );
  XNOR2X1 U467 ( .A(n21), .B(\u_div/CryTmp[3][8] ), .Y(\u_div/SumTmp[3][8] )
         );
  XNOR2X1 U468 ( .A(n31), .B(\u_div/CryTmp[4][8] ), .Y(\u_div/SumTmp[4][8] )
         );
  XNOR2X1 U469 ( .A(n42), .B(\u_div/CryTmp[11][11] ), .Y(
        \u_div/SumTmp[11][11] ) );
  XNOR2X1 U470 ( .A(n131), .B(\u_div/CryTmp[11][12] ), .Y(
        \u_div/SumTmp[11][12] ) );
  MXI2X1 U471 ( .A(n160), .B(\u_div/SumTmp[11][15] ), .S0(n275), .Y(n255) );
  XOR2X1 U472 ( .A(n160), .B(\u_div/CryTmp[11][15] ), .Y(
        \u_div/SumTmp[11][15] ) );
  XNOR2X1 U473 ( .A(n146), .B(\u_div/CryTmp[11][14] ), .Y(
        \u_div/SumTmp[11][14] ) );
  XNOR2X1 U474 ( .A(n54), .B(\u_div/CryTmp[11][13] ), .Y(
        \u_div/SumTmp[11][13] ) );
  INVX1 U475 ( .A(n254), .Y(\u_div/PartRem[12][16] ) );
  XOR2X1 U476 ( .A(\u_div/PartRem[2][6] ), .B(\u_div/CryTmp[1][6] ), .Y(n203)
         );
  XNOR2X1 U477 ( .A(\u_div/PartRem[13][16] ), .B(\u_div/CryTmp[12][16] ), .Y(
        n204) );
  XNOR2X1 U478 ( .A(\u_div/PartRem[15][16] ), .B(\u_div/CryTmp[14][16] ), .Y(
        n205) );
  MX2X1 U479 ( .A(n253), .B(n204), .S0(n274), .Y(n206) );
  INVX1 U480 ( .A(n260), .Y(\u_div/CryTmp[9][6] ) );
  MXI2X1 U481 ( .A(n2), .B(n2), .S0(n276), .Y(n260) );
  INVX1 U482 ( .A(n235), .Y(\u_div/CryTmp[1][6] ) );
  AND2X2 U483 ( .A(\u_div/CryTmp[12][7] ), .B(n88), .Y(\u_div/CryTmp[12][8] )
         );
  AND2X2 U484 ( .A(\u_div/CryTmp[12][10] ), .B(n118), .Y(
        \u_div/CryTmp[12][11] ) );
  AND2X2 U485 ( .A(\u_div/CryTmp[11][7] ), .B(n89), .Y(\u_div/CryTmp[11][8] )
         );
  AND2X2 U486 ( .A(\u_div/CryTmp[4][7] ), .B(n91), .Y(\u_div/CryTmp[4][8] ) );
  AND2X2 U487 ( .A(\u_div/CryTmp[3][7] ), .B(n90), .Y(\u_div/CryTmp[3][8] ) );
  AND2X2 U488 ( .A(\u_div/CryTmp[2][7] ), .B(n87), .Y(\u_div/CryTmp[2][8] ) );
  AND2X2 U489 ( .A(\u_div/CryTmp[12][9] ), .B(n104), .Y(\u_div/CryTmp[12][10] ) );
  AND2X2 U490 ( .A(\u_div/CryTmp[12][15] ), .B(n161), .Y(
        \u_div/CryTmp[12][16] ) );
  OR2X2 U491 ( .A(\u_div/CryTmp[12][11] ), .B(n43), .Y(\u_div/CryTmp[12][12] )
         );
  OR2X2 U492 ( .A(\u_div/CryTmp[12][12] ), .B(n132), .Y(\u_div/CryTmp[12][13] ) );
  OR2X2 U493 ( .A(\u_div/CryTmp[12][13] ), .B(n55), .Y(\u_div/CryTmp[12][14] )
         );
  OR2X2 U494 ( .A(\u_div/CryTmp[11][6] ), .B(n76), .Y(\u_div/CryTmp[11][7] )
         );
  OR2X2 U495 ( .A(\u_div/CryTmp[10][6] ), .B(n8), .Y(\u_div/CryTmp[10][7] ) );
  OR2X2 U496 ( .A(\u_div/CryTmp[8][6] ), .B(n9), .Y(\u_div/CryTmp[8][7] ) );
  OR2X2 U497 ( .A(\u_div/CryTmp[7][6] ), .B(n12), .Y(\u_div/CryTmp[7][7] ) );
  OR2X2 U498 ( .A(\u_div/CryTmp[6][6] ), .B(n10), .Y(\u_div/CryTmp[6][7] ) );
  OR2X2 U499 ( .A(\u_div/CryTmp[5][6] ), .B(n11), .Y(\u_div/CryTmp[5][7] ) );
  OR2X2 U500 ( .A(\u_div/CryTmp[2][6] ), .B(n75), .Y(\u_div/CryTmp[2][7] ) );
  OR2X2 U501 ( .A(\u_div/CryTmp[12][8] ), .B(n22), .Y(\u_div/CryTmp[12][9] )
         );
  OR2X2 U502 ( .A(\u_div/CryTmp[12][14] ), .B(n147), .Y(\u_div/CryTmp[12][15] ) );
  MXI2X1 U503 ( .A(n234), .B(n203), .S0(n264), .Y(\u_div/PartRem[1][7] ) );
  NAND2BX1 U504 ( .AN(\u_div/CryTmp[0][6] ), .B(n16), .Y(\u_div/CryTmp[0][7] )
         );
  MXI2X1 U505 ( .A(\u_div/CryTmp[2][6] ), .B(n245), .S0(n265), .Y(n234) );
  MXI2X1 U506 ( .A(n75), .B(\u_div/SumTmp[2][6] ), .S0(n265), .Y(n233) );
  XNOR2X1 U507 ( .A(n75), .B(\u_div/CryTmp[2][6] ), .Y(\u_div/SumTmp[2][6] )
         );
  MXI2X1 U508 ( .A(n87), .B(\u_div/SumTmp[2][7] ), .S0(n265), .Y(n232) );
  XOR2X1 U509 ( .A(n87), .B(\u_div/CryTmp[2][7] ), .Y(\u_div/SumTmp[2][7] ) );
  XNOR2X1 U510 ( .A(n76), .B(\u_div/CryTmp[11][6] ), .Y(\u_div/SumTmp[11][6] )
         );
  XNOR2X1 U511 ( .A(n8), .B(\u_div/CryTmp[10][6] ), .Y(\u_div/SumTmp[10][6] )
         );
  XOR2X1 U512 ( .A(n88), .B(\u_div/CryTmp[12][7] ), .Y(\u_div/SumTmp[12][7] )
         );
  XOR2X1 U513 ( .A(n89), .B(\u_div/CryTmp[11][7] ), .Y(\u_div/SumTmp[11][7] )
         );
  XNOR2X1 U514 ( .A(n9), .B(\u_div/CryTmp[8][6] ), .Y(\u_div/SumTmp[8][6] ) );
  XNOR2X1 U515 ( .A(n10), .B(\u_div/CryTmp[6][6] ), .Y(\u_div/SumTmp[6][6] )
         );
  XNOR2X1 U516 ( .A(n11), .B(\u_div/CryTmp[5][6] ), .Y(\u_div/SumTmp[5][6] )
         );
  XOR2X1 U517 ( .A(n90), .B(\u_div/CryTmp[3][7] ), .Y(\u_div/SumTmp[3][7] ) );
  XOR2X1 U518 ( .A(n91), .B(\u_div/CryTmp[4][7] ), .Y(\u_div/SumTmp[4][7] ) );
  XNOR2X1 U519 ( .A(n12), .B(\u_div/CryTmp[7][6] ), .Y(\u_div/SumTmp[7][6] )
         );
  AND2X2 U520 ( .A(\u_div/CryTmp[14][15] ), .B(n163), .Y(
        \u_div/CryTmp[14][16] ) );
  OR2X2 U521 ( .A(\u_div/CryTmp[14][13] ), .B(n135), .Y(\u_div/CryTmp[14][14] ) );
  OR2X2 U522 ( .A(\u_div/CryTmp[14][14] ), .B(n149), .Y(\u_div/CryTmp[14][15] ) );
  XNOR2X1 U523 ( .A(n22), .B(\u_div/CryTmp[12][8] ), .Y(\u_div/SumTmp[12][8] )
         );
  XOR2X1 U524 ( .A(n104), .B(\u_div/CryTmp[12][9] ), .Y(\u_div/SumTmp[12][9] )
         );
  XOR2X1 U525 ( .A(n118), .B(\u_div/CryTmp[12][10] ), .Y(
        \u_div/SumTmp[12][10] ) );
  XNOR2X1 U526 ( .A(n43), .B(\u_div/CryTmp[12][11] ), .Y(
        \u_div/SumTmp[12][11] ) );
  XNOR2X1 U527 ( .A(n132), .B(\u_div/CryTmp[12][12] ), .Y(
        \u_div/SumTmp[12][12] ) );
  MXI2X1 U528 ( .A(n161), .B(\u_div/SumTmp[12][15] ), .S0(n274), .Y(n254) );
  XOR2X1 U529 ( .A(n161), .B(\u_div/CryTmp[12][15] ), .Y(
        \u_div/SumTmp[12][15] ) );
  XNOR2X1 U530 ( .A(n147), .B(\u_div/CryTmp[12][14] ), .Y(
        \u_div/SumTmp[12][14] ) );
  XNOR2X1 U531 ( .A(n55), .B(\u_div/CryTmp[12][13] ), .Y(
        \u_div/SumTmp[12][13] ) );
  INVX1 U532 ( .A(n253), .Y(\u_div/PartRem[13][16] ) );
  INVX1 U533 ( .A(n251), .Y(\u_div/PartRem[15][16] ) );
  XNOR2X1 U534 ( .A(\u_div/PartRem[14][16] ), .B(\u_div/CryTmp[13][16] ), .Y(
        n207) );
  MX2X1 U535 ( .A(n252), .B(n207), .S0(n273), .Y(n208) );
  INVX1 U536 ( .A(n258), .Y(\u_div/CryTmp[11][6] ) );
  MXI2X1 U537 ( .A(n58), .B(n58), .S0(n274), .Y(n258) );
  INVX1 U538 ( .A(n259), .Y(\u_div/CryTmp[10][6] ) );
  MXI2X1 U539 ( .A(n165), .B(n165), .S0(n275), .Y(n259) );
  INVX1 U540 ( .A(n246), .Y(\u_div/CryTmp[8][6] ) );
  MXI2X1 U541 ( .A(n3), .B(n3), .S0(n271), .Y(n246) );
  INVX1 U542 ( .A(n247), .Y(\u_div/CryTmp[7][6] ) );
  MXI2X1 U543 ( .A(n4), .B(n4), .S0(n267), .Y(n247) );
  INVX1 U544 ( .A(n249), .Y(\u_div/CryTmp[5][6] ) );
  MXI2X1 U545 ( .A(n5), .B(n5), .S0(n263), .Y(n249) );
  INVX1 U546 ( .A(n245), .Y(\u_div/CryTmp[2][6] ) );
  MXI2X1 U547 ( .A(n171), .B(n171), .S0(n268), .Y(n245) );
  MXI2X1 U548 ( .A(n60), .B(n60), .S0(n265), .Y(n235) );
  INVX1 U549 ( .A(n248), .Y(\u_div/CryTmp[6][6] ) );
  MXI2X1 U550 ( .A(n6), .B(n6), .S0(n266), .Y(n248) );
  MX2X1 U551 ( .A(n209), .B(n209), .S0(n264), .Y(\u_div/CryTmp[0][6] ) );
  MX2X1 U552 ( .A(n71), .B(n71), .S0(n265), .Y(n209) );
  AND2X2 U553 ( .A(\u_div/CryTmp[13][7] ), .B(n92), .Y(\u_div/CryTmp[13][8] )
         );
  AND2X2 U554 ( .A(\u_div/CryTmp[13][10] ), .B(n119), .Y(
        \u_div/CryTmp[13][11] ) );
  AND2X2 U555 ( .A(\u_div/CryTmp[13][9] ), .B(n105), .Y(\u_div/CryTmp[13][10] ) );
  AND2X2 U556 ( .A(\u_div/CryTmp[13][15] ), .B(n162), .Y(
        \u_div/CryTmp[13][16] ) );
  OR2X2 U557 ( .A(\u_div/CryTmp[13][11] ), .B(n44), .Y(\u_div/CryTmp[13][12] )
         );
  OR2X2 U558 ( .A(\u_div/CryTmp[13][12] ), .B(n133), .Y(\u_div/CryTmp[13][13] ) );
  OR2X2 U559 ( .A(\u_div/CryTmp[13][13] ), .B(n56), .Y(\u_div/CryTmp[13][14] )
         );
  OR2X2 U560 ( .A(\u_div/CryTmp[13][6] ), .B(n77), .Y(\u_div/CryTmp[13][7] )
         );
  OR2X2 U561 ( .A(\u_div/CryTmp[12][6] ), .B(n13), .Y(\u_div/CryTmp[12][7] )
         );
  OR2X2 U562 ( .A(\u_div/CryTmp[4][6] ), .B(n15), .Y(\u_div/CryTmp[4][7] ) );
  OR2X2 U563 ( .A(\u_div/CryTmp[3][6] ), .B(n14), .Y(\u_div/CryTmp[3][7] ) );
  OR2X2 U564 ( .A(\u_div/CryTmp[13][8] ), .B(n32), .Y(\u_div/CryTmp[13][9] )
         );
  OR2X2 U565 ( .A(\u_div/CryTmp[13][14] ), .B(n148), .Y(\u_div/CryTmp[13][15] ) );
  XNOR2X1 U566 ( .A(n77), .B(\u_div/CryTmp[13][6] ), .Y(\u_div/SumTmp[13][6] )
         );
  XNOR2X1 U567 ( .A(n13), .B(\u_div/CryTmp[12][6] ), .Y(\u_div/SumTmp[12][6] )
         );
  XOR2X1 U568 ( .A(n92), .B(\u_div/CryTmp[13][7] ), .Y(\u_div/SumTmp[13][7] )
         );
  XNOR2X1 U569 ( .A(n14), .B(\u_div/CryTmp[3][6] ), .Y(\u_div/SumTmp[3][6] )
         );
  XNOR2X1 U570 ( .A(n15), .B(\u_div/CryTmp[4][6] ), .Y(\u_div/SumTmp[4][6] )
         );
  AND2X2 U571 ( .A(\u_div/CryTmp[14][7] ), .B(n93), .Y(\u_div/CryTmp[14][8] )
         );
  AND2X2 U572 ( .A(\u_div/CryTmp[14][9] ), .B(n106), .Y(\u_div/CryTmp[14][10] ) );
  AND2X2 U573 ( .A(\u_div/CryTmp[15][15] ), .B(a[30]), .Y(
        \u_div/CryTmp[15][16] ) );
  OR2X2 U574 ( .A(\u_div/CryTmp[14][12] ), .B(n134), .Y(\u_div/CryTmp[14][13] ) );
  OR2X2 U575 ( .A(\u_div/CryTmp[14][6] ), .B(n1), .Y(\u_div/CryTmp[14][7] ) );
  OR2X2 U576 ( .A(\u_div/CryTmp[14][8] ), .B(n23), .Y(\u_div/CryTmp[14][9] )
         );
  OR2X2 U577 ( .A(\u_div/CryTmp[15][14] ), .B(a[29]), .Y(
        \u_div/CryTmp[15][15] ) );
  XNOR2X1 U578 ( .A(n32), .B(\u_div/CryTmp[13][8] ), .Y(\u_div/SumTmp[13][8] )
         );
  XOR2X1 U579 ( .A(n105), .B(\u_div/CryTmp[13][9] ), .Y(\u_div/SumTmp[13][9] )
         );
  XOR2X1 U580 ( .A(n119), .B(\u_div/CryTmp[13][10] ), .Y(
        \u_div/SumTmp[13][10] ) );
  OR2X2 U581 ( .A(\u_div/CryTmp[15][12] ), .B(a[27]), .Y(
        \u_div/CryTmp[15][13] ) );
  OR2X2 U582 ( .A(\u_div/CryTmp[15][13] ), .B(a[28]), .Y(
        \u_div/CryTmp[15][14] ) );
  XNOR2X1 U583 ( .A(n44), .B(\u_div/CryTmp[13][11] ), .Y(
        \u_div/SumTmp[13][11] ) );
  XNOR2X1 U584 ( .A(n133), .B(\u_div/CryTmp[13][12] ), .Y(
        \u_div/SumTmp[13][12] ) );
  XNOR2X1 U585 ( .A(a[27]), .B(\u_div/CryTmp[15][12] ), .Y(
        \u_div/SumTmp[15][12] ) );
  MXI2X1 U586 ( .A(n162), .B(\u_div/SumTmp[13][15] ), .S0(n273), .Y(n253) );
  XOR2X1 U587 ( .A(n162), .B(\u_div/CryTmp[13][15] ), .Y(
        \u_div/SumTmp[13][15] ) );
  MXI2X1 U588 ( .A(a[30]), .B(\u_div/SumTmp[15][15] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n251) );
  XOR2X1 U589 ( .A(a[30]), .B(\u_div/CryTmp[15][15] ), .Y(
        \u_div/SumTmp[15][15] ) );
  XNOR2X1 U590 ( .A(a[29]), .B(\u_div/CryTmp[15][14] ), .Y(
        \u_div/SumTmp[15][14] ) );
  XNOR2X1 U591 ( .A(n148), .B(\u_div/CryTmp[13][14] ), .Y(
        \u_div/SumTmp[13][14] ) );
  XNOR2X1 U592 ( .A(n56), .B(\u_div/CryTmp[13][13] ), .Y(
        \u_div/SumTmp[13][13] ) );
  XNOR2X1 U593 ( .A(a[28]), .B(\u_div/CryTmp[15][13] ), .Y(
        \u_div/SumTmp[15][13] ) );
  INVX1 U594 ( .A(n252), .Y(\u_div/PartRem[14][16] ) );
  MX2X1 U595 ( .A(n251), .B(n205), .S0(n272), .Y(n210) );
  INVX1 U596 ( .A(n256), .Y(\u_div/CryTmp[13][6] ) );
  MXI2X1 U597 ( .A(n59), .B(n59), .S0(n272), .Y(n256) );
  INVX1 U598 ( .A(n257), .Y(\u_div/CryTmp[12][6] ) );
  MXI2X1 U599 ( .A(n166), .B(n166), .S0(n273), .Y(n257) );
  INVX1 U600 ( .A(n243), .Y(\u_div/CryTmp[4][6] ) );
  MXI2X1 U601 ( .A(n7), .B(n7), .S0(n269), .Y(n243) );
  INVX1 U602 ( .A(n244), .Y(\u_div/CryTmp[3][6] ) );
  MXI2X1 U603 ( .A(n172), .B(n172), .S0(n270), .Y(n244) );
  INVX1 U604 ( .A(n262), .Y(\u_div/CryTmp[14][6] ) );
  MXI2X1 U605 ( .A(\u_div/PartRem[19][1] ), .B(\u_div/PartRem[19][1] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n262) );
  XNOR2X1 U606 ( .A(\u_div/PartRem[21][1] ), .B(\u_div/PartRem[20][1] ), .Y(
        \u_div/SumTmp[15][6] ) );
  XNOR2X1 U607 ( .A(n1), .B(\u_div/CryTmp[14][6] ), .Y(\u_div/SumTmp[14][6] )
         );
  XOR2X1 U608 ( .A(n93), .B(\u_div/CryTmp[14][7] ), .Y(\u_div/SumTmp[14][7] )
         );
  XOR2X1 U609 ( .A(\u_div/PartRem[22][1] ), .B(\u_div/CryTmp[15][7] ), .Y(
        \u_div/SumTmp[15][7] ) );
  AND2X2 U610 ( .A(\u_div/CryTmp[14][10] ), .B(n120), .Y(
        \u_div/CryTmp[14][11] ) );
  OR2X2 U611 ( .A(\u_div/CryTmp[14][11] ), .B(n107), .Y(\u_div/CryTmp[14][12] ) );
  XOR2X1 U612 ( .A(n106), .B(\u_div/CryTmp[14][9] ), .Y(\u_div/SumTmp[14][9] )
         );
  XOR2X1 U613 ( .A(n120), .B(\u_div/CryTmp[14][10] ), .Y(
        \u_div/SumTmp[14][10] ) );
  XNOR2X1 U614 ( .A(\u_div/PartRem[23][1] ), .B(\u_div/CryTmp[15][8] ), .Y(
        \u_div/SumTmp[15][8] ) );
  XNOR2X1 U615 ( .A(n23), .B(\u_div/CryTmp[14][8] ), .Y(\u_div/SumTmp[14][8] )
         );
  OR2X2 U616 ( .A(\u_div/CryTmp[15][11] ), .B(a[26]), .Y(
        \u_div/CryTmp[15][12] ) );
  XNOR2X1 U617 ( .A(n107), .B(\u_div/CryTmp[14][11] ), .Y(
        \u_div/SumTmp[14][11] ) );
  XNOR2X1 U618 ( .A(n134), .B(\u_div/CryTmp[14][12] ), .Y(
        \u_div/SumTmp[14][12] ) );
  XNOR2X1 U619 ( .A(a[26]), .B(\u_div/CryTmp[15][11] ), .Y(
        \u_div/SumTmp[15][11] ) );
  AND2X2 U620 ( .A(\u_div/CryTmp[15][7] ), .B(\u_div/PartRem[22][1] ), .Y(
        \u_div/CryTmp[15][8] ) );
  OR2X2 U621 ( .A(\u_div/PartRem[20][1] ), .B(\u_div/PartRem[21][1] ), .Y(
        \u_div/CryTmp[15][7] ) );
  OR2X2 U622 ( .A(\u_div/CryTmp[15][8] ), .B(\u_div/PartRem[23][1] ), .Y(
        \u_div/CryTmp[15][9] ) );
  MXI2X1 U623 ( .A(n163), .B(\u_div/SumTmp[14][15] ), .S0(n272), .Y(n252) );
  XOR2X1 U624 ( .A(n163), .B(\u_div/CryTmp[14][15] ), .Y(
        \u_div/SumTmp[14][15] ) );
  XNOR2X1 U625 ( .A(n149), .B(\u_div/CryTmp[14][14] ), .Y(
        \u_div/SumTmp[14][14] ) );
  XNOR2X1 U626 ( .A(n135), .B(\u_div/CryTmp[14][13] ), .Y(
        \u_div/SumTmp[14][13] ) );
  XNOR2X1 U627 ( .A(\u_div/PartRem[31][1] ), .B(\u_div/CryTmp[15][16] ), .Y(
        n211) );
  MX2X1 U628 ( .A(\u_div/SumTmp[14][0] ), .B(\u_div/SumTmp[14][0] ), .S0(n272), 
        .Y(n212) );
  MX2X1 U629 ( .A(\u_div/SumTmp[15][0] ), .B(\u_div/SumTmp[15][0] ), .S0(
        \u_div/CryTmp[15][17] ), .Y(n213) );
  MX2X1 U630 ( .A(n250), .B(n211), .S0(\u_div/CryTmp[15][17] ), .Y(n214) );
  XOR2X1 U631 ( .A(\u_div/PartRem[24][1] ), .B(\u_div/CryTmp[15][9] ), .Y(
        \u_div/SumTmp[15][9] ) );
  AND2X2 U632 ( .A(\u_div/CryTmp[15][10] ), .B(\u_div/PartRem[25][1] ), .Y(
        \u_div/CryTmp[15][11] ) );
  INVX1 U633 ( .A(\u_div/PartRem[20][1] ), .Y(n261) );
  XOR2X1 U634 ( .A(\u_div/PartRem[25][1] ), .B(\u_div/CryTmp[15][10] ), .Y(
        \u_div/SumTmp[15][10] ) );
  AND2X2 U635 ( .A(\u_div/CryTmp[15][9] ), .B(\u_div/PartRem[24][1] ), .Y(
        \u_div/CryTmp[15][10] ) );
  MX2X1 U636 ( .A(\u_div/SumTmp[10][0] ), .B(\u_div/SumTmp[10][0] ), .S0(n276), 
        .Y(n215) );
  MX2X1 U637 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[7][0] ), .S0(n266), 
        .Y(n216) );
  MX2X1 U638 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[5][0] ), .S0(n269), 
        .Y(n217) );
  MX2X1 U639 ( .A(\u_div/SumTmp[11][0] ), .B(\u_div/SumTmp[11][0] ), .S0(n275), 
        .Y(n218) );
  MX2X1 U640 ( .A(\u_div/SumTmp[12][0] ), .B(\u_div/SumTmp[12][0] ), .S0(n274), 
        .Y(n219) );
  MX2X1 U641 ( .A(\u_div/SumTmp[13][0] ), .B(\u_div/SumTmp[13][0] ), .S0(n273), 
        .Y(n220) );
  INVX1 U642 ( .A(\u_div/PartRem[31][1] ), .Y(n250) );
  MX2X1 U643 ( .A(\u_div/SumTmp[9][0] ), .B(\u_div/SumTmp[9][0] ), .S0(n271), 
        .Y(n221) );
  MX2X1 U644 ( .A(\u_div/SumTmp[8][0] ), .B(\u_div/SumTmp[8][0] ), .S0(n267), 
        .Y(n222) );
  NAND2BX4 U645 ( .AN(\u_div/CryTmp[14][17] ), .B(n214), .Y(n272) );
  NAND2BX4 U646 ( .AN(\u_div/CryTmp[13][17] ), .B(n210), .Y(n273) );
  NAND2BX4 U647 ( .AN(\u_div/CryTmp[12][17] ), .B(n208), .Y(n274) );
  NAND2BX4 U648 ( .AN(\u_div/CryTmp[11][17] ), .B(n206), .Y(n275) );
  NAND2BX4 U649 ( .AN(\u_div/CryTmp[10][17] ), .B(n202), .Y(n276) );
  AND2X4 U650 ( .A(\u_div/CryTmp[15][16] ), .B(\u_div/PartRem[31][1] ), .Y(
        \u_div/CryTmp[15][17] ) );
endmodule


module Equation_Implementation_DW_div_uns_29 ( a, b, quotient, remainder, 
        divide_by_0 );
  input [21:0] a;
  input [11:0] b;
  output [21:0] quotient;
  output [11:0] remainder;
  output divide_by_0;
  wire   \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] , \u_div/SumTmp[1][3] ,
         \u_div/SumTmp[1][4] , \u_div/SumTmp[1][5] , \u_div/SumTmp[1][6] ,
         \u_div/SumTmp[1][7] , \u_div/SumTmp[1][8] , \u_div/SumTmp[1][9] ,
         \u_div/SumTmp[1][10] , \u_div/SumTmp[1][11] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[2][5] , \u_div/SumTmp[2][6] , \u_div/SumTmp[2][7] ,
         \u_div/SumTmp[2][8] , \u_div/SumTmp[2][9] , \u_div/SumTmp[2][10] ,
         \u_div/SumTmp[2][11] , \u_div/SumTmp[3][0] , \u_div/SumTmp[3][1] ,
         \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] , \u_div/SumTmp[3][4] ,
         \u_div/SumTmp[3][5] , \u_div/SumTmp[3][6] , \u_div/SumTmp[3][7] ,
         \u_div/SumTmp[3][8] , \u_div/SumTmp[3][9] , \u_div/SumTmp[3][10] ,
         \u_div/SumTmp[3][11] , \u_div/SumTmp[4][0] , \u_div/SumTmp[4][1] ,
         \u_div/SumTmp[4][2] , \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] ,
         \u_div/SumTmp[4][5] , \u_div/SumTmp[4][6] , \u_div/SumTmp[4][7] ,
         \u_div/SumTmp[4][8] , \u_div/SumTmp[4][9] , \u_div/SumTmp[4][10] ,
         \u_div/SumTmp[4][11] , \u_div/SumTmp[5][0] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[5][5] , \u_div/SumTmp[5][6] , \u_div/SumTmp[5][7] ,
         \u_div/SumTmp[5][8] , \u_div/SumTmp[5][9] , \u_div/SumTmp[5][10] ,
         \u_div/SumTmp[5][11] , \u_div/SumTmp[6][0] , \u_div/SumTmp[6][1] ,
         \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] , \u_div/SumTmp[6][4] ,
         \u_div/SumTmp[6][5] , \u_div/SumTmp[6][6] , \u_div/SumTmp[6][7] ,
         \u_div/SumTmp[6][8] , \u_div/SumTmp[6][9] , \u_div/SumTmp[6][10] ,
         \u_div/SumTmp[6][11] , \u_div/SumTmp[7][0] , \u_div/SumTmp[7][1] ,
         \u_div/SumTmp[7][2] , \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] ,
         \u_div/SumTmp[7][5] , \u_div/SumTmp[7][6] , \u_div/SumTmp[7][7] ,
         \u_div/SumTmp[7][8] , \u_div/SumTmp[7][9] , \u_div/SumTmp[7][10] ,
         \u_div/SumTmp[7][11] , \u_div/SumTmp[8][0] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[8][5] , \u_div/SumTmp[8][6] , \u_div/SumTmp[8][7] ,
         \u_div/SumTmp[8][8] , \u_div/SumTmp[8][9] , \u_div/SumTmp[8][10] ,
         \u_div/SumTmp[8][11] , \u_div/SumTmp[9][0] , \u_div/SumTmp[9][1] ,
         \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] , \u_div/SumTmp[9][4] ,
         \u_div/SumTmp[9][5] , \u_div/SumTmp[9][6] , \u_div/SumTmp[9][7] ,
         \u_div/SumTmp[9][8] , \u_div/SumTmp[9][9] , \u_div/SumTmp[9][10] ,
         \u_div/SumTmp[9][11] , \u_div/SumTmp[10][0] , \u_div/SumTmp[10][1] ,
         \u_div/SumTmp[10][2] , \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] ,
         \u_div/SumTmp[10][5] , \u_div/SumTmp[10][6] , \u_div/SumTmp[10][7] ,
         \u_div/SumTmp[10][8] , \u_div/SumTmp[10][9] , \u_div/SumTmp[10][10] ,
         \u_div/SumTmp[10][11] , \u_div/SumTmp[11][0] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[11][5] , \u_div/SumTmp[11][6] , \u_div/SumTmp[11][7] ,
         \u_div/SumTmp[11][8] , \u_div/SumTmp[11][9] , \u_div/SumTmp[11][10] ,
         \u_div/SumTmp[12][0] , \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] ,
         \u_div/SumTmp[12][3] , \u_div/SumTmp[12][4] , \u_div/SumTmp[12][5] ,
         \u_div/SumTmp[12][6] , \u_div/SumTmp[12][7] , \u_div/SumTmp[12][8] ,
         \u_div/SumTmp[12][9] , \u_div/SumTmp[13][0] , \u_div/SumTmp[13][1] ,
         \u_div/SumTmp[13][2] , \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] ,
         \u_div/SumTmp[13][5] , \u_div/SumTmp[13][6] , \u_div/SumTmp[13][7] ,
         \u_div/SumTmp[13][8] , \u_div/SumTmp[14][0] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[14][5] , \u_div/SumTmp[14][6] , \u_div/SumTmp[14][7] ,
         \u_div/SumTmp[15][0] , \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] ,
         \u_div/SumTmp[15][3] , \u_div/SumTmp[15][4] , \u_div/SumTmp[15][5] ,
         \u_div/SumTmp[15][6] , \u_div/SumTmp[16][0] , \u_div/SumTmp[16][1] ,
         \u_div/SumTmp[16][2] , \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] ,
         \u_div/SumTmp[16][5] , \u_div/SumTmp[17][0] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[18][0] , \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] ,
         \u_div/SumTmp[18][3] , \u_div/SumTmp[19][0] , \u_div/SumTmp[19][1] ,
         \u_div/SumTmp[19][2] , \u_div/SumTmp[20][0] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[21][0] , \u_div/CryTmp[0][2] , \u_div/CryTmp[0][3] ,
         \u_div/CryTmp[0][4] , \u_div/CryTmp[0][5] , \u_div/CryTmp[0][6] ,
         \u_div/CryTmp[0][7] , \u_div/CryTmp[0][8] , \u_div/CryTmp[0][9] ,
         \u_div/CryTmp[0][10] , \u_div/CryTmp[0][11] , \u_div/CryTmp[0][12] ,
         \u_div/CryTmp[1][2] , \u_div/CryTmp[1][3] , \u_div/CryTmp[1][4] ,
         \u_div/CryTmp[1][5] , \u_div/CryTmp[1][6] , \u_div/CryTmp[1][7] ,
         \u_div/CryTmp[1][8] , \u_div/CryTmp[1][9] , \u_div/CryTmp[1][10] ,
         \u_div/CryTmp[1][11] , \u_div/CryTmp[1][12] , \u_div/CryTmp[2][1] ,
         \u_div/CryTmp[2][2] , \u_div/CryTmp[2][3] , \u_div/CryTmp[2][4] ,
         \u_div/CryTmp[2][5] , \u_div/CryTmp[2][6] , \u_div/CryTmp[2][7] ,
         \u_div/CryTmp[2][8] , \u_div/CryTmp[2][9] , \u_div/CryTmp[2][10] ,
         \u_div/CryTmp[2][11] , \u_div/CryTmp[2][12] , \u_div/CryTmp[3][1] ,
         \u_div/CryTmp[3][2] , \u_div/CryTmp[3][3] , \u_div/CryTmp[3][4] ,
         \u_div/CryTmp[3][5] , \u_div/CryTmp[3][6] , \u_div/CryTmp[3][7] ,
         \u_div/CryTmp[3][8] , \u_div/CryTmp[3][9] , \u_div/CryTmp[3][10] ,
         \u_div/CryTmp[3][11] , \u_div/CryTmp[3][12] , \u_div/CryTmp[4][1] ,
         \u_div/CryTmp[4][2] , \u_div/CryTmp[4][3] , \u_div/CryTmp[4][4] ,
         \u_div/CryTmp[4][5] , \u_div/CryTmp[4][6] , \u_div/CryTmp[4][7] ,
         \u_div/CryTmp[4][8] , \u_div/CryTmp[4][9] , \u_div/CryTmp[4][10] ,
         \u_div/CryTmp[4][11] , \u_div/CryTmp[4][12] , \u_div/CryTmp[5][1] ,
         \u_div/CryTmp[5][2] , \u_div/CryTmp[5][3] , \u_div/CryTmp[5][4] ,
         \u_div/CryTmp[5][5] , \u_div/CryTmp[5][6] , \u_div/CryTmp[5][7] ,
         \u_div/CryTmp[5][8] , \u_div/CryTmp[5][9] , \u_div/CryTmp[5][10] ,
         \u_div/CryTmp[5][11] , \u_div/CryTmp[5][12] , \u_div/CryTmp[6][1] ,
         \u_div/CryTmp[6][2] , \u_div/CryTmp[6][3] , \u_div/CryTmp[6][4] ,
         \u_div/CryTmp[6][5] , \u_div/CryTmp[6][6] , \u_div/CryTmp[6][7] ,
         \u_div/CryTmp[6][8] , \u_div/CryTmp[6][9] , \u_div/CryTmp[6][10] ,
         \u_div/CryTmp[6][11] , \u_div/CryTmp[6][12] , \u_div/CryTmp[7][1] ,
         \u_div/CryTmp[7][2] , \u_div/CryTmp[7][3] , \u_div/CryTmp[7][4] ,
         \u_div/CryTmp[7][5] , \u_div/CryTmp[7][6] , \u_div/CryTmp[7][7] ,
         \u_div/CryTmp[7][8] , \u_div/CryTmp[7][9] , \u_div/CryTmp[7][10] ,
         \u_div/CryTmp[7][11] , \u_div/CryTmp[7][12] , \u_div/CryTmp[8][1] ,
         \u_div/CryTmp[8][2] , \u_div/CryTmp[8][3] , \u_div/CryTmp[8][4] ,
         \u_div/CryTmp[8][5] , \u_div/CryTmp[8][6] , \u_div/CryTmp[8][7] ,
         \u_div/CryTmp[8][8] , \u_div/CryTmp[8][9] , \u_div/CryTmp[8][10] ,
         \u_div/CryTmp[8][11] , \u_div/CryTmp[8][12] , \u_div/CryTmp[9][1] ,
         \u_div/CryTmp[9][2] , \u_div/CryTmp[9][3] , \u_div/CryTmp[9][4] ,
         \u_div/CryTmp[9][5] , \u_div/CryTmp[9][6] , \u_div/CryTmp[9][7] ,
         \u_div/CryTmp[9][8] , \u_div/CryTmp[9][9] , \u_div/CryTmp[9][10] ,
         \u_div/CryTmp[9][11] , \u_div/CryTmp[9][12] , \u_div/CryTmp[10][1] ,
         \u_div/CryTmp[10][2] , \u_div/CryTmp[10][3] , \u_div/CryTmp[10][4] ,
         \u_div/CryTmp[10][5] , \u_div/CryTmp[10][6] , \u_div/CryTmp[10][7] ,
         \u_div/CryTmp[10][8] , \u_div/CryTmp[10][9] , \u_div/CryTmp[10][10] ,
         \u_div/CryTmp[10][11] , \u_div/CryTmp[10][12] , \u_div/CryTmp[11][1] ,
         \u_div/CryTmp[11][2] , \u_div/CryTmp[11][3] , \u_div/CryTmp[11][4] ,
         \u_div/CryTmp[11][5] , \u_div/CryTmp[11][6] , \u_div/CryTmp[11][7] ,
         \u_div/CryTmp[11][8] , \u_div/CryTmp[11][9] , \u_div/CryTmp[11][10] ,
         \u_div/CryTmp[11][11] , \u_div/CryTmp[12][1] , \u_div/CryTmp[12][2] ,
         \u_div/CryTmp[12][3] , \u_div/CryTmp[12][4] , \u_div/CryTmp[12][5] ,
         \u_div/CryTmp[12][6] , \u_div/CryTmp[12][7] , \u_div/CryTmp[12][8] ,
         \u_div/CryTmp[12][9] , \u_div/CryTmp[12][10] , \u_div/CryTmp[13][1] ,
         \u_div/CryTmp[13][2] , \u_div/CryTmp[13][3] , \u_div/CryTmp[13][4] ,
         \u_div/CryTmp[13][5] , \u_div/CryTmp[13][6] , \u_div/CryTmp[13][7] ,
         \u_div/CryTmp[13][8] , \u_div/CryTmp[13][9] , \u_div/CryTmp[14][1] ,
         \u_div/CryTmp[14][2] , \u_div/CryTmp[14][3] , \u_div/CryTmp[14][4] ,
         \u_div/CryTmp[14][5] , \u_div/CryTmp[14][6] , \u_div/CryTmp[14][7] ,
         \u_div/CryTmp[14][8] , \u_div/CryTmp[15][1] , \u_div/CryTmp[15][2] ,
         \u_div/CryTmp[15][3] , \u_div/CryTmp[15][4] , \u_div/CryTmp[15][5] ,
         \u_div/CryTmp[15][6] , \u_div/CryTmp[15][7] , \u_div/CryTmp[16][1] ,
         \u_div/CryTmp[16][2] , \u_div/CryTmp[16][3] , \u_div/CryTmp[16][4] ,
         \u_div/CryTmp[16][5] , \u_div/CryTmp[16][6] , \u_div/CryTmp[17][1] ,
         \u_div/CryTmp[17][2] , \u_div/CryTmp[17][3] , \u_div/CryTmp[17][4] ,
         \u_div/CryTmp[17][5] , \u_div/CryTmp[18][1] , \u_div/CryTmp[18][2] ,
         \u_div/CryTmp[18][3] , \u_div/CryTmp[18][4] , \u_div/CryTmp[19][1] ,
         \u_div/CryTmp[19][2] , \u_div/CryTmp[19][3] , \u_div/CryTmp[20][1] ,
         \u_div/CryTmp[20][2] , \u_div/CryTmp[21][1] , \u_div/PartRem[1][2] ,
         \u_div/PartRem[1][3] , \u_div/PartRem[1][4] , \u_div/PartRem[1][5] ,
         \u_div/PartRem[1][6] , \u_div/PartRem[1][7] , \u_div/PartRem[1][8] ,
         \u_div/PartRem[1][9] , \u_div/PartRem[1][10] , \u_div/PartRem[1][11] ,
         \u_div/PartRem[2][1] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[2][4] , \u_div/PartRem[2][5] , \u_div/PartRem[2][6] ,
         \u_div/PartRem[2][7] , \u_div/PartRem[2][8] , \u_div/PartRem[2][9] ,
         \u_div/PartRem[2][10] , \u_div/PartRem[2][11] ,
         \u_div/PartRem[3][11] , \u_div/PartRem[4][11] ,
         \u_div/PartRem[5][11] , \u_div/PartRem[6][11] ,
         \u_div/PartRem[7][11] , \u_div/PartRem[8][11] ,
         \u_div/PartRem[9][11] , \u_div/PartRem[10][11] ,
         \u_div/PartRem[11][11] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227;
  wire   [11:0] \u_div/BInv ;

  ADDFX2 \u_div/u_fa_PartRem_0_3_1  ( .A(n2), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[3][2] ), .S(
        \u_div/SumTmp[3][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_1  ( .A(n11), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[4][1] ), .CO(\u_div/CryTmp[4][2] ), .S(
        \u_div/SumTmp[4][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_2  ( .A(n157), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[3][2] ), .CO(\u_div/CryTmp[3][3] ), .S(
        \u_div/SumTmp[3][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_2  ( .A(n148), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[4][2] ), .CO(\u_div/CryTmp[4][3] ), .S(
        \u_div/SumTmp[4][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_1  ( .A(n10), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[5][1] ), .CO(\u_div/CryTmp[5][2] ), .S(
        \u_div/SumTmp[5][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_1  ( .A(n9), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[6][1] ), .CO(\u_div/CryTmp[6][2] ), .S(
        \u_div/SumTmp[6][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_1  ( .A(n8), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[7][1] ), .CO(\u_div/CryTmp[7][2] ), .S(
        \u_div/SumTmp[7][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_1  ( .A(n7), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[8][1] ), .CO(\u_div/CryTmp[8][2] ), .S(
        \u_div/SumTmp[8][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_1  ( .A(n15), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[9][1] ), .CO(\u_div/CryTmp[9][2] ), .S(
        \u_div/SumTmp[9][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_1  ( .A(n6), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[10][1] ), .CO(\u_div/CryTmp[10][2] ), .S(
        \u_div/SumTmp[10][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_1  ( .A(n13), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[18][1] ), .CO(\u_div/CryTmp[18][2] ), .S(
        \u_div/SumTmp[18][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_1  ( .A(n18), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[19][1] ), .CO(\u_div/CryTmp[19][2] ), .S(
        \u_div/SumTmp[19][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_1  ( .A(n17), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[20][1] ), .CO(\u_div/CryTmp[20][2] ), .S(
        \u_div/SumTmp[20][1] ) );
  CMPR32X1 \u_div/u_fa_PartRem_0_2_1  ( .A(n1), .B(\u_div/BInv [1]), .C(
        \u_div/CryTmp[2][1] ), .CO(\u_div/CryTmp[2][2] ), .S(
        \u_div/SumTmp[2][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_3  ( .A(n155), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[3][3] ), .CO(\u_div/CryTmp[3][4] ), .S(
        \u_div/SumTmp[3][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_3  ( .A(n128), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[4][3] ), .CO(\u_div/CryTmp[4][4] ), .S(
        \u_div/SumTmp[4][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/BInv [2]), .CI(\u_div/CryTmp[1][2] ), .CO(\u_div/CryTmp[1][3] ), 
        .S(\u_div/SumTmp[1][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_2  ( .A(n158), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[2][2] ), .CO(\u_div/CryTmp[2][3] ), .S(
        \u_div/SumTmp[2][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_2  ( .A(n147), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[5][2] ), .CO(\u_div/CryTmp[5][3] ), .S(
        \u_div/SumTmp[5][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_2  ( .A(n146), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[6][2] ), .CO(\u_div/CryTmp[6][3] ), .S(
        \u_div/SumTmp[6][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_2  ( .A(n145), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[7][2] ), .CO(\u_div/CryTmp[7][3] ), .S(
        \u_div/SumTmp[7][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_2  ( .A(n144), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[8][2] ), .CO(\u_div/CryTmp[8][3] ), .S(
        \u_div/SumTmp[8][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_2  ( .A(n118), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[10][2] ), .CO(\u_div/CryTmp[10][3] ), .S(
        \u_div/SumTmp[10][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_2  ( .A(n149), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[9][2] ), .CO(\u_div/CryTmp[9][3] ), .S(
        \u_div/SumTmp[9][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_2  ( .A(n153), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[18][2] ), .CO(\u_div/CryTmp[18][3] ), .S(
        \u_div/SumTmp[18][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_1  ( .A(n14), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[12][1] ), .CO(\u_div/CryTmp[12][2] ), .S(
        \u_div/SumTmp[12][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_1  ( .A(n12), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[11][2] ), .S(
        \u_div/SumTmp[11][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_1  ( .A(n4), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[13][1] ), .CO(\u_div/CryTmp[13][2] ), .S(
        \u_div/SumTmp[13][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_1  ( .A(n16), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[14][1] ), .CO(\u_div/CryTmp[14][2] ), .S(
        \u_div/SumTmp[14][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_1  ( .A(n19), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[15][1] ), .CO(\u_div/CryTmp[15][2] ), .S(
        \u_div/SumTmp[15][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_1  ( .A(n3), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[16][1] ), .CO(\u_div/CryTmp[16][2] ), .S(
        \u_div/SumTmp[16][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_1  ( .A(n5), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[17][1] ), .CO(\u_div/CryTmp[17][2] ), .S(
        \u_div/SumTmp[17][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_2  ( .A(n154), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[19][2] ), .CO(\u_div/CryTmp[19][3] ), .S(
        \u_div/SumTmp[19][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_9  ( .A(\u_div/PartRem[1][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[0][9] ), .CO(\u_div/CryTmp[0][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_10  ( .A(\u_div/PartRem[1][10] ), .B(
        \u_div/BInv [10]), .CI(\u_div/CryTmp[0][10] ), .CO(
        \u_div/CryTmp[0][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_10  ( .A(n114), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[10][10] ), .CO(\u_div/CryTmp[10][11] ), .S(
        \u_div/SumTmp[10][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_10  ( .A(n112), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[9][10] ), .CO(\u_div/CryTmp[9][11] ), .S(
        \u_div/SumTmp[9][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_10  ( .A(n110), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[8][10] ), .CO(\u_div/CryTmp[8][11] ), .S(
        \u_div/SumTmp[8][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_10  ( .A(n109), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[7][10] ), .CO(\u_div/CryTmp[7][11] ), .S(
        \u_div/SumTmp[7][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_10  ( .A(n108), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[6][10] ), .CO(\u_div/CryTmp[6][11] ), .S(
        \u_div/SumTmp[6][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_10  ( .A(n107), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[5][10] ), .CO(\u_div/CryTmp[5][11] ), .S(
        \u_div/SumTmp[5][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_10  ( .A(n106), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[4][10] ), .CO(\u_div/CryTmp[4][11] ), .S(
        \u_div/SumTmp[4][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_10  ( .A(n105), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[3][10] ), .CO(\u_div/CryTmp[3][11] ), .S(
        \u_div/SumTmp[3][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_10  ( .A(n104), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[2][10] ), .CO(\u_div/CryTmp[2][11] ), .S(
        \u_div/SumTmp[2][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_10  ( .A(\u_div/PartRem[2][10] ), .B(
        \u_div/BInv [10]), .CI(\u_div/CryTmp[1][10] ), .CO(
        \u_div/CryTmp[1][11] ), .S(\u_div/SumTmp[1][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_9  ( .A(\u_div/PartRem[2][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[1][9] ), .CO(\u_div/CryTmp[1][10] ), .S(\u_div/SumTmp[1][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_9  ( .A(n113), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[10][9] ), .CO(\u_div/CryTmp[10][10] ), .S(
        \u_div/SumTmp[10][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_9  ( .A(n111), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[9][9] ), .CO(\u_div/CryTmp[9][10] ), .S(
        \u_div/SumTmp[9][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_9  ( .A(n103), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[8][9] ), .CO(\u_div/CryTmp[8][10] ), .S(
        \u_div/SumTmp[8][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_9  ( .A(n102), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[7][9] ), .CO(\u_div/CryTmp[7][10] ), .S(
        \u_div/SumTmp[7][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_9  ( .A(n101), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[6][9] ), .CO(\u_div/CryTmp[6][10] ), .S(
        \u_div/SumTmp[6][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_9  ( .A(n100), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[5][9] ), .CO(\u_div/CryTmp[5][10] ), .S(
        \u_div/SumTmp[5][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_9  ( .A(n99), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[4][9] ), .CO(\u_div/CryTmp[4][10] ), .S(
        \u_div/SumTmp[4][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_9  ( .A(n98), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[3][9] ), .CO(\u_div/CryTmp[3][10] ), .S(
        \u_div/SumTmp[3][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_9  ( .A(n97), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[2][9] ), .CO(\u_div/CryTmp[2][10] ), .S(
        \u_div/SumTmp[2][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_9  ( .A(n142), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[11][9] ), .CO(\u_div/CryTmp[11][10] ), .S(
        \u_div/SumTmp[11][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_7  ( .A(\u_div/PartRem[1][7] ), .B(
        \u_div/BInv [7]), .CI(\u_div/CryTmp[0][7] ), .CO(\u_div/CryTmp[0][8] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_8  ( .A(\u_div/PartRem[1][8] ), .B(
        \u_div/BInv [8]), .CI(\u_div/CryTmp[0][8] ), .CO(\u_div/CryTmp[0][9] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_8  ( .A(\u_div/PartRem[2][8] ), .B(
        \u_div/BInv [8]), .CI(\u_div/CryTmp[1][8] ), .CO(\u_div/CryTmp[1][9] ), 
        .S(\u_div/SumTmp[1][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_8  ( .A(n82), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[2][8] ), .CO(\u_div/CryTmp[2][9] ), .S(
        \u_div/SumTmp[2][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_8  ( .A(n88), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[10][8] ), .CO(\u_div/CryTmp[10][9] ), .S(
        \u_div/SumTmp[10][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_8  ( .A(n85), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[9][8] ), .CO(\u_div/CryTmp[9][9] ), .S(
        \u_div/SumTmp[9][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_8  ( .A(n80), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[8][8] ), .CO(\u_div/CryTmp[8][9] ), .S(
        \u_div/SumTmp[8][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_8  ( .A(n79), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[7][8] ), .CO(\u_div/CryTmp[7][9] ), .S(
        \u_div/SumTmp[7][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_8  ( .A(n78), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[6][8] ), .CO(\u_div/CryTmp[6][9] ), .S(
        \u_div/SumTmp[6][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_8  ( .A(n77), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[5][8] ), .CO(\u_div/CryTmp[5][9] ), .S(
        \u_div/SumTmp[5][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_8  ( .A(n76), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[4][8] ), .CO(\u_div/CryTmp[4][9] ), .S(
        \u_div/SumTmp[4][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_8  ( .A(n75), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[3][8] ), .CO(\u_div/CryTmp[3][9] ), .S(
        \u_div/SumTmp[3][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_8  ( .A(n141), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[11][8] ), .CO(\u_div/CryTmp[11][9] ), .S(
        \u_div/SumTmp[11][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_8  ( .A(n91), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[12][8] ), .CO(\u_div/CryTmp[12][9] ), .S(
        \u_div/SumTmp[12][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_7  ( .A(\u_div/PartRem[2][7] ), .B(
        \u_div/BInv [7]), .CI(\u_div/CryTmp[1][7] ), .CO(\u_div/CryTmp[1][8] ), 
        .S(\u_div/SumTmp[1][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_7  ( .A(n81), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[2][7] ), .CO(\u_div/CryTmp[2][8] ), .S(
        \u_div/SumTmp[2][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_7  ( .A(n73), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[3][7] ), .CO(\u_div/CryTmp[3][8] ), .S(
        \u_div/SumTmp[3][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_7  ( .A(n87), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[10][7] ), .CO(\u_div/CryTmp[10][8] ), .S(
        \u_div/SumTmp[10][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_7  ( .A(n84), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[9][7] ), .CO(\u_div/CryTmp[9][8] ), .S(
        \u_div/SumTmp[9][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_7  ( .A(n71), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[8][7] ), .CO(\u_div/CryTmp[8][8] ), .S(
        \u_div/SumTmp[8][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_7  ( .A(n70), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[7][7] ), .CO(\u_div/CryTmp[7][8] ), .S(
        \u_div/SumTmp[7][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_7  ( .A(n69), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[6][7] ), .CO(\u_div/CryTmp[6][8] ), .S(
        \u_div/SumTmp[6][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_7  ( .A(n68), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[5][7] ), .CO(\u_div/CryTmp[5][8] ), .S(
        \u_div/SumTmp[5][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_7  ( .A(n67), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[4][7] ), .CO(\u_div/CryTmp[4][8] ), .S(
        \u_div/SumTmp[4][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_7  ( .A(n140), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[11][7] ), .CO(\u_div/CryTmp[11][8] ), .S(
        \u_div/SumTmp[11][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_7  ( .A(n90), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[12][7] ), .CO(\u_div/CryTmp[12][8] ), .S(
        \u_div/SumTmp[12][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_7  ( .A(n93), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[13][7] ), .CO(\u_div/CryTmp[13][8] ), .S(
        \u_div/SumTmp[13][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_5  ( .A(\u_div/PartRem[1][5] ), .B(
        \u_div/BInv [5]), .CI(\u_div/CryTmp[0][5] ), .CO(\u_div/CryTmp[0][6] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_6  ( .A(\u_div/PartRem[1][6] ), .B(
        \u_div/BInv [6]), .CI(\u_div/CryTmp[0][6] ), .CO(\u_div/CryTmp[0][7] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_6  ( .A(\u_div/PartRem[2][6] ), .B(
        \u_div/BInv [6]), .CI(\u_div/CryTmp[1][6] ), .CO(\u_div/CryTmp[1][7] ), 
        .S(\u_div/SumTmp[1][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_6  ( .A(n74), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[2][6] ), .CO(\u_div/CryTmp[2][7] ), .S(
        \u_div/SumTmp[2][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_6  ( .A(n72), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[3][6] ), .CO(\u_div/CryTmp[3][7] ), .S(
        \u_div/SumTmp[3][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_6  ( .A(n66), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[4][6] ), .CO(\u_div/CryTmp[4][7] ), .S(
        \u_div/SumTmp[4][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_6  ( .A(n139), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[11][6] ), .CO(\u_div/CryTmp[11][7] ), .S(
        \u_div/SumTmp[11][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_6  ( .A(n86), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[10][6] ), .CO(\u_div/CryTmp[10][7] ), .S(
        \u_div/SumTmp[10][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_6  ( .A(n83), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[9][6] ), .CO(\u_div/CryTmp[9][7] ), .S(
        \u_div/SumTmp[9][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_6  ( .A(n65), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[8][6] ), .CO(\u_div/CryTmp[8][7] ), .S(
        \u_div/SumTmp[8][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_6  ( .A(n64), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[7][6] ), .CO(\u_div/CryTmp[7][7] ), .S(
        \u_div/SumTmp[7][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_6  ( .A(n63), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[6][6] ), .CO(\u_div/CryTmp[6][7] ), .S(
        \u_div/SumTmp[6][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_6  ( .A(n62), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[5][6] ), .CO(\u_div/CryTmp[5][7] ), .S(
        \u_div/SumTmp[5][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_6  ( .A(n89), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[12][6] ), .CO(\u_div/CryTmp[12][7] ), .S(
        \u_div/SumTmp[12][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_6  ( .A(n92), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[13][6] ), .CO(\u_div/CryTmp[13][7] ), .S(
        \u_div/SumTmp[13][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_6  ( .A(n94), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[14][6] ), .CO(\u_div/CryTmp[14][7] ), .S(
        \u_div/SumTmp[14][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_5  ( .A(\u_div/PartRem[2][5] ), .B(
        \u_div/BInv [5]), .CI(\u_div/CryTmp[1][5] ), .CO(\u_div/CryTmp[1][6] ), 
        .S(\u_div/SumTmp[1][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_5  ( .A(n42), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[2][5] ), .CO(\u_div/CryTmp[2][6] ), .S(
        \u_div/SumTmp[2][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_5  ( .A(n41), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[3][5] ), .CO(\u_div/CryTmp[3][6] ), .S(
        \u_div/SumTmp[3][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_5  ( .A(n40), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[4][5] ), .CO(\u_div/CryTmp[4][6] ), .S(
        \u_div/SumTmp[4][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_5  ( .A(n38), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[5][5] ), .CO(\u_div/CryTmp[5][6] ), .S(
        \u_div/SumTmp[5][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_5  ( .A(n138), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[11][5] ), .CO(\u_div/CryTmp[11][6] ), .S(
        \u_div/SumTmp[11][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_5  ( .A(n47), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[10][5] ), .CO(\u_div/CryTmp[10][6] ), .S(
        \u_div/SumTmp[10][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_5  ( .A(n44), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[9][5] ), .CO(\u_div/CryTmp[9][6] ), .S(
        \u_div/SumTmp[9][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_5  ( .A(n36), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[8][5] ), .CO(\u_div/CryTmp[8][6] ), .S(
        \u_div/SumTmp[8][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_5  ( .A(n35), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[7][5] ), .CO(\u_div/CryTmp[7][6] ), .S(
        \u_div/SumTmp[7][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_5  ( .A(n34), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[6][5] ), .CO(\u_div/CryTmp[6][6] ), .S(
        \u_div/SumTmp[6][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_5  ( .A(n50), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[12][5] ), .CO(\u_div/CryTmp[12][6] ), .S(
        \u_div/SumTmp[12][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_5  ( .A(n53), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[13][5] ), .CO(\u_div/CryTmp[13][6] ), .S(
        \u_div/SumTmp[13][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_5  ( .A(n56), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[14][5] ), .CO(\u_div/CryTmp[14][6] ), .S(
        \u_div/SumTmp[14][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_5  ( .A(n58), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[15][5] ), .CO(\u_div/CryTmp[15][6] ), .S(
        \u_div/SumTmp[15][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/BInv [4]), .CI(\u_div/CryTmp[1][4] ), .CO(\u_div/CryTmp[1][5] ), 
        .S(\u_div/SumTmp[1][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_4  ( .A(n130), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[2][4] ), .CO(\u_div/CryTmp[2][5] ), .S(
        \u_div/SumTmp[2][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_4  ( .A(n129), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[3][4] ), .CO(\u_div/CryTmp[3][5] ), .S(
        \u_div/SumTmp[3][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_4  ( .A(n39), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[4][4] ), .CO(\u_div/CryTmp[4][5] ), .S(
        \u_div/SumTmp[4][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_4  ( .A(n37), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[5][4] ), .CO(\u_div/CryTmp[5][5] ), .S(
        \u_div/SumTmp[5][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_4  ( .A(n33), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[6][4] ), .CO(\u_div/CryTmp[6][5] ), .S(
        \u_div/SumTmp[6][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_4  ( .A(n137), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[11][4] ), .CO(\u_div/CryTmp[11][5] ), .S(
        \u_div/SumTmp[11][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_4  ( .A(n46), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[10][4] ), .CO(\u_div/CryTmp[10][5] ), .S(
        \u_div/SumTmp[10][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_4  ( .A(n43), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[9][4] ), .CO(\u_div/CryTmp[9][5] ), .S(
        \u_div/SumTmp[9][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_4  ( .A(n32), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[8][4] ), .CO(\u_div/CryTmp[8][5] ), .S(
        \u_div/SumTmp[8][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_4  ( .A(n31), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[7][4] ), .CO(\u_div/CryTmp[7][5] ), .S(
        \u_div/SumTmp[7][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_4  ( .A(n49), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[12][4] ), .CO(\u_div/CryTmp[12][5] ), .S(
        \u_div/SumTmp[12][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_4  ( .A(n52), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[13][4] ), .CO(\u_div/CryTmp[13][5] ), .S(
        \u_div/SumTmp[13][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_4  ( .A(n55), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[14][4] ), .CO(\u_div/CryTmp[14][5] ), .S(
        \u_div/SumTmp[14][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_4  ( .A(n57), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[15][4] ), .CO(\u_div/CryTmp[15][5] ), .S(
        \u_div/SumTmp[15][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_4  ( .A(n59), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[16][4] ), .CO(\u_div/CryTmp[16][5] ), .S(
        \u_div/SumTmp[16][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_3  ( .A(\u_div/PartRem[1][3] ), .B(
        \u_div/BInv [3]), .CI(\u_div/CryTmp[0][3] ), .CO(\u_div/CryTmp[0][4] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_4  ( .A(\u_div/PartRem[1][4] ), .B(
        \u_div/BInv [4]), .CI(\u_div/CryTmp[0][4] ), .CO(\u_div/CryTmp[0][5] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/BInv [3]), .CI(\u_div/CryTmp[1][3] ), .CO(\u_div/CryTmp[1][4] ), 
        .S(\u_div/SumTmp[1][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_3  ( .A(n156), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[2][3] ), .CO(\u_div/CryTmp[2][4] ), .S(
        \u_div/SumTmp[2][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_3  ( .A(n127), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[5][3] ), .CO(\u_div/CryTmp[5][4] ), .S(
        \u_div/SumTmp[5][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_3  ( .A(n126), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[6][3] ), .CO(\u_div/CryTmp[6][4] ), .S(
        \u_div/SumTmp[6][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_3  ( .A(n125), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[7][3] ), .CO(\u_div/CryTmp[7][4] ), .S(
        \u_div/SumTmp[7][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_3  ( .A(n136), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[11][3] ), .CO(\u_div/CryTmp[11][4] ), .S(
        \u_div/SumTmp[11][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_3  ( .A(n45), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[10][3] ), .CO(\u_div/CryTmp[10][4] ), .S(
        \u_div/SumTmp[10][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_3  ( .A(n131), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[9][3] ), .CO(\u_div/CryTmp[9][4] ), .S(
        \u_div/SumTmp[9][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_3  ( .A(n124), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[8][3] ), .CO(\u_div/CryTmp[8][4] ), .S(
        \u_div/SumTmp[8][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_3  ( .A(n48), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[12][3] ), .CO(\u_div/CryTmp[12][4] ), .S(
        \u_div/SumTmp[12][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_3  ( .A(n51), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[13][3] ), .CO(\u_div/CryTmp[13][4] ), .S(
        \u_div/SumTmp[13][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_3  ( .A(n54), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[14][3] ), .CO(\u_div/CryTmp[14][4] ), .S(
        \u_div/SumTmp[14][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_3  ( .A(n132), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[15][3] ), .CO(\u_div/CryTmp[15][4] ), .S(
        \u_div/SumTmp[15][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_3  ( .A(n133), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[16][3] ), .CO(\u_div/CryTmp[16][4] ), .S(
        \u_div/SumTmp[16][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_3  ( .A(n134), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[17][3] ), .CO(\u_div/CryTmp[17][4] ), .S(
        \u_div/SumTmp[17][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_2  ( .A(n123), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[11][2] ), .CO(\u_div/CryTmp[11][3] ), .S(
        \u_div/SumTmp[11][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_2  ( .A(n119), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[12][2] ), .CO(\u_div/CryTmp[12][3] ), .S(
        \u_div/SumTmp[12][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_2  ( .A(n120), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[13][2] ), .CO(\u_div/CryTmp[13][3] ), .S(
        \u_div/SumTmp[13][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_2  ( .A(n121), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[14][2] ), .CO(\u_div/CryTmp[14][3] ), .S(
        \u_div/SumTmp[14][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_2  ( .A(n122), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[15][2] ), .CO(\u_div/CryTmp[15][3] ), .S(
        \u_div/SumTmp[15][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_2  ( .A(n151), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[16][2] ), .CO(\u_div/CryTmp[16][3] ), .S(
        \u_div/SumTmp[16][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_2  ( .A(n152), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[17][2] ), .CO(\u_div/CryTmp[17][3] ), .S(
        \u_div/SumTmp[17][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_5  ( .A(n60), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[16][5] ), .CO(\u_div/CryTmp[16][6] ), .S(
        \u_div/SumTmp[16][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_3  ( .A(n135), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[18][3] ), .CO(\u_div/CryTmp[18][4] ), .S(
        \u_div/SumTmp[18][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_10  ( .A(n143), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[11][10] ), .CO(\u_div/CryTmp[11][11] ), .S(
        \u_div/SumTmp[11][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_8  ( .A(n116), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[13][8] ), .CO(\u_div/CryTmp[13][9] ), .S(
        \u_div/SumTmp[13][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_6  ( .A(n96), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[15][6] ), .CO(\u_div/CryTmp[15][7] ), .S(
        \u_div/SumTmp[15][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_7  ( .A(n95), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[14][7] ), .CO(\u_div/CryTmp[14][8] ), .S(
        \u_div/SumTmp[14][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_4  ( .A(n61), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[17][4] ), .CO(\u_div/CryTmp[17][5] ), .S(
        \u_div/SumTmp[17][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_1  ( .A(n30), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[2][1] ), .CO(\u_div/CryTmp[0][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/BInv [2]), .CI(\u_div/CryTmp[0][2] ), .CO(\u_div/CryTmp[0][3] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_12_9  ( .A(n115), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[12][9] ), .CO(\u_div/CryTmp[12][10] ), .S(
        \u_div/SumTmp[12][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_11  ( .A(\u_div/PartRem[10][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[9][11] ), .CO(
        \u_div/CryTmp[9][12] ), .S(\u_div/SumTmp[9][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_11  ( .A(\u_div/PartRem[9][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[8][11] ), .CO(
        \u_div/CryTmp[8][12] ), .S(\u_div/SumTmp[8][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_11  ( .A(\u_div/PartRem[8][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[7][11] ), .CO(
        \u_div/CryTmp[7][12] ), .S(\u_div/SumTmp[7][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_11  ( .A(\u_div/PartRem[7][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[6][11] ), .CO(
        \u_div/CryTmp[6][12] ), .S(\u_div/SumTmp[6][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_11  ( .A(\u_div/PartRem[6][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[5][11] ), .CO(
        \u_div/CryTmp[5][12] ), .S(\u_div/SumTmp[5][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_11  ( .A(\u_div/PartRem[5][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[4][11] ), .CO(
        \u_div/CryTmp[4][12] ), .S(\u_div/SumTmp[4][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_11  ( .A(\u_div/PartRem[4][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[3][11] ), .CO(
        \u_div/CryTmp[3][12] ), .S(\u_div/SumTmp[3][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_11  ( .A(\u_div/PartRem[3][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[2][11] ), .CO(
        \u_div/CryTmp[2][12] ), .S(\u_div/SumTmp[2][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_11  ( .A(\u_div/PartRem[2][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[1][11] ), .CO(
        \u_div/CryTmp[1][12] ), .S(\u_div/SumTmp[1][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_11  ( .A(\u_div/PartRem[1][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[0][11] ), .CO(
        \u_div/CryTmp[0][12] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        \u_div/BInv [1]), .CI(\u_div/CryTmp[2][1] ), .CO(\u_div/CryTmp[1][2] ), 
        .S(\u_div/SumTmp[1][1] ) );
  ADDFX4 \u_div/u_fa_PartRem_0_10_11  ( .A(\u_div/PartRem[11][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[10][11] ), .CO(
        \u_div/CryTmp[10][12] ), .S(\u_div/SumTmp[10][11] ) );
  INVX4 U1 ( .A(b[2]), .Y(\u_div/BInv [2]) );
  INVX4 U2 ( .A(b[4]), .Y(\u_div/BInv [4]) );
  INVX4 U3 ( .A(b[3]), .Y(\u_div/BInv [3]) );
  INVX4 U4 ( .A(b[6]), .Y(\u_div/BInv [6]) );
  INVX4 U5 ( .A(b[5]), .Y(\u_div/BInv [5]) );
  MX2X1 U6 ( .A(a[3]), .B(\u_div/SumTmp[3][0] ), .S0(quotient[3]), .Y(n1) );
  MX2X1 U7 ( .A(a[4]), .B(\u_div/SumTmp[4][0] ), .S0(quotient[4]), .Y(n2) );
  MX2X1 U8 ( .A(a[17]), .B(\u_div/SumTmp[17][0] ), .S0(n203), .Y(n3) );
  MX2X1 U9 ( .A(a[14]), .B(\u_div/SumTmp[14][0] ), .S0(n117), .Y(n4) );
  MX2X1 U10 ( .A(a[18]), .B(\u_div/SumTmp[18][0] ), .S0(n204), .Y(n5) );
  MX2X1 U11 ( .A(a[11]), .B(\u_div/SumTmp[11][0] ), .S0(n198), .Y(n6) );
  MX2X1 U12 ( .A(a[9]), .B(\u_div/SumTmp[9][0] ), .S0(quotient[9]), .Y(n7) );
  MX2X1 U13 ( .A(a[8]), .B(\u_div/SumTmp[8][0] ), .S0(quotient[8]), .Y(n8) );
  MX2X1 U14 ( .A(a[7]), .B(\u_div/SumTmp[7][0] ), .S0(quotient[7]), .Y(n9) );
  MX2X1 U15 ( .A(a[6]), .B(\u_div/SumTmp[6][0] ), .S0(quotient[6]), .Y(n10) );
  MX2X1 U16 ( .A(a[5]), .B(\u_div/SumTmp[5][0] ), .S0(quotient[5]), .Y(n11) );
  MX2X1 U17 ( .A(a[12]), .B(\u_div/SumTmp[12][0] ), .S0(n227), .Y(n12) );
  MX2X1 U18 ( .A(a[19]), .B(\u_div/SumTmp[19][0] ), .S0(n206), .Y(n13) );
  MX2X1 U19 ( .A(a[13]), .B(\u_div/SumTmp[13][0] ), .S0(n200), .Y(n14) );
  MX2X1 U20 ( .A(a[10]), .B(\u_div/SumTmp[10][0] ), .S0(\u_div/CryTmp[10][12] ), .Y(n15) );
  MX2X1 U21 ( .A(a[15]), .B(\u_div/SumTmp[15][0] ), .S0(n201), .Y(n16) );
  MX2X1 U22 ( .A(a[21]), .B(\u_div/SumTmp[21][0] ), .S0(n208), .Y(n17) );
  MX2X1 U23 ( .A(a[20]), .B(\u_div/SumTmp[20][0] ), .S0(n207), .Y(n18) );
  MX2X1 U24 ( .A(a[16]), .B(\u_div/SumTmp[16][0] ), .S0(n202), .Y(n19) );
  MX2X1 U25 ( .A(n184), .B(n194), .S0(quotient[1]), .Y(n20) );
  MX2X1 U26 ( .A(n173), .B(n183), .S0(quotient[2]), .Y(n21) );
  MX2X1 U27 ( .A(n159), .B(n160), .S0(quotient[9]), .Y(n22) );
  MX2X1 U28 ( .A(n161), .B(n162), .S0(quotient[8]), .Y(n23) );
  MX2X1 U29 ( .A(n163), .B(n164), .S0(quotient[7]), .Y(n24) );
  MX2X1 U30 ( .A(n165), .B(n166), .S0(quotient[6]), .Y(n25) );
  MX2X1 U31 ( .A(n167), .B(n168), .S0(quotient[5]), .Y(n26) );
  MX2X1 U32 ( .A(n171), .B(n172), .S0(quotient[3]), .Y(n27) );
  MX2X1 U33 ( .A(n169), .B(n170), .S0(quotient[4]), .Y(n28) );
  MX2X1 U34 ( .A(n197), .B(n205), .S0(\u_div/CryTmp[10][12] ), .Y(n29) );
  XNOR2XL U35 ( .A(\u_div/CryTmp[2][1] ), .B(a[4]), .Y(\u_div/SumTmp[4][0] )
         );
  CLKINVX3 U36 ( .A(b[7]), .Y(\u_div/BInv [7]) );
  CLKINVX3 U37 ( .A(b[8]), .Y(\u_div/BInv [8]) );
  CLKINVX3 U38 ( .A(b[9]), .Y(\u_div/BInv [9]) );
  INVX1 U39 ( .A(\u_div/SumTmp[4][11] ), .Y(n170) );
  INVX1 U40 ( .A(\u_div/SumTmp[5][11] ), .Y(n168) );
  INVX1 U41 ( .A(\u_div/SumTmp[6][11] ), .Y(n166) );
  INVX1 U42 ( .A(\u_div/SumTmp[7][11] ), .Y(n164) );
  INVX1 U43 ( .A(\u_div/SumTmp[8][11] ), .Y(n162) );
  INVX1 U44 ( .A(\u_div/SumTmp[9][11] ), .Y(n160) );
  INVX1 U45 ( .A(\u_div/SumTmp[10][11] ), .Y(n205) );
  INVX1 U46 ( .A(\u_div/SumTmp[2][11] ), .Y(n183) );
  INVX1 U47 ( .A(\u_div/SumTmp[3][11] ), .Y(n172) );
  NAND2X1 U48 ( .A(quotient[2]), .B(b[0]), .Y(n182) );
  NOR2BX1 U49 ( .AN(quotient[1]), .B(\u_div/CryTmp[2][1] ), .Y(n30) );
  INVX1 U50 ( .A(\u_div/SumTmp[1][11] ), .Y(n194) );
  INVX1 U51 ( .A(n197), .Y(\u_div/PartRem[11][11] ) );
  CLKINVX3 U52 ( .A(n217), .Y(n201) );
  NAND2BX1 U53 ( .AN(n218), .B(\u_div/CryTmp[15][7] ), .Y(n217) );
  INVX1 U54 ( .A(n182), .Y(\u_div/PartRem[2][1] ) );
  NAND2BX1 U55 ( .AN(\u_div/CryTmp[0][12] ), .B(n20), .Y(quotient[0]) );
  INVX1 U56 ( .A(n184), .Y(\u_div/PartRem[2][11] ) );
  INVX1 U57 ( .A(n173), .Y(\u_div/PartRem[3][11] ) );
  INVX1 U58 ( .A(n171), .Y(\u_div/PartRem[4][11] ) );
  INVX1 U59 ( .A(n169), .Y(\u_div/PartRem[5][11] ) );
  INVX1 U60 ( .A(n167), .Y(\u_div/PartRem[6][11] ) );
  INVX1 U61 ( .A(n165), .Y(\u_div/PartRem[7][11] ) );
  INVX1 U62 ( .A(n163), .Y(\u_div/PartRem[8][11] ) );
  INVX1 U63 ( .A(n161), .Y(\u_div/PartRem[9][11] ) );
  INVX1 U64 ( .A(n159), .Y(\u_div/PartRem[10][11] ) );
  MXI2X1 U65 ( .A(n130), .B(\u_div/SumTmp[2][4] ), .S0(quotient[2]), .Y(n178)
         );
  MX2X1 U66 ( .A(n124), .B(\u_div/SumTmp[8][3] ), .S0(quotient[8]), .Y(n31) );
  MX2X1 U67 ( .A(n131), .B(\u_div/SumTmp[9][3] ), .S0(quotient[9]), .Y(n32) );
  MX2X1 U68 ( .A(n125), .B(\u_div/SumTmp[7][3] ), .S0(quotient[7]), .Y(n33) );
  MX2X1 U69 ( .A(n31), .B(\u_div/SumTmp[7][4] ), .S0(quotient[7]), .Y(n34) );
  MX2X1 U70 ( .A(n32), .B(\u_div/SumTmp[8][4] ), .S0(quotient[8]), .Y(n35) );
  MX2X1 U71 ( .A(n43), .B(\u_div/SumTmp[9][4] ), .S0(quotient[9]), .Y(n36) );
  MX2X1 U72 ( .A(n126), .B(\u_div/SumTmp[6][3] ), .S0(quotient[6]), .Y(n37) );
  MX2X1 U73 ( .A(n33), .B(\u_div/SumTmp[6][4] ), .S0(quotient[6]), .Y(n38) );
  MX2X1 U74 ( .A(n127), .B(\u_div/SumTmp[5][3] ), .S0(quotient[5]), .Y(n39) );
  MX2X1 U75 ( .A(n37), .B(\u_div/SumTmp[5][4] ), .S0(quotient[5]), .Y(n40) );
  MX2X1 U76 ( .A(n39), .B(\u_div/SumTmp[4][4] ), .S0(quotient[4]), .Y(n41) );
  MX2X1 U77 ( .A(n129), .B(\u_div/SumTmp[3][4] ), .S0(quotient[3]), .Y(n42) );
  MX2X1 U78 ( .A(n45), .B(\u_div/SumTmp[10][3] ), .S0(\u_div/CryTmp[10][12] ), 
        .Y(n43) );
  MX2X1 U79 ( .A(n46), .B(\u_div/SumTmp[10][4] ), .S0(\u_div/CryTmp[10][12] ), 
        .Y(n44) );
  MX2X1 U80 ( .A(n123), .B(\u_div/SumTmp[11][2] ), .S0(n198), .Y(n45) );
  MX2X1 U81 ( .A(n136), .B(\u_div/SumTmp[11][3] ), .S0(n198), .Y(n46) );
  MX2X1 U82 ( .A(n137), .B(\u_div/SumTmp[11][4] ), .S0(n198), .Y(n47) );
  MX2X1 U83 ( .A(n120), .B(\u_div/SumTmp[13][2] ), .S0(n200), .Y(n48) );
  MX2X1 U84 ( .A(n51), .B(\u_div/SumTmp[13][3] ), .S0(n200), .Y(n49) );
  MX2X1 U85 ( .A(n52), .B(\u_div/SumTmp[13][4] ), .S0(n200), .Y(n50) );
  MX2X1 U86 ( .A(n121), .B(\u_div/SumTmp[14][2] ), .S0(n117), .Y(n51) );
  MX2X1 U87 ( .A(n54), .B(\u_div/SumTmp[14][3] ), .S0(n117), .Y(n52) );
  MX2X1 U88 ( .A(n55), .B(\u_div/SumTmp[14][4] ), .S0(n117), .Y(n53) );
  MX2X1 U89 ( .A(n122), .B(\u_div/SumTmp[15][2] ), .S0(n201), .Y(n54) );
  MX2X1 U90 ( .A(n132), .B(\u_div/SumTmp[15][3] ), .S0(n201), .Y(n55) );
  MX2X1 U91 ( .A(n57), .B(\u_div/SumTmp[15][4] ), .S0(n201), .Y(n56) );
  MX2X1 U92 ( .A(n133), .B(\u_div/SumTmp[16][3] ), .S0(n202), .Y(n57) );
  MX2X1 U93 ( .A(n59), .B(\u_div/SumTmp[16][4] ), .S0(n202), .Y(n58) );
  MX2X1 U94 ( .A(n134), .B(\u_div/SumTmp[17][3] ), .S0(n203), .Y(n59) );
  MX2X1 U95 ( .A(n61), .B(\u_div/SumTmp[17][4] ), .S0(n203), .Y(n60) );
  MX2X1 U96 ( .A(n135), .B(\u_div/SumTmp[18][3] ), .S0(n204), .Y(n61) );
  MXI2X1 U97 ( .A(n42), .B(\u_div/SumTmp[2][5] ), .S0(quotient[2]), .Y(n177)
         );
  MXI2X1 U98 ( .A(n81), .B(\u_div/SumTmp[2][7] ), .S0(quotient[2]), .Y(n175)
         );
  MXI2X1 U99 ( .A(n74), .B(\u_div/SumTmp[2][6] ), .S0(quotient[2]), .Y(n176)
         );
  MXI2X1 U100 ( .A(n179), .B(n190), .S0(quotient[1]), .Y(\u_div/PartRem[1][5] ) );
  INVX1 U101 ( .A(\u_div/SumTmp[1][4] ), .Y(n190) );
  MXI2X1 U102 ( .A(n177), .B(n188), .S0(quotient[1]), .Y(\u_div/PartRem[1][7] ) );
  INVX1 U103 ( .A(\u_div/SumTmp[1][6] ), .Y(n188) );
  MX2X1 U104 ( .A(n34), .B(\u_div/SumTmp[6][5] ), .S0(quotient[6]), .Y(n62) );
  MX2X1 U105 ( .A(n35), .B(\u_div/SumTmp[7][5] ), .S0(quotient[7]), .Y(n63) );
  MX2X1 U106 ( .A(n36), .B(\u_div/SumTmp[8][5] ), .S0(quotient[8]), .Y(n64) );
  MX2X1 U107 ( .A(n44), .B(\u_div/SumTmp[9][5] ), .S0(quotient[9]), .Y(n65) );
  MX2X1 U108 ( .A(n38), .B(\u_div/SumTmp[5][5] ), .S0(quotient[5]), .Y(n66) );
  MX2X1 U109 ( .A(n62), .B(\u_div/SumTmp[5][6] ), .S0(quotient[5]), .Y(n67) );
  MX2X1 U110 ( .A(n63), .B(\u_div/SumTmp[6][6] ), .S0(quotient[6]), .Y(n68) );
  MX2X1 U111 ( .A(n64), .B(\u_div/SumTmp[7][6] ), .S0(quotient[7]), .Y(n69) );
  MX2X1 U112 ( .A(n65), .B(\u_div/SumTmp[8][6] ), .S0(quotient[8]), .Y(n70) );
  MX2X1 U113 ( .A(n83), .B(\u_div/SumTmp[9][6] ), .S0(quotient[9]), .Y(n71) );
  MX2X1 U114 ( .A(n40), .B(\u_div/SumTmp[4][5] ), .S0(quotient[4]), .Y(n72) );
  MX2X1 U115 ( .A(n66), .B(\u_div/SumTmp[4][6] ), .S0(quotient[4]), .Y(n73) );
  MX2X1 U116 ( .A(n41), .B(\u_div/SumTmp[3][5] ), .S0(quotient[3]), .Y(n74) );
  MX2X1 U117 ( .A(n67), .B(\u_div/SumTmp[4][7] ), .S0(quotient[4]), .Y(n75) );
  MX2X1 U118 ( .A(n68), .B(\u_div/SumTmp[5][7] ), .S0(quotient[5]), .Y(n76) );
  MX2X1 U119 ( .A(n69), .B(\u_div/SumTmp[6][7] ), .S0(quotient[6]), .Y(n77) );
  MX2X1 U120 ( .A(n70), .B(\u_div/SumTmp[7][7] ), .S0(quotient[7]), .Y(n78) );
  MX2X1 U121 ( .A(n71), .B(\u_div/SumTmp[8][7] ), .S0(quotient[8]), .Y(n79) );
  MX2X1 U122 ( .A(n84), .B(\u_div/SumTmp[9][7] ), .S0(quotient[9]), .Y(n80) );
  MX2X1 U123 ( .A(n72), .B(\u_div/SumTmp[3][6] ), .S0(quotient[3]), .Y(n81) );
  MX2X1 U124 ( .A(n73), .B(\u_div/SumTmp[3][7] ), .S0(quotient[3]), .Y(n82) );
  MX2X1 U125 ( .A(n47), .B(\u_div/SumTmp[10][5] ), .S0(\u_div/CryTmp[10][12] ), 
        .Y(n83) );
  MX2X1 U126 ( .A(n86), .B(\u_div/SumTmp[10][6] ), .S0(\u_div/CryTmp[10][12] ), 
        .Y(n84) );
  MX2X1 U127 ( .A(n87), .B(\u_div/SumTmp[10][7] ), .S0(\u_div/CryTmp[10][12] ), 
        .Y(n85) );
  MX2X1 U128 ( .A(n138), .B(\u_div/SumTmp[11][5] ), .S0(n198), .Y(n86) );
  MX2X1 U129 ( .A(n139), .B(\u_div/SumTmp[11][6] ), .S0(n198), .Y(n87) );
  MX2X1 U130 ( .A(n140), .B(\u_div/SumTmp[11][7] ), .S0(n198), .Y(n88) );
  MX2X1 U131 ( .A(n53), .B(\u_div/SumTmp[13][5] ), .S0(n200), .Y(n89) );
  MX2X1 U132 ( .A(n92), .B(\u_div/SumTmp[13][6] ), .S0(n200), .Y(n90) );
  MX2X1 U133 ( .A(n93), .B(\u_div/SumTmp[13][7] ), .S0(n200), .Y(n91) );
  MX2X1 U134 ( .A(n56), .B(\u_div/SumTmp[14][5] ), .S0(n117), .Y(n92) );
  MX2X1 U135 ( .A(n94), .B(\u_div/SumTmp[14][6] ), .S0(n117), .Y(n93) );
  MX2X1 U136 ( .A(n58), .B(\u_div/SumTmp[15][5] ), .S0(n201), .Y(n94) );
  MX2X1 U137 ( .A(n96), .B(\u_div/SumTmp[15][6] ), .S0(n201), .Y(n95) );
  MX2X1 U138 ( .A(n60), .B(\u_div/SumTmp[16][5] ), .S0(n202), .Y(n96) );
  MXI2X1 U139 ( .A(n105), .B(\u_div/SumTmp[3][10] ), .S0(quotient[3]), .Y(n173) );
  MXI2X1 U140 ( .A(n106), .B(\u_div/SumTmp[4][10] ), .S0(quotient[4]), .Y(n171) );
  MXI2X1 U141 ( .A(n107), .B(\u_div/SumTmp[5][10] ), .S0(quotient[5]), .Y(n169) );
  MXI2X1 U142 ( .A(n108), .B(\u_div/SumTmp[6][10] ), .S0(quotient[6]), .Y(n167) );
  MXI2X1 U143 ( .A(n109), .B(\u_div/SumTmp[7][10] ), .S0(quotient[7]), .Y(n165) );
  MXI2X1 U144 ( .A(n110), .B(\u_div/SumTmp[8][10] ), .S0(quotient[8]), .Y(n163) );
  MXI2X1 U145 ( .A(n112), .B(\u_div/SumTmp[9][10] ), .S0(quotient[9]), .Y(n161) );
  MXI2X1 U146 ( .A(n97), .B(\u_div/SumTmp[2][9] ), .S0(quotient[2]), .Y(n185)
         );
  MXI2X1 U147 ( .A(n82), .B(\u_div/SumTmp[2][8] ), .S0(quotient[2]), .Y(n174)
         );
  MXI2X1 U148 ( .A(n104), .B(\u_div/SumTmp[2][10] ), .S0(quotient[2]), .Y(n184) );
  MXI2X1 U149 ( .A(n114), .B(\u_div/SumTmp[10][10] ), .S0(
        \u_div/CryTmp[10][12] ), .Y(n159) );
  MXI2X1 U150 ( .A(n143), .B(\u_div/SumTmp[11][10] ), .S0(n198), .Y(n197) );
  MXI2X1 U151 ( .A(n175), .B(n186), .S0(quotient[1]), .Y(\u_div/PartRem[1][9] ) );
  INVX1 U152 ( .A(\u_div/SumTmp[1][8] ), .Y(n186) );
  MX2X1 U153 ( .A(n75), .B(\u_div/SumTmp[3][8] ), .S0(quotient[3]), .Y(n97) );
  MX2X1 U154 ( .A(n76), .B(\u_div/SumTmp[4][8] ), .S0(quotient[4]), .Y(n98) );
  MX2X1 U155 ( .A(n77), .B(\u_div/SumTmp[5][8] ), .S0(quotient[5]), .Y(n99) );
  MX2X1 U156 ( .A(n78), .B(\u_div/SumTmp[6][8] ), .S0(quotient[6]), .Y(n100)
         );
  MX2X1 U157 ( .A(n79), .B(\u_div/SumTmp[7][8] ), .S0(quotient[7]), .Y(n101)
         );
  MX2X1 U158 ( .A(n80), .B(\u_div/SumTmp[8][8] ), .S0(quotient[8]), .Y(n102)
         );
  MX2X1 U159 ( .A(n85), .B(\u_div/SumTmp[9][8] ), .S0(quotient[9]), .Y(n103)
         );
  MX2X1 U160 ( .A(n98), .B(\u_div/SumTmp[3][9] ), .S0(quotient[3]), .Y(n104)
         );
  MX2X1 U161 ( .A(n99), .B(\u_div/SumTmp[4][9] ), .S0(quotient[4]), .Y(n105)
         );
  MX2X1 U162 ( .A(n100), .B(\u_div/SumTmp[5][9] ), .S0(quotient[5]), .Y(n106)
         );
  MX2X1 U163 ( .A(n101), .B(\u_div/SumTmp[6][9] ), .S0(quotient[6]), .Y(n107)
         );
  MX2X1 U164 ( .A(n102), .B(\u_div/SumTmp[7][9] ), .S0(quotient[7]), .Y(n108)
         );
  MX2X1 U165 ( .A(n103), .B(\u_div/SumTmp[8][9] ), .S0(quotient[8]), .Y(n109)
         );
  MX2X1 U166 ( .A(n111), .B(\u_div/SumTmp[9][9] ), .S0(quotient[9]), .Y(n110)
         );
  MX2X1 U167 ( .A(n88), .B(\u_div/SumTmp[10][8] ), .S0(\u_div/CryTmp[10][12] ), 
        .Y(n111) );
  MX2X1 U168 ( .A(n113), .B(\u_div/SumTmp[10][9] ), .S0(\u_div/CryTmp[10][12] ), .Y(n112) );
  MX2X1 U169 ( .A(n141), .B(\u_div/SumTmp[11][8] ), .S0(n198), .Y(n113) );
  MX2X1 U170 ( .A(n142), .B(\u_div/SumTmp[11][9] ), .S0(n198), .Y(n114) );
  MX2X1 U171 ( .A(n116), .B(\u_div/SumTmp[13][8] ), .S0(n200), .Y(n115) );
  MX2X1 U172 ( .A(n95), .B(\u_div/SumTmp[14][7] ), .S0(n117), .Y(n116) );
  MXI2X1 U173 ( .A(n185), .B(n195), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][11] ) );
  INVX1 U174 ( .A(\u_div/SumTmp[1][10] ), .Y(n195) );
  CLKINVX3 U175 ( .A(n213), .Y(n198) );
  NAND2BX1 U176 ( .AN(b[11]), .B(\u_div/CryTmp[11][11] ), .Y(n213) );
  CLKINVX3 U177 ( .A(n215), .Y(n200) );
  NAND2BX1 U178 ( .AN(n216), .B(\u_div/CryTmp[13][9] ), .Y(n215) );
  AND2X2 U179 ( .A(\u_div/CryTmp[14][8] ), .B(n150), .Y(n117) );
  CLKINVX3 U180 ( .A(n219), .Y(n202) );
  NAND3BX1 U181 ( .AN(n218), .B(\u_div/BInv [6]), .C(\u_div/CryTmp[16][6] ), 
        .Y(n219) );
  INVX1 U182 ( .A(n220), .Y(n203) );
  NAND2BX1 U183 ( .AN(n221), .B(\u_div/CryTmp[17][5] ), .Y(n220) );
  INVX1 U184 ( .A(n222), .Y(n204) );
  NAND3BX1 U185 ( .AN(n221), .B(\u_div/BInv [4]), .C(\u_div/CryTmp[18][4] ), 
        .Y(n222) );
  NAND2X1 U186 ( .A(n150), .B(\u_div/BInv [7]), .Y(n218) );
  INVX1 U187 ( .A(n223), .Y(n206) );
  NAND2BX1 U188 ( .AN(n209), .B(\u_div/CryTmp[19][3] ), .Y(n223) );
  MX2X1 U189 ( .A(n12), .B(\u_div/SumTmp[11][1] ), .S0(n198), .Y(n118) );
  MX2X1 U190 ( .A(n4), .B(\u_div/SumTmp[13][1] ), .S0(n200), .Y(n119) );
  MX2X1 U191 ( .A(n16), .B(\u_div/SumTmp[14][1] ), .S0(n117), .Y(n120) );
  MX2X1 U192 ( .A(n19), .B(\u_div/SumTmp[15][1] ), .S0(n201), .Y(n121) );
  MX2X1 U193 ( .A(n3), .B(\u_div/SumTmp[16][1] ), .S0(n202), .Y(n122) );
  MX2X1 U194 ( .A(n14), .B(\u_div/SumTmp[12][1] ), .S0(n227), .Y(n123) );
  MXI2X1 U195 ( .A(n182), .B(n193), .S0(quotient[1]), .Y(\u_div/PartRem[1][2] ) );
  INVX1 U196 ( .A(\u_div/SumTmp[1][1] ), .Y(n193) );
  INVX1 U197 ( .A(n180), .Y(\u_div/PartRem[2][3] ) );
  MXI2X1 U198 ( .A(n180), .B(n191), .S0(quotient[1]), .Y(\u_div/PartRem[1][4] ) );
  INVX1 U199 ( .A(\u_div/SumTmp[1][3] ), .Y(n191) );
  INVX1 U200 ( .A(n179), .Y(\u_div/PartRem[2][4] ) );
  INVX1 U201 ( .A(n178), .Y(\u_div/PartRem[2][5] ) );
  INVX1 U202 ( .A(n177), .Y(\u_div/PartRem[2][6] ) );
  MXI2X1 U203 ( .A(n178), .B(n189), .S0(quotient[1]), .Y(\u_div/PartRem[1][6] ) );
  INVX1 U204 ( .A(\u_div/SumTmp[1][5] ), .Y(n189) );
  INVX1 U205 ( .A(n176), .Y(\u_div/PartRem[2][7] ) );
  INVX1 U206 ( .A(n175), .Y(\u_div/PartRem[2][8] ) );
  MXI2X1 U207 ( .A(n176), .B(n187), .S0(quotient[1]), .Y(\u_div/PartRem[1][8] ) );
  INVX1 U208 ( .A(\u_div/SumTmp[1][7] ), .Y(n187) );
  INVX1 U209 ( .A(n174), .Y(\u_div/PartRem[2][9] ) );
  INVX1 U210 ( .A(n185), .Y(\u_div/PartRem[2][10] ) );
  MXI2X1 U211 ( .A(n174), .B(n196), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][10] ) );
  INVX1 U212 ( .A(\u_div/SumTmp[1][9] ), .Y(n196) );
  MXI2X1 U213 ( .A(n156), .B(\u_div/SumTmp[2][3] ), .S0(quotient[2]), .Y(n179)
         );
  MX2X1 U214 ( .A(n149), .B(\u_div/SumTmp[9][2] ), .S0(quotient[9]), .Y(n124)
         );
  MX2X1 U215 ( .A(n144), .B(\u_div/SumTmp[8][2] ), .S0(quotient[8]), .Y(n125)
         );
  MX2X1 U216 ( .A(n145), .B(\u_div/SumTmp[7][2] ), .S0(quotient[7]), .Y(n126)
         );
  MX2X1 U217 ( .A(n146), .B(\u_div/SumTmp[6][2] ), .S0(quotient[6]), .Y(n127)
         );
  MX2X1 U218 ( .A(n147), .B(\u_div/SumTmp[5][2] ), .S0(quotient[5]), .Y(n128)
         );
  MX2X1 U219 ( .A(n128), .B(\u_div/SumTmp[4][3] ), .S0(quotient[4]), .Y(n129)
         );
  MX2X1 U220 ( .A(n155), .B(\u_div/SumTmp[3][3] ), .S0(quotient[3]), .Y(n130)
         );
  MX2X1 U221 ( .A(n118), .B(\u_div/SumTmp[10][2] ), .S0(\u_div/CryTmp[10][12] ), .Y(n131) );
  MX2X1 U222 ( .A(n151), .B(\u_div/SumTmp[16][2] ), .S0(n202), .Y(n132) );
  MX2X1 U223 ( .A(n152), .B(\u_div/SumTmp[17][2] ), .S0(n203), .Y(n133) );
  MX2X1 U224 ( .A(n153), .B(\u_div/SumTmp[18][2] ), .S0(n204), .Y(n134) );
  MX2X1 U225 ( .A(n154), .B(\u_div/SumTmp[19][2] ), .S0(n206), .Y(n135) );
  MX2X1 U226 ( .A(n119), .B(\u_div/SumTmp[12][2] ), .S0(n227), .Y(n136) );
  MX2X1 U227 ( .A(n48), .B(\u_div/SumTmp[12][3] ), .S0(n227), .Y(n137) );
  MX2X1 U228 ( .A(n49), .B(\u_div/SumTmp[12][4] ), .S0(n227), .Y(n138) );
  MX2X1 U229 ( .A(n50), .B(\u_div/SumTmp[12][5] ), .S0(n227), .Y(n139) );
  MX2X1 U230 ( .A(n89), .B(\u_div/SumTmp[12][6] ), .S0(n227), .Y(n140) );
  MX2X1 U231 ( .A(n90), .B(\u_div/SumTmp[12][7] ), .S0(n227), .Y(n141) );
  MX2X1 U232 ( .A(n91), .B(\u_div/SumTmp[12][8] ), .S0(n227), .Y(n142) );
  MX2X1 U233 ( .A(n115), .B(\u_div/SumTmp[12][9] ), .S0(n227), .Y(n143) );
  INVX4 U234 ( .A(n226), .Y(\u_div/BInv [1]) );
  CLKINVX3 U235 ( .A(b[11]), .Y(\u_div/BInv [11]) );
  NAND2BX1 U236 ( .AN(n221), .B(n224), .Y(n209) );
  NOR2X1 U237 ( .A(b[4]), .B(b[3]), .Y(n224) );
  NAND2BX1 U238 ( .AN(n218), .B(n225), .Y(n221) );
  NOR2X1 U239 ( .A(b[6]), .B(b[5]), .Y(n225) );
  XNOR2X1 U240 ( .A(\u_div/CryTmp[2][1] ), .B(a[12]), .Y(\u_div/SumTmp[12][0] ) );
  INVX1 U241 ( .A(n212), .Y(n207) );
  NAND3BX1 U242 ( .AN(n209), .B(\u_div/BInv [2]), .C(\u_div/CryTmp[20][2] ), 
        .Y(n212) );
  MX2X1 U243 ( .A(n15), .B(\u_div/SumTmp[9][1] ), .S0(quotient[9]), .Y(n144)
         );
  MX2X1 U244 ( .A(n7), .B(\u_div/SumTmp[8][1] ), .S0(quotient[8]), .Y(n145) );
  MX2X1 U245 ( .A(n8), .B(\u_div/SumTmp[7][1] ), .S0(quotient[7]), .Y(n146) );
  MX2X1 U246 ( .A(n9), .B(\u_div/SumTmp[6][1] ), .S0(quotient[6]), .Y(n147) );
  MX2X1 U247 ( .A(n10), .B(\u_div/SumTmp[5][1] ), .S0(quotient[5]), .Y(n148)
         );
  MX2X1 U248 ( .A(n6), .B(\u_div/SumTmp[10][1] ), .S0(\u_div/CryTmp[10][12] ), 
        .Y(n149) );
  XNOR2X1 U249 ( .A(\u_div/CryTmp[2][1] ), .B(a[11]), .Y(\u_div/SumTmp[11][0] ) );
  XNOR2X1 U250 ( .A(\u_div/CryTmp[2][1] ), .B(a[13]), .Y(\u_div/SumTmp[13][0] ) );
  NOR2X1 U251 ( .A(b[8]), .B(n216), .Y(n150) );
  XNOR2X1 U252 ( .A(\u_div/CryTmp[2][1] ), .B(a[14]), .Y(\u_div/SumTmp[14][0] ) );
  XNOR2X1 U253 ( .A(\u_div/CryTmp[2][1] ), .B(a[15]), .Y(\u_div/SumTmp[15][0] ) );
  XNOR2X1 U254 ( .A(\u_div/CryTmp[2][1] ), .B(a[16]), .Y(\u_div/SumTmp[16][0] ) );
  XNOR2X1 U255 ( .A(\u_div/CryTmp[2][1] ), .B(a[17]), .Y(\u_div/SumTmp[17][0] ) );
  MX2X1 U256 ( .A(n5), .B(\u_div/SumTmp[17][1] ), .S0(n203), .Y(n151) );
  MX2X1 U257 ( .A(n13), .B(\u_div/SumTmp[18][1] ), .S0(n204), .Y(n152) );
  MX2X1 U258 ( .A(n18), .B(\u_div/SumTmp[19][1] ), .S0(n206), .Y(n153) );
  MX2X1 U259 ( .A(n17), .B(\u_div/SumTmp[20][1] ), .S0(n207), .Y(n154) );
  OR3XL U260 ( .A(b[9]), .B(b[10]), .C(b[11]), .Y(n216) );
  BUFX3 U261 ( .A(n199), .Y(n227) );
  NOR3X1 U262 ( .A(n214), .B(b[11]), .C(b[10]), .Y(n199) );
  INVX1 U263 ( .A(\u_div/CryTmp[12][10] ), .Y(n214) );
  OR2X2 U264 ( .A(a[17]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[17][1] )
         );
  OR2X2 U265 ( .A(a[16]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[16][1] )
         );
  OR2X2 U266 ( .A(a[15]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[15][1] )
         );
  OR2X2 U267 ( .A(a[14]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[14][1] )
         );
  OR2X2 U268 ( .A(a[13]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[13][1] )
         );
  OR2X2 U269 ( .A(a[11]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[11][1] )
         );
  OR2X2 U270 ( .A(a[12]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[12][1] )
         );
  INVX1 U271 ( .A(n181), .Y(\u_div/PartRem[2][2] ) );
  MXI2X1 U272 ( .A(n158), .B(\u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(n180)
         );
  MXI2X1 U273 ( .A(n181), .B(n192), .S0(quotient[1]), .Y(\u_div/PartRem[1][3] ) );
  INVX1 U274 ( .A(\u_div/SumTmp[1][2] ), .Y(n192) );
  MX2X1 U275 ( .A(n148), .B(\u_div/SumTmp[4][2] ), .S0(quotient[4]), .Y(n155)
         );
  MX2X1 U276 ( .A(n157), .B(\u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(n156)
         );
  BUFX3 U277 ( .A(b[1]), .Y(n226) );
  CLKINVX3 U278 ( .A(b[10]), .Y(\u_div/BInv [10]) );
  MXI2X1 U279 ( .A(n1), .B(\u_div/SumTmp[2][1] ), .S0(quotient[2]), .Y(n181)
         );
  XNOR2X1 U280 ( .A(\u_div/CryTmp[2][1] ), .B(a[9]), .Y(\u_div/SumTmp[9][0] )
         );
  XNOR2X1 U281 ( .A(\u_div/CryTmp[2][1] ), .B(a[8]), .Y(\u_div/SumTmp[8][0] )
         );
  XNOR2X1 U282 ( .A(\u_div/CryTmp[2][1] ), .B(a[7]), .Y(\u_div/SumTmp[7][0] )
         );
  XNOR2X1 U283 ( .A(\u_div/CryTmp[2][1] ), .B(a[6]), .Y(\u_div/SumTmp[6][0] )
         );
  XNOR2X1 U284 ( .A(\u_div/CryTmp[2][1] ), .B(a[5]), .Y(\u_div/SumTmp[5][0] )
         );
  MX2X1 U285 ( .A(n11), .B(\u_div/SumTmp[4][1] ), .S0(quotient[4]), .Y(n157)
         );
  MX2X1 U286 ( .A(n2), .B(\u_div/SumTmp[3][1] ), .S0(quotient[3]), .Y(n158) );
  XNOR2X1 U287 ( .A(\u_div/CryTmp[2][1] ), .B(a[10]), .Y(\u_div/SumTmp[10][0] ) );
  XNOR2X1 U288 ( .A(\u_div/CryTmp[2][1] ), .B(a[21]), .Y(\u_div/SumTmp[21][0] ) );
  NOR2X1 U289 ( .A(n209), .B(n210), .Y(n208) );
  XNOR2X1 U290 ( .A(\u_div/CryTmp[2][1] ), .B(a[20]), .Y(\u_div/SumTmp[20][0] ) );
  XNOR2X1 U291 ( .A(\u_div/CryTmp[2][1] ), .B(a[19]), .Y(\u_div/SumTmp[19][0] ) );
  XNOR2X1 U292 ( .A(\u_div/CryTmp[2][1] ), .B(a[18]), .Y(\u_div/SumTmp[18][0] ) );
  OR2XL U293 ( .A(a[20]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[20][1] )
         );
  OR2XL U294 ( .A(a[19]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[19][1] )
         );
  OR2XL U295 ( .A(a[18]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[18][1] )
         );
  OR2XL U296 ( .A(a[10]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[10][1] )
         );
  OR2XL U297 ( .A(a[9]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[9][1] ) );
  OR2XL U298 ( .A(a[8]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[8][1] ) );
  OR2XL U299 ( .A(a[7]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[7][1] ) );
  OR2XL U300 ( .A(a[6]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[6][1] ) );
  OR2XL U301 ( .A(a[5]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[5][1] ) );
  NAND2X1 U302 ( .A(\u_div/CryTmp[21][1] ), .B(n211), .Y(n210) );
  NOR2X1 U303 ( .A(b[2]), .B(n226), .Y(n211) );
  OR2XL U304 ( .A(a[21]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[21][1] )
         );
  XNOR2X1 U305 ( .A(\u_div/CryTmp[2][1] ), .B(a[3]), .Y(\u_div/SumTmp[3][0] )
         );
  OR2XL U306 ( .A(a[4]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[4][1] ) );
  OR2XL U307 ( .A(a[3]), .B(\u_div/CryTmp[2][1] ), .Y(\u_div/CryTmp[3][1] ) );
  NAND2BX4 U308 ( .AN(\u_div/CryTmp[9][12] ), .B(n29), .Y(quotient[9]) );
  NAND2BX4 U309 ( .AN(\u_div/CryTmp[8][12] ), .B(n22), .Y(quotient[8]) );
  NAND2BX4 U310 ( .AN(\u_div/CryTmp[7][12] ), .B(n23), .Y(quotient[7]) );
  NAND2BX4 U311 ( .AN(\u_div/CryTmp[6][12] ), .B(n24), .Y(quotient[6]) );
  NAND2BX4 U312 ( .AN(\u_div/CryTmp[5][12] ), .B(n25), .Y(quotient[5]) );
  NAND2BX4 U313 ( .AN(\u_div/CryTmp[4][12] ), .B(n26), .Y(quotient[4]) );
  NAND2BX4 U314 ( .AN(\u_div/CryTmp[3][12] ), .B(n28), .Y(quotient[3]) );
  NAND2BX4 U315 ( .AN(\u_div/CryTmp[2][12] ), .B(n27), .Y(quotient[2]) );
  NAND2BX4 U316 ( .AN(\u_div/CryTmp[1][12] ), .B(n21), .Y(quotient[1]) );
  CLKINVX8 U317 ( .A(b[0]), .Y(\u_div/CryTmp[2][1] ) );
endmodule


module Equation_Implementation_DW_div_uns_34 ( a, b, quotient, remainder, 
        divide_by_0 );
  input [22:0] a;
  input [11:0] b;
  output [22:0] quotient;
  output [11:0] remainder;
  output divide_by_0;
  wire   n242, \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] , \u_div/SumTmp[1][5] ,
         \u_div/SumTmp[1][6] , \u_div/SumTmp[1][7] , \u_div/SumTmp[1][8] ,
         \u_div/SumTmp[1][9] , \u_div/SumTmp[1][10] , \u_div/SumTmp[1][11] ,
         \u_div/SumTmp[2][1] , \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] ,
         \u_div/SumTmp[2][4] , \u_div/SumTmp[2][5] , \u_div/SumTmp[2][6] ,
         \u_div/SumTmp[2][7] , \u_div/SumTmp[2][8] , \u_div/SumTmp[2][9] ,
         \u_div/SumTmp[2][10] , \u_div/SumTmp[2][11] , \u_div/SumTmp[3][1] ,
         \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] , \u_div/SumTmp[3][4] ,
         \u_div/SumTmp[3][5] , \u_div/SumTmp[3][6] , \u_div/SumTmp[3][7] ,
         \u_div/SumTmp[3][8] , \u_div/SumTmp[3][9] , \u_div/SumTmp[3][10] ,
         \u_div/SumTmp[3][11] , \u_div/SumTmp[4][0] , \u_div/SumTmp[4][1] ,
         \u_div/SumTmp[4][2] , \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] ,
         \u_div/SumTmp[4][5] , \u_div/SumTmp[4][6] , \u_div/SumTmp[4][7] ,
         \u_div/SumTmp[4][8] , \u_div/SumTmp[4][9] , \u_div/SumTmp[4][10] ,
         \u_div/SumTmp[4][11] , \u_div/SumTmp[5][0] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[5][5] , \u_div/SumTmp[5][6] , \u_div/SumTmp[5][7] ,
         \u_div/SumTmp[5][8] , \u_div/SumTmp[5][9] , \u_div/SumTmp[5][10] ,
         \u_div/SumTmp[5][11] , \u_div/SumTmp[6][0] , \u_div/SumTmp[6][1] ,
         \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] , \u_div/SumTmp[6][4] ,
         \u_div/SumTmp[6][5] , \u_div/SumTmp[6][6] , \u_div/SumTmp[6][7] ,
         \u_div/SumTmp[6][8] , \u_div/SumTmp[6][9] , \u_div/SumTmp[6][10] ,
         \u_div/SumTmp[6][11] , \u_div/SumTmp[7][0] , \u_div/SumTmp[7][1] ,
         \u_div/SumTmp[7][2] , \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] ,
         \u_div/SumTmp[7][5] , \u_div/SumTmp[7][6] , \u_div/SumTmp[7][7] ,
         \u_div/SumTmp[7][8] , \u_div/SumTmp[7][9] , \u_div/SumTmp[7][10] ,
         \u_div/SumTmp[7][11] , \u_div/SumTmp[8][0] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[8][5] , \u_div/SumTmp[8][6] , \u_div/SumTmp[8][7] ,
         \u_div/SumTmp[8][8] , \u_div/SumTmp[8][9] , \u_div/SumTmp[8][10] ,
         \u_div/SumTmp[8][11] , \u_div/SumTmp[9][0] , \u_div/SumTmp[9][1] ,
         \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] , \u_div/SumTmp[9][4] ,
         \u_div/SumTmp[9][5] , \u_div/SumTmp[9][6] , \u_div/SumTmp[9][7] ,
         \u_div/SumTmp[9][8] , \u_div/SumTmp[9][9] , \u_div/SumTmp[9][10] ,
         \u_div/SumTmp[9][11] , \u_div/SumTmp[10][0] , \u_div/SumTmp[10][1] ,
         \u_div/SumTmp[10][2] , \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] ,
         \u_div/SumTmp[10][5] , \u_div/SumTmp[10][6] , \u_div/SumTmp[10][7] ,
         \u_div/SumTmp[10][8] , \u_div/SumTmp[10][9] , \u_div/SumTmp[10][10] ,
         \u_div/SumTmp[10][11] , \u_div/SumTmp[11][0] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[11][5] , \u_div/SumTmp[11][6] , \u_div/SumTmp[11][7] ,
         \u_div/SumTmp[11][8] , \u_div/SumTmp[11][9] , \u_div/SumTmp[11][10] ,
         \u_div/SumTmp[11][11] , \u_div/SumTmp[12][0] , \u_div/SumTmp[12][1] ,
         \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] , \u_div/SumTmp[12][4] ,
         \u_div/SumTmp[12][5] , \u_div/SumTmp[12][6] , \u_div/SumTmp[12][7] ,
         \u_div/SumTmp[12][8] , \u_div/SumTmp[12][9] , \u_div/SumTmp[12][10] ,
         \u_div/SumTmp[13][0] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[13][5] ,
         \u_div/SumTmp[13][6] , \u_div/SumTmp[13][7] , \u_div/SumTmp[13][8] ,
         \u_div/SumTmp[13][9] , \u_div/SumTmp[14][0] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[14][5] , \u_div/SumTmp[14][6] , \u_div/SumTmp[14][7] ,
         \u_div/SumTmp[14][8] , \u_div/SumTmp[15][0] , \u_div/SumTmp[15][1] ,
         \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] , \u_div/SumTmp[15][4] ,
         \u_div/SumTmp[15][5] , \u_div/SumTmp[15][6] , \u_div/SumTmp[15][7] ,
         \u_div/SumTmp[16][0] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] , \u_div/SumTmp[16][5] ,
         \u_div/SumTmp[16][6] , \u_div/SumTmp[17][0] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] ,
         \u_div/SumTmp[17][5] , \u_div/SumTmp[18][0] , \u_div/SumTmp[18][1] ,
         \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] , \u_div/SumTmp[18][4] ,
         \u_div/SumTmp[19][0] , \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] ,
         \u_div/SumTmp[19][3] , \u_div/SumTmp[20][0] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[21][0] , \u_div/SumTmp[21][1] ,
         \u_div/SumTmp[22][0] , \u_div/CryTmp[0][2] , \u_div/CryTmp[0][3] ,
         \u_div/CryTmp[0][4] , \u_div/CryTmp[0][5] , \u_div/CryTmp[0][6] ,
         \u_div/CryTmp[0][7] , \u_div/CryTmp[0][8] , \u_div/CryTmp[0][9] ,
         \u_div/CryTmp[0][10] , \u_div/CryTmp[0][11] , \u_div/CryTmp[0][12] ,
         \u_div/CryTmp[1][2] , \u_div/CryTmp[1][3] , \u_div/CryTmp[1][4] ,
         \u_div/CryTmp[1][5] , \u_div/CryTmp[1][6] , \u_div/CryTmp[1][7] ,
         \u_div/CryTmp[1][8] , \u_div/CryTmp[1][9] , \u_div/CryTmp[1][10] ,
         \u_div/CryTmp[1][11] , \u_div/CryTmp[1][12] , \u_div/CryTmp[2][2] ,
         \u_div/CryTmp[2][3] , \u_div/CryTmp[2][4] , \u_div/CryTmp[2][5] ,
         \u_div/CryTmp[2][6] , \u_div/CryTmp[2][7] , \u_div/CryTmp[2][8] ,
         \u_div/CryTmp[2][9] , \u_div/CryTmp[2][10] , \u_div/CryTmp[2][11] ,
         \u_div/CryTmp[2][12] , \u_div/CryTmp[3][1] , \u_div/CryTmp[3][2] ,
         \u_div/CryTmp[3][3] , \u_div/CryTmp[3][4] , \u_div/CryTmp[3][5] ,
         \u_div/CryTmp[3][6] , \u_div/CryTmp[3][7] , \u_div/CryTmp[3][8] ,
         \u_div/CryTmp[3][9] , \u_div/CryTmp[3][10] , \u_div/CryTmp[3][11] ,
         \u_div/CryTmp[3][12] , \u_div/CryTmp[4][1] , \u_div/CryTmp[4][2] ,
         \u_div/CryTmp[4][3] , \u_div/CryTmp[4][4] , \u_div/CryTmp[4][5] ,
         \u_div/CryTmp[4][6] , \u_div/CryTmp[4][7] , \u_div/CryTmp[4][8] ,
         \u_div/CryTmp[4][9] , \u_div/CryTmp[4][10] , \u_div/CryTmp[4][11] ,
         \u_div/CryTmp[4][12] , \u_div/CryTmp[5][1] , \u_div/CryTmp[5][2] ,
         \u_div/CryTmp[5][3] , \u_div/CryTmp[5][4] , \u_div/CryTmp[5][5] ,
         \u_div/CryTmp[5][6] , \u_div/CryTmp[5][7] , \u_div/CryTmp[5][8] ,
         \u_div/CryTmp[5][9] , \u_div/CryTmp[5][10] , \u_div/CryTmp[5][11] ,
         \u_div/CryTmp[5][12] , \u_div/CryTmp[6][1] , \u_div/CryTmp[6][2] ,
         \u_div/CryTmp[6][3] , \u_div/CryTmp[6][4] , \u_div/CryTmp[6][5] ,
         \u_div/CryTmp[6][6] , \u_div/CryTmp[6][7] , \u_div/CryTmp[6][8] ,
         \u_div/CryTmp[6][9] , \u_div/CryTmp[6][10] , \u_div/CryTmp[6][11] ,
         \u_div/CryTmp[6][12] , \u_div/CryTmp[7][1] , \u_div/CryTmp[7][2] ,
         \u_div/CryTmp[7][3] , \u_div/CryTmp[7][4] , \u_div/CryTmp[7][5] ,
         \u_div/CryTmp[7][6] , \u_div/CryTmp[7][7] , \u_div/CryTmp[7][8] ,
         \u_div/CryTmp[7][9] , \u_div/CryTmp[7][10] , \u_div/CryTmp[7][11] ,
         \u_div/CryTmp[7][12] , \u_div/CryTmp[8][1] , \u_div/CryTmp[8][2] ,
         \u_div/CryTmp[8][3] , \u_div/CryTmp[8][4] , \u_div/CryTmp[8][5] ,
         \u_div/CryTmp[8][6] , \u_div/CryTmp[8][7] , \u_div/CryTmp[8][8] ,
         \u_div/CryTmp[8][9] , \u_div/CryTmp[8][10] , \u_div/CryTmp[8][11] ,
         \u_div/CryTmp[8][12] , \u_div/CryTmp[9][1] , \u_div/CryTmp[9][2] ,
         \u_div/CryTmp[9][3] , \u_div/CryTmp[9][4] , \u_div/CryTmp[9][5] ,
         \u_div/CryTmp[9][6] , \u_div/CryTmp[9][7] , \u_div/CryTmp[9][8] ,
         \u_div/CryTmp[9][9] , \u_div/CryTmp[9][10] , \u_div/CryTmp[9][11] ,
         \u_div/CryTmp[9][12] , \u_div/CryTmp[10][1] , \u_div/CryTmp[10][2] ,
         \u_div/CryTmp[10][3] , \u_div/CryTmp[10][4] , \u_div/CryTmp[10][5] ,
         \u_div/CryTmp[10][6] , \u_div/CryTmp[10][7] , \u_div/CryTmp[10][8] ,
         \u_div/CryTmp[10][9] , \u_div/CryTmp[10][10] , \u_div/CryTmp[10][11] ,
         \u_div/CryTmp[10][12] , \u_div/CryTmp[11][1] , \u_div/CryTmp[11][2] ,
         \u_div/CryTmp[11][3] , \u_div/CryTmp[11][4] , \u_div/CryTmp[11][5] ,
         \u_div/CryTmp[11][6] , \u_div/CryTmp[11][7] , \u_div/CryTmp[11][8] ,
         \u_div/CryTmp[11][9] , \u_div/CryTmp[11][10] , \u_div/CryTmp[11][11] ,
         \u_div/CryTmp[11][12] , \u_div/CryTmp[12][1] , \u_div/CryTmp[12][2] ,
         \u_div/CryTmp[12][3] , \u_div/CryTmp[12][4] , \u_div/CryTmp[12][5] ,
         \u_div/CryTmp[12][6] , \u_div/CryTmp[12][7] , \u_div/CryTmp[12][8] ,
         \u_div/CryTmp[12][9] , \u_div/CryTmp[12][10] , \u_div/CryTmp[12][11] ,
         \u_div/CryTmp[13][1] , \u_div/CryTmp[13][2] , \u_div/CryTmp[13][3] ,
         \u_div/CryTmp[13][4] , \u_div/CryTmp[13][5] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[13][7] , \u_div/CryTmp[13][8] , \u_div/CryTmp[13][9] ,
         \u_div/CryTmp[13][10] , \u_div/CryTmp[14][1] , \u_div/CryTmp[14][2] ,
         \u_div/CryTmp[14][3] , \u_div/CryTmp[14][4] , \u_div/CryTmp[14][5] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[14][7] , \u_div/CryTmp[14][8] ,
         \u_div/CryTmp[14][9] , \u_div/CryTmp[15][1] , \u_div/CryTmp[15][2] ,
         \u_div/CryTmp[15][3] , \u_div/CryTmp[15][4] , \u_div/CryTmp[15][5] ,
         \u_div/CryTmp[15][6] , \u_div/CryTmp[15][7] , \u_div/CryTmp[15][8] ,
         \u_div/CryTmp[16][1] , \u_div/CryTmp[16][2] , \u_div/CryTmp[16][3] ,
         \u_div/CryTmp[16][4] , \u_div/CryTmp[16][5] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[16][7] , \u_div/CryTmp[17][1] , \u_div/CryTmp[17][2] ,
         \u_div/CryTmp[17][3] , \u_div/CryTmp[17][4] , \u_div/CryTmp[17][5] ,
         \u_div/CryTmp[17][6] , \u_div/CryTmp[18][1] , \u_div/CryTmp[18][2] ,
         \u_div/CryTmp[18][3] , \u_div/CryTmp[18][4] , \u_div/CryTmp[18][5] ,
         \u_div/CryTmp[19][1] , \u_div/CryTmp[19][2] , \u_div/CryTmp[19][3] ,
         \u_div/CryTmp[19][4] , \u_div/CryTmp[20][1] , \u_div/CryTmp[20][2] ,
         \u_div/CryTmp[20][3] , \u_div/CryTmp[21][1] , \u_div/CryTmp[21][2] ,
         \u_div/CryTmp[22][1] , \u_div/PartRem[1][2] , \u_div/PartRem[1][3] ,
         \u_div/PartRem[1][4] , \u_div/PartRem[1][5] , \u_div/PartRem[1][6] ,
         \u_div/PartRem[1][7] , \u_div/PartRem[1][8] , \u_div/PartRem[1][9] ,
         \u_div/PartRem[1][10] , \u_div/PartRem[1][11] , \u_div/PartRem[2][1] ,
         \u_div/PartRem[2][2] , \u_div/PartRem[2][3] , \u_div/PartRem[2][4] ,
         \u_div/PartRem[2][5] , \u_div/PartRem[2][6] , \u_div/PartRem[2][7] ,
         \u_div/PartRem[2][8] , \u_div/PartRem[2][9] , \u_div/PartRem[2][10] ,
         \u_div/PartRem[2][11] , \u_div/PartRem[3][11] ,
         \u_div/PartRem[4][11] , \u_div/PartRem[5][11] ,
         \u_div/PartRem[6][11] , \u_div/PartRem[7][11] ,
         \u_div/PartRem[8][11] , \u_div/PartRem[9][11] ,
         \u_div/PartRem[10][11] , \u_div/PartRem[11][11] ,
         \u_div/PartRem[12][11] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241;
  wire   [11:0] \u_div/BInv ;

  ADDFX2 \u_div/u_fa_PartRem_0_4_1  ( .A(n10), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[4][1] ), .CO(\u_div/CryTmp[4][2] ), .S(
        \u_div/SumTmp[4][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_1  ( .A(n9), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[5][1] ), .CO(\u_div/CryTmp[5][2] ), .S(
        \u_div/SumTmp[5][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_2  ( .A(n167), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[4][2] ), .CO(\u_div/CryTmp[4][3] ), .S(
        \u_div/SumTmp[4][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_2  ( .A(n157), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[5][2] ), .CO(\u_div/CryTmp[5][3] ), .S(
        \u_div/SumTmp[5][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_1  ( .A(n8), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[6][1] ), .CO(\u_div/CryTmp[6][2] ), .S(
        \u_div/SumTmp[6][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_1  ( .A(n7), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[7][1] ), .CO(\u_div/CryTmp[7][2] ), .S(
        \u_div/SumTmp[7][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_1  ( .A(n6), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[8][1] ), .CO(\u_div/CryTmp[8][2] ), .S(
        \u_div/SumTmp[8][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_1  ( .A(n12), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[9][1] ), .CO(\u_div/CryTmp[9][2] ), .S(
        \u_div/SumTmp[9][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_1  ( .A(n4), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[11][2] ), .S(
        \u_div/SumTmp[11][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_1  ( .A(n14), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[10][1] ), .CO(\u_div/CryTmp[10][2] ), .S(
        \u_div/SumTmp[10][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_1  ( .A(n19), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[19][1] ), .CO(\u_div/CryTmp[19][2] ), .S(
        \u_div/SumTmp[19][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_1  ( .A(n17), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[20][1] ), .CO(\u_div/CryTmp[20][2] ), .S(
        \u_div/SumTmp[20][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_21_1  ( .A(n16), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[21][1] ), .CO(\u_div/CryTmp[21][2] ), .S(
        \u_div/SumTmp[21][1] ) );
  CMPR32X1 \u_div/u_fa_PartRem_0_3_1  ( .A(n5), .B(\u_div/BInv [1]), .C(
        \u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[3][2] ), .S(
        \u_div/SumTmp[3][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_3  ( .A(n165), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[4][3] ), .CO(\u_div/CryTmp[4][4] ), .S(
        \u_div/SumTmp[4][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_3  ( .A(n136), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[5][3] ), .CO(\u_div/CryTmp[5][4] ), .S(
        \u_div/SumTmp[5][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_2  ( .A(n169), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[2][2] ), .CO(\u_div/CryTmp[2][3] ), .S(
        \u_div/SumTmp[2][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_2  ( .A(n168), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[3][2] ), .CO(\u_div/CryTmp[3][3] ), .S(
        \u_div/SumTmp[3][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_2  ( .A(n156), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[6][2] ), .CO(\u_div/CryTmp[6][3] ), .S(
        \u_div/SumTmp[6][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_2  ( .A(n155), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[7][2] ), .CO(\u_div/CryTmp[7][3] ), .S(
        \u_div/SumTmp[7][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_2  ( .A(n154), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[8][2] ), .CO(\u_div/CryTmp[8][3] ), .S(
        \u_div/SumTmp[8][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_2  ( .A(n126), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[11][2] ), .CO(\u_div/CryTmp[11][3] ), .S(
        \u_div/SumTmp[11][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_2  ( .A(n160), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[10][2] ), .CO(\u_div/CryTmp[10][3] ), .S(
        \u_div/SumTmp[10][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_2  ( .A(n159), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[9][2] ), .CO(\u_div/CryTmp[9][3] ), .S(
        \u_div/SumTmp[9][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_2  ( .A(n163), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[19][2] ), .CO(\u_div/CryTmp[19][3] ), .S(
        \u_div/SumTmp[19][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_1  ( .A(n13), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[13][1] ), .CO(\u_div/CryTmp[13][2] ), .S(
        \u_div/SumTmp[13][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_1  ( .A(n11), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[12][1] ), .CO(\u_div/CryTmp[12][2] ), .S(
        \u_div/SumTmp[12][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_1  ( .A(n2), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[14][1] ), .CO(\u_div/CryTmp[14][2] ), .S(
        \u_div/SumTmp[14][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_1  ( .A(n15), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[15][1] ), .CO(\u_div/CryTmp[15][2] ), .S(
        \u_div/SumTmp[15][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_1  ( .A(n18), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[16][1] ), .CO(\u_div/CryTmp[16][2] ), .S(
        \u_div/SumTmp[16][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_1  ( .A(n1), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[17][1] ), .CO(\u_div/CryTmp[17][2] ), .S(
        \u_div/SumTmp[17][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_1  ( .A(n3), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[18][1] ), .CO(\u_div/CryTmp[18][2] ), .S(
        \u_div/SumTmp[18][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_20_2  ( .A(n164), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[20][2] ), .CO(\u_div/CryTmp[20][3] ), .S(
        \u_div/SumTmp[20][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_9  ( .A(\u_div/PartRem[1][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[0][9] ), .CO(\u_div/CryTmp[0][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_10  ( .A(\u_div/PartRem[1][10] ), .B(
        \u_div/BInv [10]), .CI(\u_div/CryTmp[0][10] ), .CO(
        \u_div/CryTmp[0][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_10  ( .A(n123), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[10][10] ), .CO(\u_div/CryTmp[10][11] ), .S(
        \u_div/SumTmp[10][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_10  ( .A(n122), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[9][10] ), .CO(\u_div/CryTmp[9][11] ), .S(
        \u_div/SumTmp[9][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_10  ( .A(n120), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[8][10] ), .CO(\u_div/CryTmp[8][11] ), .S(
        \u_div/SumTmp[8][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_10  ( .A(n119), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[7][10] ), .CO(\u_div/CryTmp[7][11] ), .S(
        \u_div/SumTmp[7][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_10  ( .A(n118), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[6][10] ), .CO(\u_div/CryTmp[6][11] ), .S(
        \u_div/SumTmp[6][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_10  ( .A(n117), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[5][10] ), .CO(\u_div/CryTmp[5][11] ), .S(
        \u_div/SumTmp[5][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_10  ( .A(n116), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[4][10] ), .CO(\u_div/CryTmp[4][11] ), .S(
        \u_div/SumTmp[4][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_10  ( .A(n115), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[3][10] ), .CO(\u_div/CryTmp[3][11] ), .S(
        \u_div/SumTmp[3][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_10  ( .A(n121), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[2][10] ), .CO(\u_div/CryTmp[2][11] ), .S(
        \u_div/SumTmp[2][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_10  ( .A(\u_div/PartRem[2][10] ), .B(
        \u_div/BInv [10]), .CI(\u_div/CryTmp[1][10] ), .CO(
        \u_div/CryTmp[1][11] ), .S(\u_div/SumTmp[1][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_10  ( .A(n124), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[11][10] ), .CO(\u_div/CryTmp[11][11] ), .S(
        \u_div/SumTmp[11][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_9  ( .A(\u_div/PartRem[2][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[1][9] ), .CO(\u_div/CryTmp[1][10] ), .S(\u_div/SumTmp[1][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_9  ( .A(n103), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[11][9] ), .CO(\u_div/CryTmp[11][10] ), .S(
        \u_div/SumTmp[11][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_9  ( .A(n100), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[10][9] ), .CO(\u_div/CryTmp[10][10] ), .S(
        \u_div/SumTmp[10][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_9  ( .A(n97), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[9][9] ), .CO(\u_div/CryTmp[9][10] ), .S(
        \u_div/SumTmp[9][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_9  ( .A(n91), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[8][9] ), .CO(\u_div/CryTmp[8][10] ), .S(
        \u_div/SumTmp[8][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_9  ( .A(n90), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[7][9] ), .CO(\u_div/CryTmp[7][10] ), .S(
        \u_div/SumTmp[7][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_9  ( .A(n89), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[6][9] ), .CO(\u_div/CryTmp[6][10] ), .S(
        \u_div/SumTmp[6][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_9  ( .A(n88), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[5][9] ), .CO(\u_div/CryTmp[5][10] ), .S(
        \u_div/SumTmp[5][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_9  ( .A(n87), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[4][9] ), .CO(\u_div/CryTmp[4][10] ), .S(
        \u_div/SumTmp[4][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_9  ( .A(n114), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[3][9] ), .CO(\u_div/CryTmp[3][10] ), .S(
        \u_div/SumTmp[3][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_9  ( .A(n94), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[2][9] ), .CO(\u_div/CryTmp[2][10] ), .S(
        \u_div/SumTmp[2][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_9  ( .A(n151), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[12][9] ), .CO(\u_div/CryTmp[12][10] ), .S(
        \u_div/SumTmp[12][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_8  ( .A(\u_div/PartRem[2][8] ), .B(
        \u_div/BInv [8]), .CI(\u_div/CryTmp[1][8] ), .CO(\u_div/CryTmp[1][9] ), 
        .S(\u_div/SumTmp[1][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_8  ( .A(n93), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[2][8] ), .CO(\u_div/CryTmp[2][9] ), .S(
        \u_div/SumTmp[2][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_8  ( .A(n102), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[11][8] ), .CO(\u_div/CryTmp[11][9] ), .S(
        \u_div/SumTmp[11][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_8  ( .A(n99), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[10][8] ), .CO(\u_div/CryTmp[10][9] ), .S(
        \u_div/SumTmp[10][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_8  ( .A(n96), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[9][8] ), .CO(\u_div/CryTmp[9][9] ), .S(
        \u_div/SumTmp[9][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_8  ( .A(n86), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[8][8] ), .CO(\u_div/CryTmp[8][9] ), .S(
        \u_div/SumTmp[8][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_8  ( .A(n85), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[7][8] ), .CO(\u_div/CryTmp[7][9] ), .S(
        \u_div/SumTmp[7][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_8  ( .A(n84), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[6][8] ), .CO(\u_div/CryTmp[6][9] ), .S(
        \u_div/SumTmp[6][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_8  ( .A(n83), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[5][8] ), .CO(\u_div/CryTmp[5][9] ), .S(
        \u_div/SumTmp[5][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_8  ( .A(n82), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[4][8] ), .CO(\u_div/CryTmp[4][9] ), .S(
        \u_div/SumTmp[4][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_8  ( .A(n81), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[3][8] ), .CO(\u_div/CryTmp[3][9] ), .S(
        \u_div/SumTmp[3][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_8  ( .A(n150), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[12][8] ), .CO(\u_div/CryTmp[12][9] ), .S(
        \u_div/SumTmp[12][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_8  ( .A(n106), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[13][8] ), .CO(\u_div/CryTmp[13][9] ), .S(
        \u_div/SumTmp[13][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_7  ( .A(\u_div/PartRem[1][7] ), .B(
        \u_div/BInv [7]), .CI(\u_div/CryTmp[0][7] ), .CO(\u_div/CryTmp[0][8] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_8  ( .A(\u_div/PartRem[1][8] ), .B(
        \u_div/BInv [8]), .CI(\u_div/CryTmp[0][8] ), .CO(\u_div/CryTmp[0][9] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_7  ( .A(\u_div/PartRem[2][7] ), .B(
        \u_div/BInv [7]), .CI(\u_div/CryTmp[1][7] ), .CO(\u_div/CryTmp[1][8] ), 
        .S(\u_div/SumTmp[1][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_7  ( .A(n92), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[2][7] ), .CO(\u_div/CryTmp[2][8] ), .S(
        \u_div/SumTmp[2][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_7  ( .A(n80), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[3][7] ), .CO(\u_div/CryTmp[3][8] ), .S(
        \u_div/SumTmp[3][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_7  ( .A(n101), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[11][7] ), .CO(\u_div/CryTmp[11][8] ), .S(
        \u_div/SumTmp[11][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_7  ( .A(n98), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[10][7] ), .CO(\u_div/CryTmp[10][8] ), .S(
        \u_div/SumTmp[10][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_7  ( .A(n95), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[9][7] ), .CO(\u_div/CryTmp[9][8] ), .S(
        \u_div/SumTmp[9][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_7  ( .A(n78), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[8][7] ), .CO(\u_div/CryTmp[8][8] ), .S(
        \u_div/SumTmp[8][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_7  ( .A(n77), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[7][7] ), .CO(\u_div/CryTmp[7][8] ), .S(
        \u_div/SumTmp[7][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_7  ( .A(n76), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[6][7] ), .CO(\u_div/CryTmp[6][8] ), .S(
        \u_div/SumTmp[6][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_7  ( .A(n75), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[5][7] ), .CO(\u_div/CryTmp[5][8] ), .S(
        \u_div/SumTmp[5][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_7  ( .A(n74), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[4][7] ), .CO(\u_div/CryTmp[4][8] ), .S(
        \u_div/SumTmp[4][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_7  ( .A(n149), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[12][7] ), .CO(\u_div/CryTmp[12][8] ), .S(
        \u_div/SumTmp[12][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_7  ( .A(n105), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[13][7] ), .CO(\u_div/CryTmp[13][8] ), .S(
        \u_div/SumTmp[13][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_7  ( .A(n109), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[14][7] ), .CO(\u_div/CryTmp[14][8] ), .S(
        \u_div/SumTmp[14][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_6  ( .A(\u_div/PartRem[2][6] ), .B(
        \u_div/BInv [6]), .CI(\u_div/CryTmp[1][6] ), .CO(\u_div/CryTmp[1][7] ), 
        .S(\u_div/SumTmp[1][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_6  ( .A(n50), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[2][6] ), .CO(\u_div/CryTmp[2][7] ), .S(
        \u_div/SumTmp[2][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_6  ( .A(n79), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[3][6] ), .CO(\u_div/CryTmp[3][7] ), .S(
        \u_div/SumTmp[3][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_6  ( .A(n47), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[4][6] ), .CO(\u_div/CryTmp[4][7] ), .S(
        \u_div/SumTmp[4][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_6  ( .A(n60), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[11][6] ), .CO(\u_div/CryTmp[11][7] ), .S(
        \u_div/SumTmp[11][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_6  ( .A(n56), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[10][6] ), .CO(\u_div/CryTmp[10][7] ), .S(
        \u_div/SumTmp[10][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_6  ( .A(n53), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[9][6] ), .CO(\u_div/CryTmp[9][7] ), .S(
        \u_div/SumTmp[9][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_6  ( .A(n45), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[8][6] ), .CO(\u_div/CryTmp[8][7] ), .S(
        \u_div/SumTmp[8][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_6  ( .A(n44), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[7][6] ), .CO(\u_div/CryTmp[7][7] ), .S(
        \u_div/SumTmp[7][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_6  ( .A(n43), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[6][6] ), .CO(\u_div/CryTmp[6][7] ), .S(
        \u_div/SumTmp[6][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_6  ( .A(n42), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[5][6] ), .CO(\u_div/CryTmp[5][7] ), .S(
        \u_div/SumTmp[5][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_6  ( .A(n148), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[12][6] ), .CO(\u_div/CryTmp[12][7] ), .S(
        \u_div/SumTmp[12][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_6  ( .A(n104), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[13][6] ), .CO(\u_div/CryTmp[13][7] ), .S(
        \u_div/SumTmp[13][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_6  ( .A(n108), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[14][6] ), .CO(\u_div/CryTmp[14][7] ), .S(
        \u_div/SumTmp[14][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_6  ( .A(n111), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[15][6] ), .CO(\u_div/CryTmp[15][7] ), .S(
        \u_div/SumTmp[15][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_5  ( .A(\u_div/PartRem[1][5] ), .B(
        \u_div/BInv [5]), .CI(\u_div/CryTmp[0][5] ), .CO(\u_div/CryTmp[0][6] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_6  ( .A(\u_div/PartRem[1][6] ), .B(
        \u_div/BInv [6]), .CI(\u_div/CryTmp[0][6] ), .CO(\u_div/CryTmp[0][7] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_5  ( .A(\u_div/PartRem[2][5] ), .B(
        \u_div/BInv [5]), .CI(\u_div/CryTmp[1][5] ), .CO(\u_div/CryTmp[1][6] ), 
        .S(\u_div/SumTmp[1][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_5  ( .A(n49), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[2][5] ), .CO(\u_div/CryTmp[2][6] ), .S(
        \u_div/SumTmp[2][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_5  ( .A(n48), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[3][5] ), .CO(\u_div/CryTmp[3][6] ), .S(
        \u_div/SumTmp[3][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_5  ( .A(n46), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[4][5] ), .CO(\u_div/CryTmp[4][6] ), .S(
        \u_div/SumTmp[4][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_5  ( .A(n41), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[5][5] ), .CO(\u_div/CryTmp[5][6] ), .S(
        \u_div/SumTmp[5][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_5  ( .A(n59), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[11][5] ), .CO(\u_div/CryTmp[11][6] ), .S(
        \u_div/SumTmp[11][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_5  ( .A(n55), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[10][5] ), .CO(\u_div/CryTmp[10][6] ), .S(
        \u_div/SumTmp[10][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_5  ( .A(n52), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[9][5] ), .CO(\u_div/CryTmp[9][6] ), .S(
        \u_div/SumTmp[9][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_5  ( .A(n39), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[8][5] ), .CO(\u_div/CryTmp[8][6] ), .S(
        \u_div/SumTmp[8][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_5  ( .A(n38), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[7][5] ), .CO(\u_div/CryTmp[7][6] ), .S(
        \u_div/SumTmp[7][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_5  ( .A(n37), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[6][5] ), .CO(\u_div/CryTmp[6][6] ), .S(
        \u_div/SumTmp[6][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_5  ( .A(n147), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[12][5] ), .CO(\u_div/CryTmp[12][6] ), .S(
        \u_div/SumTmp[12][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_5  ( .A(n63), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[13][5] ), .CO(\u_div/CryTmp[13][6] ), .S(
        \u_div/SumTmp[13][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_5  ( .A(n66), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[14][5] ), .CO(\u_div/CryTmp[14][6] ), .S(
        \u_div/SumTmp[14][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_5  ( .A(n69), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[15][5] ), .CO(\u_div/CryTmp[15][6] ), .S(
        \u_div/SumTmp[15][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_5  ( .A(n71), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[16][5] ), .CO(\u_div/CryTmp[16][6] ), .S(
        \u_div/SumTmp[16][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/BInv [4]), .CI(\u_div/CryTmp[1][4] ), .CO(\u_div/CryTmp[1][5] ), 
        .S(\u_div/SumTmp[1][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_4  ( .A(n139), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[2][4] ), .CO(\u_div/CryTmp[2][5] ), .S(
        \u_div/SumTmp[2][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_4  ( .A(n138), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[3][4] ), .CO(\u_div/CryTmp[3][5] ), .S(
        \u_div/SumTmp[3][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_4  ( .A(n137), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[4][4] ), .CO(\u_div/CryTmp[4][5] ), .S(
        \u_div/SumTmp[4][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_4  ( .A(n40), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[5][4] ), .CO(\u_div/CryTmp[5][5] ), .S(
        \u_div/SumTmp[5][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_4  ( .A(n36), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[6][4] ), .CO(\u_div/CryTmp[6][5] ), .S(
        \u_div/SumTmp[6][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_4  ( .A(n146), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[12][4] ), .CO(\u_div/CryTmp[12][5] ), .S(
        \u_div/SumTmp[12][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_4  ( .A(n58), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[11][4] ), .CO(\u_div/CryTmp[11][5] ), .S(
        \u_div/SumTmp[11][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_4  ( .A(n54), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[10][4] ), .CO(\u_div/CryTmp[10][5] ), .S(
        \u_div/SumTmp[10][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_4  ( .A(n51), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[9][4] ), .CO(\u_div/CryTmp[9][5] ), .S(
        \u_div/SumTmp[9][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_4  ( .A(n35), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[8][4] ), .CO(\u_div/CryTmp[8][5] ), .S(
        \u_div/SumTmp[8][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_4  ( .A(n34), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[7][4] ), .CO(\u_div/CryTmp[7][5] ), .S(
        \u_div/SumTmp[7][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_4  ( .A(n62), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[13][4] ), .CO(\u_div/CryTmp[13][5] ), .S(
        \u_div/SumTmp[13][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_4  ( .A(n65), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[14][4] ), .CO(\u_div/CryTmp[14][5] ), .S(
        \u_div/SumTmp[14][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_4  ( .A(n68), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[15][4] ), .CO(\u_div/CryTmp[15][5] ), .S(
        \u_div/SumTmp[15][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_4  ( .A(n70), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[16][4] ), .CO(\u_div/CryTmp[16][5] ), .S(
        \u_div/SumTmp[16][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_4  ( .A(n72), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[17][4] ), .CO(\u_div/CryTmp[17][5] ), .S(
        \u_div/SumTmp[17][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_3  ( .A(\u_div/PartRem[1][3] ), .B(
        \u_div/BInv [3]), .CI(\u_div/CryTmp[0][3] ), .CO(\u_div/CryTmp[0][4] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_4  ( .A(\u_div/PartRem[1][4] ), .B(
        \u_div/BInv [4]), .CI(\u_div/CryTmp[0][4] ), .CO(\u_div/CryTmp[0][5] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/BInv [3]), .CI(\u_div/CryTmp[1][3] ), .CO(\u_div/CryTmp[1][4] ), 
        .S(\u_div/SumTmp[1][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_3  ( .A(n158), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[2][3] ), .CO(\u_div/CryTmp[2][4] ), .S(
        \u_div/SumTmp[2][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_3  ( .A(n166), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[3][3] ), .CO(\u_div/CryTmp[3][4] ), .S(
        \u_div/SumTmp[3][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_3  ( .A(n135), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[6][3] ), .CO(\u_div/CryTmp[6][4] ), .S(
        \u_div/SumTmp[6][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_3  ( .A(n134), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[7][3] ), .CO(\u_div/CryTmp[7][4] ), .S(
        \u_div/SumTmp[7][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_3  ( .A(n145), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[12][3] ), .CO(\u_div/CryTmp[12][4] ), .S(
        \u_div/SumTmp[12][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_3  ( .A(n57), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[11][3] ), .CO(\u_div/CryTmp[11][4] ), .S(
        \u_div/SumTmp[11][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_3  ( .A(n141), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[10][3] ), .CO(\u_div/CryTmp[10][4] ), .S(
        \u_div/SumTmp[10][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_3  ( .A(n140), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[9][3] ), .CO(\u_div/CryTmp[9][4] ), .S(
        \u_div/SumTmp[9][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_3  ( .A(n133), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[8][3] ), .CO(\u_div/CryTmp[8][4] ), .S(
        \u_div/SumTmp[8][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_3  ( .A(n61), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[13][3] ), .CO(\u_div/CryTmp[13][4] ), .S(
        \u_div/SumTmp[13][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_3  ( .A(n64), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[14][3] ), .CO(\u_div/CryTmp[14][4] ), .S(
        \u_div/SumTmp[14][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_3  ( .A(n67), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[15][3] ), .CO(\u_div/CryTmp[15][4] ), .S(
        \u_div/SumTmp[15][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_3  ( .A(n142), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[16][3] ), .CO(\u_div/CryTmp[16][4] ), .S(
        \u_div/SumTmp[16][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_3  ( .A(n143), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[17][3] ), .CO(\u_div/CryTmp[17][4] ), .S(
        \u_div/SumTmp[17][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_3  ( .A(n132), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[18][3] ), .CO(\u_div/CryTmp[18][4] ), .S(
        \u_div/SumTmp[18][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/BInv [2]), .CI(\u_div/CryTmp[1][2] ), .CO(\u_div/CryTmp[1][3] ), 
        .S(\u_div/SumTmp[1][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_2  ( .A(n131), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[12][2] ), .CO(\u_div/CryTmp[12][3] ), .S(
        \u_div/SumTmp[12][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_2  ( .A(n127), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[13][2] ), .CO(\u_div/CryTmp[13][3] ), .S(
        \u_div/SumTmp[13][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_2  ( .A(n128), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[14][2] ), .CO(\u_div/CryTmp[14][3] ), .S(
        \u_div/SumTmp[14][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_2  ( .A(n129), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[15][2] ), .CO(\u_div/CryTmp[15][3] ), .S(
        \u_div/SumTmp[15][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_2  ( .A(n130), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[16][2] ), .CO(\u_div/CryTmp[16][3] ), .S(
        \u_div/SumTmp[16][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_2  ( .A(n162), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[17][2] ), .CO(\u_div/CryTmp[17][3] ), .S(
        \u_div/SumTmp[17][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_2  ( .A(n153), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[18][2] ), .CO(\u_div/CryTmp[18][3] ), .S(
        \u_div/SumTmp[18][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_5  ( .A(n73), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[17][5] ), .CO(\u_div/CryTmp[17][6] ), .S(
        \u_div/SumTmp[17][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_19_3  ( .A(n144), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[19][3] ), .CO(\u_div/CryTmp[19][4] ), .S(
        \u_div/SumTmp[19][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_10  ( .A(n152), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[12][10] ), .CO(\u_div/CryTmp[12][11] ), .S(
        \u_div/SumTmp[12][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_8  ( .A(n110), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[14][8] ), .CO(\u_div/CryTmp[14][9] ), .S(
        \u_div/SumTmp[14][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_6  ( .A(n113), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[16][6] ), .CO(\u_div/CryTmp[16][7] ), .S(
        \u_div/SumTmp[16][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_7  ( .A(n112), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[15][7] ), .CO(\u_div/CryTmp[15][8] ), .S(
        \u_div/SumTmp[15][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_4  ( .A(n33), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[18][4] ), .CO(\u_div/CryTmp[18][5] ), .S(
        \u_div/SumTmp[18][4] ) );
  CMPR32X1 \u_div/u_fa_PartRem_0_0_1  ( .A(n32), .B(\u_div/BInv [1]), .C(
        \u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[0][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/BInv [2]), .CI(\u_div/CryTmp[0][2] ), .CO(\u_div/CryTmp[0][3] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_13_9  ( .A(n107), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[13][9] ), .CO(\u_div/CryTmp[13][10] ), .S(
        \u_div/SumTmp[13][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_11  ( .A(\u_div/PartRem[11][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[10][11] ), .CO(
        \u_div/CryTmp[10][12] ), .S(\u_div/SumTmp[10][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_11  ( .A(\u_div/PartRem[10][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[9][11] ), .CO(
        \u_div/CryTmp[9][12] ), .S(\u_div/SumTmp[9][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_11  ( .A(\u_div/PartRem[9][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[8][11] ), .CO(
        \u_div/CryTmp[8][12] ), .S(\u_div/SumTmp[8][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_11  ( .A(\u_div/PartRem[8][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[7][11] ), .CO(
        \u_div/CryTmp[7][12] ), .S(\u_div/SumTmp[7][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_11  ( .A(\u_div/PartRem[7][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[6][11] ), .CO(
        \u_div/CryTmp[6][12] ), .S(\u_div/SumTmp[6][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_11  ( .A(\u_div/PartRem[6][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[5][11] ), .CO(
        \u_div/CryTmp[5][12] ), .S(\u_div/SumTmp[5][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_11  ( .A(\u_div/PartRem[5][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[4][11] ), .CO(
        \u_div/CryTmp[4][12] ), .S(\u_div/SumTmp[4][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_11  ( .A(\u_div/PartRem[4][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[3][11] ), .CO(
        \u_div/CryTmp[3][12] ), .S(\u_div/SumTmp[3][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_11  ( .A(\u_div/PartRem[3][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[2][11] ), .CO(
        \u_div/CryTmp[2][12] ), .S(\u_div/SumTmp[2][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_11  ( .A(\u_div/PartRem[2][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[1][11] ), .CO(
        \u_div/CryTmp[1][12] ), .S(\u_div/SumTmp[1][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_11  ( .A(\u_div/PartRem[1][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[0][11] ), .CO(
        \u_div/CryTmp[0][12] ) );
  CMPR32X1 \u_div/u_fa_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        \u_div/BInv [1]), .C(\u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[1][2] ), 
        .S(\u_div/SumTmp[1][1] ) );
  CMPR32X1 \u_div/u_fa_PartRem_0_2_1  ( .A(n31), .B(\u_div/BInv [1]), .C(
        \u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[2][2] ), .S(
        \u_div/SumTmp[2][1] ) );
  ADDFX4 \u_div/u_fa_PartRem_0_11_11  ( .A(\u_div/PartRem[12][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[11][11] ), .CO(
        \u_div/CryTmp[11][12] ), .S(\u_div/SumTmp[11][11] ) );
  INVX1 U1 ( .A(n226), .Y(n217) );
  INVX4 U2 ( .A(b[4]), .Y(\u_div/BInv [4]) );
  INVX4 U3 ( .A(b[3]), .Y(\u_div/BInv [3]) );
  INVX4 U4 ( .A(b[6]), .Y(\u_div/BInv [6]) );
  INVX4 U5 ( .A(b[5]), .Y(\u_div/BInv [5]) );
  INVX4 U6 ( .A(b[7]), .Y(\u_div/BInv [7]) );
  MX2X1 U7 ( .A(a[18]), .B(\u_div/SumTmp[18][0] ), .S0(n215), .Y(n1) );
  MX2X1 U8 ( .A(a[15]), .B(\u_div/SumTmp[15][0] ), .S0(n125), .Y(n2) );
  MX2X1 U9 ( .A(a[19]), .B(\u_div/SumTmp[19][0] ), .S0(n216), .Y(n3) );
  MX2X1 U10 ( .A(a[12]), .B(\u_div/SumTmp[12][0] ), .S0(n210), .Y(n4) );
  MX2X1 U11 ( .A(a[4]), .B(\u_div/SumTmp[4][0] ), .S0(quotient[4]), .Y(n5) );
  MX2X1 U12 ( .A(a[9]), .B(\u_div/SumTmp[9][0] ), .S0(quotient[9]), .Y(n6) );
  MX2X1 U13 ( .A(a[8]), .B(\u_div/SumTmp[8][0] ), .S0(quotient[8]), .Y(n7) );
  MX2X1 U14 ( .A(a[7]), .B(\u_div/SumTmp[7][0] ), .S0(quotient[7]), .Y(n8) );
  MX2X1 U15 ( .A(a[6]), .B(\u_div/SumTmp[6][0] ), .S0(quotient[6]), .Y(n9) );
  MX2X1 U16 ( .A(a[5]), .B(\u_div/SumTmp[5][0] ), .S0(quotient[5]), .Y(n10) );
  MX2X1 U17 ( .A(a[13]), .B(\u_div/SumTmp[13][0] ), .S0(n241), .Y(n11) );
  MX2X1 U18 ( .A(a[10]), .B(\u_div/SumTmp[10][0] ), .S0(n242), .Y(n12) );
  MX2X1 U19 ( .A(a[14]), .B(\u_div/SumTmp[14][0] ), .S0(n212), .Y(n13) );
  MX2X1 U20 ( .A(a[11]), .B(\u_div/SumTmp[11][0] ), .S0(\u_div/CryTmp[11][12] ), .Y(n14) );
  MX2X1 U21 ( .A(a[16]), .B(\u_div/SumTmp[16][0] ), .S0(n213), .Y(n15) );
  MX2X1 U22 ( .A(a[22]), .B(\u_div/SumTmp[22][0] ), .S0(n219), .Y(n16) );
  MX2X1 U23 ( .A(a[21]), .B(\u_div/SumTmp[21][0] ), .S0(n218), .Y(n17) );
  MX2X1 U24 ( .A(a[17]), .B(\u_div/SumTmp[17][0] ), .S0(n214), .Y(n18) );
  MX2X1 U25 ( .A(a[20]), .B(\u_div/SumTmp[20][0] ), .S0(n217), .Y(n19) );
  MX2X1 U26 ( .A(n195), .B(n205), .S0(quotient[1]), .Y(n20) );
  MX2X1 U27 ( .A(n184), .B(n194), .S0(quotient[2]), .Y(n21) );
  MX2X1 U28 ( .A(n170), .B(n171), .S0(quotient[9]), .Y(n22) );
  MX2X1 U29 ( .A(n172), .B(n173), .S0(quotient[8]), .Y(n23) );
  MX2X1 U30 ( .A(n174), .B(n175), .S0(quotient[7]), .Y(n24) );
  MX2X1 U31 ( .A(n176), .B(n177), .S0(quotient[6]), .Y(n25) );
  MX2X1 U32 ( .A(n178), .B(n179), .S0(quotient[5]), .Y(n26) );
  MX2X1 U33 ( .A(n180), .B(n181), .S0(quotient[4]), .Y(n27) );
  MX2X1 U34 ( .A(n182), .B(n183), .S0(quotient[3]), .Y(n28) );
  MX2X1 U35 ( .A(n223), .B(n224), .S0(n242), .Y(n29) );
  MX2X1 U36 ( .A(n208), .B(n209), .S0(\u_div/CryTmp[11][12] ), .Y(n30) );
  CLKINVX3 U37 ( .A(b[8]), .Y(\u_div/BInv [8]) );
  CLKINVX3 U38 ( .A(b[9]), .Y(\u_div/BInv [9]) );
  CLKINVX3 U39 ( .A(b[10]), .Y(\u_div/BInv [10]) );
  INVX1 U40 ( .A(\u_div/SumTmp[5][11] ), .Y(n179) );
  INVX1 U41 ( .A(\u_div/SumTmp[6][11] ), .Y(n177) );
  INVX1 U42 ( .A(\u_div/SumTmp[7][11] ), .Y(n175) );
  INVX1 U43 ( .A(\u_div/SumTmp[8][11] ), .Y(n173) );
  INVX1 U44 ( .A(\u_div/SumTmp[9][11] ), .Y(n171) );
  INVX1 U45 ( .A(\u_div/SumTmp[10][11] ), .Y(n224) );
  INVX1 U46 ( .A(\u_div/SumTmp[2][11] ), .Y(n194) );
  INVX1 U47 ( .A(\u_div/SumTmp[3][11] ), .Y(n183) );
  INVX1 U48 ( .A(\u_div/SumTmp[4][11] ), .Y(n181) );
  INVX1 U49 ( .A(\u_div/SumTmp[11][11] ), .Y(n209) );
  MXI2X1 U50 ( .A(n31), .B(\u_div/SumTmp[2][1] ), .S0(quotient[2]), .Y(n192)
         );
  NAND2X1 U51 ( .A(quotient[2]), .B(b[0]), .Y(n193) );
  NOR2BX1 U52 ( .AN(quotient[3]), .B(\u_div/CryTmp[3][1] ), .Y(n31) );
  NOR2BX1 U53 ( .AN(quotient[1]), .B(\u_div/CryTmp[3][1] ), .Y(n32) );
  INVX1 U54 ( .A(\u_div/SumTmp[1][11] ), .Y(n205) );
  INVX1 U55 ( .A(n208), .Y(\u_div/PartRem[12][11] ) );
  CLKINVX3 U56 ( .A(n233), .Y(n213) );
  NAND2BX1 U57 ( .AN(n234), .B(\u_div/CryTmp[16][7] ), .Y(n233) );
  INVX1 U58 ( .A(n193), .Y(\u_div/PartRem[2][1] ) );
  NAND2BX1 U59 ( .AN(\u_div/CryTmp[0][12] ), .B(n20), .Y(quotient[0]) );
  INVX1 U60 ( .A(n195), .Y(\u_div/PartRem[2][11] ) );
  INVX1 U61 ( .A(n184), .Y(\u_div/PartRem[3][11] ) );
  INVX1 U62 ( .A(n182), .Y(\u_div/PartRem[4][11] ) );
  INVX1 U63 ( .A(n180), .Y(\u_div/PartRem[5][11] ) );
  INVX1 U64 ( .A(n178), .Y(\u_div/PartRem[6][11] ) );
  INVX1 U65 ( .A(n176), .Y(\u_div/PartRem[7][11] ) );
  INVX1 U66 ( .A(n174), .Y(\u_div/PartRem[8][11] ) );
  INVX1 U67 ( .A(n172), .Y(\u_div/PartRem[9][11] ) );
  INVX1 U68 ( .A(n170), .Y(\u_div/PartRem[10][11] ) );
  INVX1 U69 ( .A(n223), .Y(\u_div/PartRem[11][11] ) );
  MXI2X1 U70 ( .A(n139), .B(\u_div/SumTmp[2][4] ), .S0(quotient[2]), .Y(n189)
         );
  MXI2X1 U71 ( .A(n192), .B(n203), .S0(quotient[1]), .Y(\u_div/PartRem[1][3] )
         );
  INVX1 U72 ( .A(\u_div/SumTmp[1][2] ), .Y(n203) );
  MX2X1 U73 ( .A(n144), .B(\u_div/SumTmp[19][3] ), .S0(n216), .Y(n33) );
  MX2X1 U74 ( .A(n133), .B(\u_div/SumTmp[8][3] ), .S0(quotient[8]), .Y(n34) );
  MX2X1 U75 ( .A(n140), .B(\u_div/SumTmp[9][3] ), .S0(quotient[9]), .Y(n35) );
  MX2X1 U76 ( .A(n134), .B(\u_div/SumTmp[7][3] ), .S0(quotient[7]), .Y(n36) );
  MX2X1 U77 ( .A(n34), .B(\u_div/SumTmp[7][4] ), .S0(quotient[7]), .Y(n37) );
  MX2X1 U78 ( .A(n35), .B(\u_div/SumTmp[8][4] ), .S0(quotient[8]), .Y(n38) );
  MX2X1 U79 ( .A(n51), .B(\u_div/SumTmp[9][4] ), .S0(quotient[9]), .Y(n39) );
  MX2X1 U80 ( .A(n135), .B(\u_div/SumTmp[6][3] ), .S0(quotient[6]), .Y(n40) );
  MX2X1 U81 ( .A(n36), .B(\u_div/SumTmp[6][4] ), .S0(quotient[6]), .Y(n41) );
  MX2X1 U82 ( .A(n37), .B(\u_div/SumTmp[6][5] ), .S0(quotient[6]), .Y(n42) );
  MX2X1 U83 ( .A(n38), .B(\u_div/SumTmp[7][5] ), .S0(quotient[7]), .Y(n43) );
  MX2X1 U84 ( .A(n39), .B(\u_div/SumTmp[8][5] ), .S0(quotient[8]), .Y(n44) );
  MX2X1 U85 ( .A(n52), .B(\u_div/SumTmp[9][5] ), .S0(quotient[9]), .Y(n45) );
  MX2X1 U86 ( .A(n40), .B(\u_div/SumTmp[5][4] ), .S0(quotient[5]), .Y(n46) );
  MX2X1 U87 ( .A(n41), .B(\u_div/SumTmp[5][5] ), .S0(quotient[5]), .Y(n47) );
  MX2X1 U88 ( .A(n137), .B(\u_div/SumTmp[4][4] ), .S0(quotient[4]), .Y(n48) );
  MX2X1 U89 ( .A(n138), .B(\u_div/SumTmp[3][4] ), .S0(quotient[3]), .Y(n49) );
  MX2X1 U90 ( .A(n48), .B(\u_div/SumTmp[3][5] ), .S0(quotient[3]), .Y(n50) );
  MX2X1 U91 ( .A(n141), .B(\u_div/SumTmp[10][3] ), .S0(n242), .Y(n51) );
  MX2X1 U92 ( .A(n54), .B(\u_div/SumTmp[10][4] ), .S0(n242), .Y(n52) );
  MX2X1 U93 ( .A(n55), .B(\u_div/SumTmp[10][5] ), .S0(n242), .Y(n53) );
  MX2X1 U94 ( .A(n57), .B(\u_div/SumTmp[11][3] ), .S0(\u_div/CryTmp[11][12] ), 
        .Y(n54) );
  MX2X1 U95 ( .A(n58), .B(\u_div/SumTmp[11][4] ), .S0(\u_div/CryTmp[11][12] ), 
        .Y(n55) );
  MX2X1 U96 ( .A(n59), .B(\u_div/SumTmp[11][5] ), .S0(\u_div/CryTmp[11][12] ), 
        .Y(n56) );
  MX2X1 U97 ( .A(n131), .B(\u_div/SumTmp[12][2] ), .S0(n210), .Y(n57) );
  MX2X1 U98 ( .A(n145), .B(\u_div/SumTmp[12][3] ), .S0(n210), .Y(n58) );
  MX2X1 U99 ( .A(n146), .B(\u_div/SumTmp[12][4] ), .S0(n210), .Y(n59) );
  MX2X1 U100 ( .A(n147), .B(\u_div/SumTmp[12][5] ), .S0(n210), .Y(n60) );
  MX2X1 U101 ( .A(n128), .B(\u_div/SumTmp[14][2] ), .S0(n212), .Y(n61) );
  MX2X1 U102 ( .A(n64), .B(\u_div/SumTmp[14][3] ), .S0(n212), .Y(n62) );
  MX2X1 U103 ( .A(n65), .B(\u_div/SumTmp[14][4] ), .S0(n212), .Y(n63) );
  MX2X1 U104 ( .A(n129), .B(\u_div/SumTmp[15][2] ), .S0(n125), .Y(n64) );
  MX2X1 U105 ( .A(n67), .B(\u_div/SumTmp[15][3] ), .S0(n125), .Y(n65) );
  MX2X1 U106 ( .A(n68), .B(\u_div/SumTmp[15][4] ), .S0(n125), .Y(n66) );
  MX2X1 U107 ( .A(n130), .B(\u_div/SumTmp[16][2] ), .S0(n213), .Y(n67) );
  MX2X1 U108 ( .A(n142), .B(\u_div/SumTmp[16][3] ), .S0(n213), .Y(n68) );
  MX2X1 U109 ( .A(n70), .B(\u_div/SumTmp[16][4] ), .S0(n213), .Y(n69) );
  MX2X1 U110 ( .A(n143), .B(\u_div/SumTmp[17][3] ), .S0(n214), .Y(n70) );
  MX2X1 U111 ( .A(n72), .B(\u_div/SumTmp[17][4] ), .S0(n214), .Y(n71) );
  MX2X1 U112 ( .A(n132), .B(\u_div/SumTmp[18][3] ), .S0(n215), .Y(n72) );
  MX2X1 U113 ( .A(n33), .B(\u_div/SumTmp[18][4] ), .S0(n215), .Y(n73) );
  MXI2X1 U114 ( .A(n49), .B(\u_div/SumTmp[2][5] ), .S0(quotient[2]), .Y(n188)
         );
  MXI2X1 U115 ( .A(n92), .B(\u_div/SumTmp[2][7] ), .S0(quotient[2]), .Y(n186)
         );
  MXI2X1 U116 ( .A(n50), .B(\u_div/SumTmp[2][6] ), .S0(quotient[2]), .Y(n187)
         );
  MXI2X1 U117 ( .A(n190), .B(n201), .S0(quotient[1]), .Y(\u_div/PartRem[1][5] ) );
  INVX1 U118 ( .A(\u_div/SumTmp[1][4] ), .Y(n201) );
  MXI2X1 U119 ( .A(n188), .B(n199), .S0(quotient[1]), .Y(\u_div/PartRem[1][7] ) );
  INVX1 U120 ( .A(\u_div/SumTmp[1][6] ), .Y(n199) );
  MX2X1 U121 ( .A(n42), .B(\u_div/SumTmp[5][6] ), .S0(quotient[5]), .Y(n74) );
  MX2X1 U122 ( .A(n43), .B(\u_div/SumTmp[6][6] ), .S0(quotient[6]), .Y(n75) );
  MX2X1 U123 ( .A(n44), .B(\u_div/SumTmp[7][6] ), .S0(quotient[7]), .Y(n76) );
  MX2X1 U124 ( .A(n45), .B(\u_div/SumTmp[8][6] ), .S0(quotient[8]), .Y(n77) );
  MX2X1 U125 ( .A(n53), .B(\u_div/SumTmp[9][6] ), .S0(quotient[9]), .Y(n78) );
  MX2X1 U126 ( .A(n46), .B(\u_div/SumTmp[4][5] ), .S0(quotient[4]), .Y(n79) );
  MX2X1 U127 ( .A(n47), .B(\u_div/SumTmp[4][6] ), .S0(quotient[4]), .Y(n80) );
  MX2X1 U128 ( .A(n74), .B(\u_div/SumTmp[4][7] ), .S0(quotient[4]), .Y(n81) );
  MX2X1 U129 ( .A(n75), .B(\u_div/SumTmp[5][7] ), .S0(quotient[5]), .Y(n82) );
  MX2X1 U130 ( .A(n76), .B(\u_div/SumTmp[6][7] ), .S0(quotient[6]), .Y(n83) );
  MX2X1 U131 ( .A(n77), .B(\u_div/SumTmp[7][7] ), .S0(quotient[7]), .Y(n84) );
  MX2X1 U132 ( .A(n78), .B(\u_div/SumTmp[8][7] ), .S0(quotient[8]), .Y(n85) );
  MX2X1 U133 ( .A(n95), .B(\u_div/SumTmp[9][7] ), .S0(quotient[9]), .Y(n86) );
  MX2X1 U134 ( .A(n83), .B(\u_div/SumTmp[5][8] ), .S0(quotient[5]), .Y(n87) );
  MX2X1 U135 ( .A(n84), .B(\u_div/SumTmp[6][8] ), .S0(quotient[6]), .Y(n88) );
  MX2X1 U136 ( .A(n85), .B(\u_div/SumTmp[7][8] ), .S0(quotient[7]), .Y(n89) );
  MX2X1 U137 ( .A(n86), .B(\u_div/SumTmp[8][8] ), .S0(quotient[8]), .Y(n90) );
  MX2X1 U138 ( .A(n96), .B(\u_div/SumTmp[9][8] ), .S0(quotient[9]), .Y(n91) );
  MX2X1 U139 ( .A(n79), .B(\u_div/SumTmp[3][6] ), .S0(quotient[3]), .Y(n92) );
  MX2X1 U140 ( .A(n80), .B(\u_div/SumTmp[3][7] ), .S0(quotient[3]), .Y(n93) );
  MX2X1 U141 ( .A(n81), .B(\u_div/SumTmp[3][8] ), .S0(quotient[3]), .Y(n94) );
  MX2X1 U142 ( .A(n56), .B(\u_div/SumTmp[10][6] ), .S0(n242), .Y(n95) );
  MX2X1 U143 ( .A(n98), .B(\u_div/SumTmp[10][7] ), .S0(n242), .Y(n96) );
  MX2X1 U144 ( .A(n99), .B(\u_div/SumTmp[10][8] ), .S0(n242), .Y(n97) );
  MX2X1 U145 ( .A(n60), .B(\u_div/SumTmp[11][6] ), .S0(\u_div/CryTmp[11][12] ), 
        .Y(n98) );
  MX2X1 U146 ( .A(n101), .B(\u_div/SumTmp[11][7] ), .S0(\u_div/CryTmp[11][12] ), .Y(n99) );
  MX2X1 U147 ( .A(n102), .B(\u_div/SumTmp[11][8] ), .S0(\u_div/CryTmp[11][12] ), .Y(n100) );
  MX2X1 U148 ( .A(n148), .B(\u_div/SumTmp[12][6] ), .S0(n210), .Y(n101) );
  MX2X1 U149 ( .A(n149), .B(\u_div/SumTmp[12][7] ), .S0(n210), .Y(n102) );
  MX2X1 U150 ( .A(n150), .B(\u_div/SumTmp[12][8] ), .S0(n210), .Y(n103) );
  MX2X1 U151 ( .A(n66), .B(\u_div/SumTmp[14][5] ), .S0(n212), .Y(n104) );
  MX2X1 U152 ( .A(n108), .B(\u_div/SumTmp[14][6] ), .S0(n212), .Y(n105) );
  MX2X1 U153 ( .A(n109), .B(\u_div/SumTmp[14][7] ), .S0(n212), .Y(n106) );
  MX2X1 U154 ( .A(n110), .B(\u_div/SumTmp[14][8] ), .S0(n212), .Y(n107) );
  MX2X1 U155 ( .A(n69), .B(\u_div/SumTmp[15][5] ), .S0(n125), .Y(n108) );
  MX2X1 U156 ( .A(n111), .B(\u_div/SumTmp[15][6] ), .S0(n125), .Y(n109) );
  MX2X1 U157 ( .A(n112), .B(\u_div/SumTmp[15][7] ), .S0(n125), .Y(n110) );
  MX2X1 U158 ( .A(n71), .B(\u_div/SumTmp[16][5] ), .S0(n213), .Y(n111) );
  MX2X1 U159 ( .A(n113), .B(\u_div/SumTmp[16][6] ), .S0(n213), .Y(n112) );
  MX2X1 U160 ( .A(n73), .B(\u_div/SumTmp[17][5] ), .S0(n214), .Y(n113) );
  MXI2X1 U161 ( .A(n116), .B(\u_div/SumTmp[4][10] ), .S0(quotient[4]), .Y(n182) );
  MXI2X1 U162 ( .A(n117), .B(\u_div/SumTmp[5][10] ), .S0(quotient[5]), .Y(n180) );
  MXI2X1 U163 ( .A(n118), .B(\u_div/SumTmp[6][10] ), .S0(quotient[6]), .Y(n178) );
  MXI2X1 U164 ( .A(n119), .B(\u_div/SumTmp[7][10] ), .S0(quotient[7]), .Y(n176) );
  MXI2X1 U165 ( .A(n120), .B(\u_div/SumTmp[8][10] ), .S0(quotient[8]), .Y(n174) );
  MXI2X1 U166 ( .A(n122), .B(\u_div/SumTmp[9][10] ), .S0(quotient[9]), .Y(n172) );
  MXI2X1 U167 ( .A(n94), .B(\u_div/SumTmp[2][9] ), .S0(quotient[2]), .Y(n196)
         );
  MXI2X1 U168 ( .A(n93), .B(\u_div/SumTmp[2][8] ), .S0(quotient[2]), .Y(n185)
         );
  MXI2X1 U169 ( .A(n121), .B(\u_div/SumTmp[2][10] ), .S0(quotient[2]), .Y(n195) );
  MXI2X1 U170 ( .A(n115), .B(\u_div/SumTmp[3][10] ), .S0(quotient[3]), .Y(n184) );
  MXI2X1 U171 ( .A(n123), .B(\u_div/SumTmp[10][10] ), .S0(n242), .Y(n170) );
  MXI2X1 U172 ( .A(n124), .B(\u_div/SumTmp[11][10] ), .S0(
        \u_div/CryTmp[11][12] ), .Y(n223) );
  MXI2X1 U173 ( .A(n152), .B(\u_div/SumTmp[12][10] ), .S0(n210), .Y(n208) );
  MXI2X1 U174 ( .A(n186), .B(n197), .S0(quotient[1]), .Y(\u_div/PartRem[1][9] ) );
  INVX1 U175 ( .A(\u_div/SumTmp[1][8] ), .Y(n197) );
  MX2X1 U176 ( .A(n82), .B(\u_div/SumTmp[4][8] ), .S0(quotient[4]), .Y(n114)
         );
  MX2X1 U177 ( .A(n87), .B(\u_div/SumTmp[4][9] ), .S0(quotient[4]), .Y(n115)
         );
  MX2X1 U178 ( .A(n88), .B(\u_div/SumTmp[5][9] ), .S0(quotient[5]), .Y(n116)
         );
  MX2X1 U179 ( .A(n89), .B(\u_div/SumTmp[6][9] ), .S0(quotient[6]), .Y(n117)
         );
  MX2X1 U180 ( .A(n90), .B(\u_div/SumTmp[7][9] ), .S0(quotient[7]), .Y(n118)
         );
  MX2X1 U181 ( .A(n91), .B(\u_div/SumTmp[8][9] ), .S0(quotient[8]), .Y(n119)
         );
  MX2X1 U182 ( .A(n97), .B(\u_div/SumTmp[9][9] ), .S0(quotient[9]), .Y(n120)
         );
  MX2X1 U183 ( .A(n114), .B(\u_div/SumTmp[3][9] ), .S0(quotient[3]), .Y(n121)
         );
  MX2X1 U184 ( .A(n100), .B(\u_div/SumTmp[10][9] ), .S0(n242), .Y(n122) );
  MX2X1 U185 ( .A(n103), .B(\u_div/SumTmp[11][9] ), .S0(\u_div/CryTmp[11][12] ), .Y(n123) );
  MX2X1 U186 ( .A(n151), .B(\u_div/SumTmp[12][9] ), .S0(n210), .Y(n124) );
  MXI2X1 U187 ( .A(n196), .B(n206), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][11] ) );
  INVX1 U188 ( .A(\u_div/SumTmp[1][10] ), .Y(n206) );
  CLKINVX3 U189 ( .A(n229), .Y(n210) );
  NAND2BX1 U190 ( .AN(n240), .B(\u_div/CryTmp[12][11] ), .Y(n229) );
  CLKINVX3 U191 ( .A(n231), .Y(n212) );
  NAND2BX1 U192 ( .AN(n232), .B(\u_div/CryTmp[14][9] ), .Y(n231) );
  AND2X2 U193 ( .A(\u_div/CryTmp[15][8] ), .B(n161), .Y(n125) );
  CLKINVX3 U194 ( .A(n235), .Y(n214) );
  NAND3BX1 U195 ( .AN(n234), .B(\u_div/BInv [6]), .C(\u_div/CryTmp[17][6] ), 
        .Y(n235) );
  INVX1 U196 ( .A(n236), .Y(n215) );
  NAND2BX1 U197 ( .AN(n227), .B(\u_div/CryTmp[18][5] ), .Y(n236) );
  INVX1 U198 ( .A(n237), .Y(n216) );
  NAND3BX1 U199 ( .AN(n227), .B(\u_div/BInv [4]), .C(\u_div/CryTmp[19][4] ), 
        .Y(n237) );
  NAND2X1 U200 ( .A(n161), .B(\u_div/BInv [7]), .Y(n234) );
  NAND2BX1 U201 ( .AN(n220), .B(\u_div/CryTmp[20][3] ), .Y(n226) );
  MX2X1 U202 ( .A(n11), .B(\u_div/SumTmp[12][1] ), .S0(n210), .Y(n126) );
  MX2X1 U203 ( .A(n2), .B(\u_div/SumTmp[14][1] ), .S0(n212), .Y(n127) );
  MX2X1 U204 ( .A(n15), .B(\u_div/SumTmp[15][1] ), .S0(n125), .Y(n128) );
  MX2X1 U205 ( .A(n18), .B(\u_div/SumTmp[16][1] ), .S0(n213), .Y(n129) );
  MX2X1 U206 ( .A(n1), .B(\u_div/SumTmp[17][1] ), .S0(n214), .Y(n130) );
  MX2X1 U207 ( .A(n13), .B(\u_div/SumTmp[13][1] ), .S0(n241), .Y(n131) );
  MXI2X1 U208 ( .A(n193), .B(n204), .S0(quotient[1]), .Y(\u_div/PartRem[1][2] ) );
  INVX1 U209 ( .A(\u_div/SumTmp[1][1] ), .Y(n204) );
  INVX1 U210 ( .A(n192), .Y(\u_div/PartRem[2][2] ) );
  INVX1 U211 ( .A(n191), .Y(\u_div/PartRem[2][3] ) );
  MXI2X1 U212 ( .A(n191), .B(n202), .S0(quotient[1]), .Y(\u_div/PartRem[1][4] ) );
  INVX1 U213 ( .A(\u_div/SumTmp[1][3] ), .Y(n202) );
  INVX1 U214 ( .A(n190), .Y(\u_div/PartRem[2][4] ) );
  INVX1 U215 ( .A(n189), .Y(\u_div/PartRem[2][5] ) );
  MXI2X1 U216 ( .A(n189), .B(n200), .S0(quotient[1]), .Y(\u_div/PartRem[1][6] ) );
  INVX1 U217 ( .A(\u_div/SumTmp[1][5] ), .Y(n200) );
  INVX1 U218 ( .A(n188), .Y(\u_div/PartRem[2][6] ) );
  INVX1 U219 ( .A(n187), .Y(\u_div/PartRem[2][7] ) );
  MXI2X1 U220 ( .A(n187), .B(n198), .S0(quotient[1]), .Y(\u_div/PartRem[1][8] ) );
  INVX1 U221 ( .A(\u_div/SumTmp[1][7] ), .Y(n198) );
  INVX1 U222 ( .A(n186), .Y(\u_div/PartRem[2][8] ) );
  INVX1 U223 ( .A(n185), .Y(\u_div/PartRem[2][9] ) );
  INVX1 U224 ( .A(n196), .Y(\u_div/PartRem[2][10] ) );
  MXI2X1 U225 ( .A(n185), .B(n207), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][10] ) );
  INVX1 U226 ( .A(\u_div/SumTmp[1][9] ), .Y(n207) );
  MXI2X1 U227 ( .A(n158), .B(\u_div/SumTmp[2][3] ), .S0(quotient[2]), .Y(n190)
         );
  MX2X1 U228 ( .A(n163), .B(\u_div/SumTmp[19][2] ), .S0(n216), .Y(n132) );
  MX2X1 U229 ( .A(n159), .B(\u_div/SumTmp[9][2] ), .S0(quotient[9]), .Y(n133)
         );
  MX2X1 U230 ( .A(n154), .B(\u_div/SumTmp[8][2] ), .S0(quotient[8]), .Y(n134)
         );
  MX2X1 U231 ( .A(n155), .B(\u_div/SumTmp[7][2] ), .S0(quotient[7]), .Y(n135)
         );
  MX2X1 U232 ( .A(n156), .B(\u_div/SumTmp[6][2] ), .S0(quotient[6]), .Y(n136)
         );
  MX2X1 U233 ( .A(n136), .B(\u_div/SumTmp[5][3] ), .S0(quotient[5]), .Y(n137)
         );
  MX2X1 U234 ( .A(n165), .B(\u_div/SumTmp[4][3] ), .S0(quotient[4]), .Y(n138)
         );
  MX2X1 U235 ( .A(n166), .B(\u_div/SumTmp[3][3] ), .S0(quotient[3]), .Y(n139)
         );
  MX2X1 U236 ( .A(n160), .B(\u_div/SumTmp[10][2] ), .S0(n242), .Y(n140) );
  MX2X1 U237 ( .A(n126), .B(\u_div/SumTmp[11][2] ), .S0(\u_div/CryTmp[11][12] ), .Y(n141) );
  MX2X1 U238 ( .A(n162), .B(\u_div/SumTmp[17][2] ), .S0(n214), .Y(n142) );
  MX2X1 U239 ( .A(n153), .B(\u_div/SumTmp[18][2] ), .S0(n215), .Y(n143) );
  MX2X1 U240 ( .A(n164), .B(\u_div/SumTmp[20][2] ), .S0(n217), .Y(n144) );
  MX2X1 U241 ( .A(n127), .B(\u_div/SumTmp[13][2] ), .S0(n241), .Y(n145) );
  MX2X1 U242 ( .A(n61), .B(\u_div/SumTmp[13][3] ), .S0(n241), .Y(n146) );
  MX2X1 U243 ( .A(n62), .B(\u_div/SumTmp[13][4] ), .S0(n241), .Y(n147) );
  MX2X1 U244 ( .A(n63), .B(\u_div/SumTmp[13][5] ), .S0(n241), .Y(n148) );
  MX2X1 U245 ( .A(n104), .B(\u_div/SumTmp[13][6] ), .S0(n241), .Y(n149) );
  MX2X1 U246 ( .A(n105), .B(\u_div/SumTmp[13][7] ), .S0(n241), .Y(n150) );
  MX2X1 U247 ( .A(n106), .B(\u_div/SumTmp[13][8] ), .S0(n241), .Y(n151) );
  MX2X1 U248 ( .A(n107), .B(\u_div/SumTmp[13][9] ), .S0(n241), .Y(n152) );
  CLKINVX3 U249 ( .A(n240), .Y(\u_div/BInv [11]) );
  NAND2BX1 U250 ( .AN(n227), .B(n228), .Y(n220) );
  NOR2X1 U251 ( .A(b[4]), .B(b[3]), .Y(n228) );
  NAND2BX1 U252 ( .AN(n234), .B(n238), .Y(n227) );
  NOR2X1 U253 ( .A(b[6]), .B(b[5]), .Y(n238) );
  MX2X1 U254 ( .A(n19), .B(\u_div/SumTmp[19][1] ), .S0(n216), .Y(n153) );
  INVX1 U255 ( .A(n225), .Y(n218) );
  NAND3BX1 U256 ( .AN(n220), .B(\u_div/BInv [2]), .C(\u_div/CryTmp[21][2] ), 
        .Y(n225) );
  BUFX3 U257 ( .A(n211), .Y(n241) );
  NOR3X1 U258 ( .A(n230), .B(n240), .C(b[10]), .Y(n211) );
  INVX1 U259 ( .A(\u_div/CryTmp[13][10] ), .Y(n230) );
  MX2X1 U260 ( .A(n12), .B(\u_div/SumTmp[9][1] ), .S0(quotient[9]), .Y(n154)
         );
  MX2X1 U261 ( .A(n6), .B(\u_div/SumTmp[8][1] ), .S0(quotient[8]), .Y(n155) );
  MX2X1 U262 ( .A(n7), .B(\u_div/SumTmp[7][1] ), .S0(quotient[7]), .Y(n156) );
  MX2X1 U263 ( .A(n8), .B(\u_div/SumTmp[6][1] ), .S0(quotient[6]), .Y(n157) );
  MX2X1 U264 ( .A(n168), .B(\u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(n158)
         );
  MX2X1 U265 ( .A(n14), .B(\u_div/SumTmp[10][1] ), .S0(n242), .Y(n159) );
  MX2X1 U266 ( .A(n4), .B(\u_div/SumTmp[11][1] ), .S0(\u_div/CryTmp[11][12] ), 
        .Y(n160) );
  XNOR2X1 U267 ( .A(\u_div/CryTmp[3][1] ), .B(a[12]), .Y(\u_div/SumTmp[12][0] ) );
  XNOR2X1 U268 ( .A(\u_div/CryTmp[3][1] ), .B(a[14]), .Y(\u_div/SumTmp[14][0] ) );
  NOR2X1 U269 ( .A(b[8]), .B(n232), .Y(n161) );
  XNOR2X1 U270 ( .A(\u_div/CryTmp[3][1] ), .B(a[15]), .Y(\u_div/SumTmp[15][0] ) );
  XNOR2X1 U271 ( .A(\u_div/CryTmp[3][1] ), .B(a[16]), .Y(\u_div/SumTmp[16][0] ) );
  XNOR2X1 U272 ( .A(\u_div/CryTmp[3][1] ), .B(a[17]), .Y(\u_div/SumTmp[17][0] ) );
  XNOR2X1 U273 ( .A(\u_div/CryTmp[3][1] ), .B(a[18]), .Y(\u_div/SumTmp[18][0] ) );
  MX2X1 U274 ( .A(n3), .B(\u_div/SumTmp[18][1] ), .S0(n215), .Y(n162) );
  XNOR2X1 U275 ( .A(\u_div/CryTmp[3][1] ), .B(a[13]), .Y(\u_div/SumTmp[13][0] ) );
  MX2X1 U276 ( .A(n17), .B(\u_div/SumTmp[20][1] ), .S0(n217), .Y(n163) );
  MX2X1 U277 ( .A(n16), .B(\u_div/SumTmp[21][1] ), .S0(n218), .Y(n164) );
  OR3XL U278 ( .A(b[9]), .B(b[10]), .C(n240), .Y(n232) );
  BUFX3 U279 ( .A(b[11]), .Y(n240) );
  OR2XL U280 ( .A(a[18]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[18][1] )
         );
  OR2XL U281 ( .A(a[17]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[17][1] )
         );
  OR2XL U282 ( .A(a[16]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[16][1] )
         );
  OR2XL U283 ( .A(a[15]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[15][1] )
         );
  OR2XL U284 ( .A(a[14]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[14][1] )
         );
  OR2XL U285 ( .A(a[12]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[12][1] )
         );
  OR2XL U286 ( .A(a[13]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[13][1] )
         );
  MXI2X1 U287 ( .A(n169), .B(\u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(n191)
         );
  MX2X1 U288 ( .A(n157), .B(\u_div/SumTmp[5][2] ), .S0(quotient[5]), .Y(n165)
         );
  MX2X1 U289 ( .A(n167), .B(\u_div/SumTmp[4][2] ), .S0(quotient[4]), .Y(n166)
         );
  BUFX3 U290 ( .A(b[1]), .Y(n239) );
  XNOR2X1 U291 ( .A(\u_div/CryTmp[3][1] ), .B(a[21]), .Y(\u_div/SumTmp[21][0] ) );
  XNOR2X1 U292 ( .A(\u_div/CryTmp[3][1] ), .B(a[19]), .Y(\u_div/SumTmp[19][0] ) );
  XNOR2X1 U293 ( .A(\u_div/CryTmp[3][1] ), .B(a[9]), .Y(\u_div/SumTmp[9][0] )
         );
  XNOR2X1 U294 ( .A(\u_div/CryTmp[3][1] ), .B(a[8]), .Y(\u_div/SumTmp[8][0] )
         );
  XNOR2X1 U295 ( .A(\u_div/CryTmp[3][1] ), .B(a[7]), .Y(\u_div/SumTmp[7][0] )
         );
  XNOR2X1 U296 ( .A(\u_div/CryTmp[3][1] ), .B(a[6]), .Y(\u_div/SumTmp[6][0] )
         );
  MX2X1 U297 ( .A(n9), .B(\u_div/SumTmp[5][1] ), .S0(quotient[5]), .Y(n167) );
  MX2X1 U298 ( .A(n10), .B(\u_div/SumTmp[4][1] ), .S0(quotient[4]), .Y(n168)
         );
  MX2X1 U299 ( .A(n5), .B(\u_div/SumTmp[3][1] ), .S0(quotient[3]), .Y(n169) );
  XNOR2X1 U300 ( .A(\u_div/CryTmp[3][1] ), .B(a[10]), .Y(\u_div/SumTmp[10][0] ) );
  XNOR2X1 U301 ( .A(\u_div/CryTmp[3][1] ), .B(a[11]), .Y(\u_div/SumTmp[11][0] ) );
  XNOR2X1 U302 ( .A(\u_div/CryTmp[3][1] ), .B(a[22]), .Y(\u_div/SumTmp[22][0] ) );
  NOR2X1 U303 ( .A(n220), .B(n221), .Y(n219) );
  XNOR2X1 U304 ( .A(\u_div/CryTmp[3][1] ), .B(a[20]), .Y(\u_div/SumTmp[20][0] ) );
  NAND2X1 U305 ( .A(\u_div/CryTmp[22][1] ), .B(n222), .Y(n221) );
  NOR2X1 U306 ( .A(b[2]), .B(n239), .Y(n222) );
  OR2XL U307 ( .A(a[22]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[22][1] )
         );
  OR2XL U308 ( .A(a[21]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[21][1] )
         );
  OR2XL U309 ( .A(a[20]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[20][1] )
         );
  OR2XL U310 ( .A(a[19]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[19][1] )
         );
  OR2XL U311 ( .A(a[10]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[10][1] )
         );
  OR2XL U312 ( .A(a[11]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[11][1] )
         );
  OR2XL U313 ( .A(a[9]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[9][1] ) );
  OR2XL U314 ( .A(a[8]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[8][1] ) );
  OR2XL U315 ( .A(a[7]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[7][1] ) );
  OR2XL U316 ( .A(a[6]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[6][1] ) );
  XNOR2X1 U317 ( .A(\u_div/CryTmp[3][1] ), .B(a[5]), .Y(\u_div/SumTmp[5][0] )
         );
  XNOR2X1 U318 ( .A(\u_div/CryTmp[3][1] ), .B(a[4]), .Y(\u_div/SumTmp[4][0] )
         );
  OR2XL U319 ( .A(a[5]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[5][1] ) );
  OR2XL U320 ( .A(a[4]), .B(\u_div/CryTmp[3][1] ), .Y(\u_div/CryTmp[4][1] ) );
  NAND2BX4 U321 ( .AN(\u_div/CryTmp[10][12] ), .B(n30), .Y(n242) );
  NAND2BX4 U322 ( .AN(\u_div/CryTmp[9][12] ), .B(n29), .Y(quotient[9]) );
  NAND2BX4 U323 ( .AN(\u_div/CryTmp[8][12] ), .B(n22), .Y(quotient[8]) );
  NAND2BX4 U324 ( .AN(\u_div/CryTmp[7][12] ), .B(n23), .Y(quotient[7]) );
  NAND2BX4 U325 ( .AN(\u_div/CryTmp[6][12] ), .B(n24), .Y(quotient[6]) );
  NAND2BX4 U326 ( .AN(\u_div/CryTmp[5][12] ), .B(n25), .Y(quotient[5]) );
  NAND2BX4 U327 ( .AN(\u_div/CryTmp[4][12] ), .B(n26), .Y(quotient[4]) );
  NAND2BX4 U328 ( .AN(\u_div/CryTmp[3][12] ), .B(n27), .Y(quotient[3]) );
  NAND2BX4 U329 ( .AN(\u_div/CryTmp[2][12] ), .B(n28), .Y(quotient[2]) );
  NAND2BX4 U330 ( .AN(\u_div/CryTmp[1][12] ), .B(n21), .Y(quotient[1]) );
  CLKINVX8 U331 ( .A(b[2]), .Y(\u_div/BInv [2]) );
  CLKINVX8 U332 ( .A(n239), .Y(\u_div/BInv [1]) );
  CLKINVX8 U333 ( .A(b[0]), .Y(\u_div/CryTmp[3][1] ) );
endmodule


module Equation_Implementation_DW_div_uns_46 ( a, b, quotient, remainder, 
        divide_by_0 );
  input [15:0] a;
  input [6:0] b;
  output [15:0] quotient;
  output [6:0] remainder;
  output divide_by_0;
  wire   \u_div/SumTmp[2][0] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[2][5] , \u_div/SumTmp[3][0] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[3][5] , \u_div/SumTmp[4][0] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[4][5] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[5][5] , \u_div/SumTmp[6][0] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[6][5] , \u_div/SumTmp[7][0] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[7][5] ,
         \u_div/SumTmp[8][0] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[8][5] , \u_div/SumTmp[9][0] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[9][5] , \u_div/CryTmp[0][3] ,
         \u_div/CryTmp[0][4] , \u_div/CryTmp[0][5] , \u_div/CryTmp[1][3] ,
         \u_div/CryTmp[1][4] , \u_div/CryTmp[1][5] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[1][7] , \u_div/CryTmp[2][3] , \u_div/CryTmp[2][4] ,
         \u_div/CryTmp[2][5] , \u_div/CryTmp[2][6] , \u_div/CryTmp[2][7] ,
         \u_div/CryTmp[3][3] , \u_div/CryTmp[3][4] , \u_div/CryTmp[3][5] ,
         \u_div/CryTmp[3][6] , \u_div/CryTmp[3][7] , \u_div/CryTmp[4][3] ,
         \u_div/CryTmp[4][4] , \u_div/CryTmp[4][5] , \u_div/CryTmp[4][6] ,
         \u_div/CryTmp[4][7] , \u_div/CryTmp[5][3] , \u_div/CryTmp[5][4] ,
         \u_div/CryTmp[5][5] , \u_div/CryTmp[5][6] , \u_div/CryTmp[5][7] ,
         \u_div/CryTmp[6][3] , \u_div/CryTmp[6][4] , \u_div/CryTmp[6][5] ,
         \u_div/CryTmp[6][6] , \u_div/CryTmp[6][7] , \u_div/CryTmp[7][3] ,
         \u_div/CryTmp[7][4] , \u_div/CryTmp[7][5] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[7][7] , \u_div/CryTmp[8][3] , \u_div/CryTmp[8][4] ,
         \u_div/CryTmp[8][5] , \u_div/CryTmp[8][6] , \u_div/CryTmp[8][7] ,
         \u_div/CryTmp[9][4] , \u_div/CryTmp[9][5] , \u_div/CryTmp[9][6] ,
         \u_div/PartRem[1][5] , \u_div/PartRem[2][3] , \u_div/PartRem[2][4] ,
         \u_div/PartRem[2][5] , \u_div/PartRem[2][6] , \u_div/PartRem[2][7] ,
         \u_div/PartRem[3][6] , \u_div/PartRem[3][7] , \u_div/PartRem[4][6] ,
         \u_div/PartRem[4][7] , \u_div/PartRem[5][6] , \u_div/PartRem[5][7] ,
         \u_div/PartRem[6][6] , \u_div/PartRem[6][7] , \u_div/PartRem[7][6] ,
         \u_div/PartRem[7][7] , \u_div/PartRem[8][6] , \u_div/PartRem[8][7] ,
         \u_div/PartRem[9][6] , \u_div/PartRem[9][7] , \u_div/PartRem[12][1] ,
         \u_div/PartRem[13][1] , \u_div/PartRem[14][1] ,
         \u_div/PartRem[15][1] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68;
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/PartRem[12][1]  = a[12];
  assign \u_div/PartRem[13][1]  = a[13];
  assign \u_div/PartRem[14][1]  = a[14];
  assign \u_div/PartRem[15][1]  = a[15];

  AND2X2 U1 ( .A(\u_div/CryTmp[8][6] ), .B(\u_div/PartRem[9][6] ), .Y(
        \u_div/CryTmp[8][7] ) );
  AND2X2 U2 ( .A(\u_div/CryTmp[1][6] ), .B(\u_div/PartRem[2][6] ), .Y(
        \u_div/CryTmp[1][7] ) );
  AND2X2 U3 ( .A(\u_div/CryTmp[2][6] ), .B(\u_div/PartRem[3][6] ), .Y(
        \u_div/CryTmp[2][7] ) );
  AND2X2 U4 ( .A(\u_div/CryTmp[3][6] ), .B(\u_div/PartRem[4][6] ), .Y(
        \u_div/CryTmp[3][7] ) );
  AND2X2 U5 ( .A(\u_div/CryTmp[4][6] ), .B(\u_div/PartRem[5][6] ), .Y(
        \u_div/CryTmp[4][7] ) );
  AND2X2 U6 ( .A(\u_div/CryTmp[5][6] ), .B(\u_div/PartRem[6][6] ), .Y(
        \u_div/CryTmp[5][7] ) );
  AND2X2 U7 ( .A(\u_div/CryTmp[6][6] ), .B(\u_div/PartRem[7][6] ), .Y(
        \u_div/CryTmp[6][7] ) );
  AND2X2 U8 ( .A(\u_div/CryTmp[7][6] ), .B(\u_div/PartRem[8][6] ), .Y(
        \u_div/CryTmp[7][7] ) );
  MX2X1 U9 ( .A(n60), .B(\u_div/CryTmp[1][3] ), .S0(quotient[1]), .Y(n1) );
  MX2X1 U10 ( .A(a[11]), .B(n68), .S0(quotient[9]), .Y(n2) );
  MX2X1 U11 ( .A(n59), .B(n25), .S0(quotient[1]), .Y(n3) );
  MX2X1 U12 ( .A(n56), .B(n27), .S0(quotient[1]), .Y(n4) );
  MX2X1 U13 ( .A(\u_div/CryTmp[3][3] ), .B(n64), .S0(quotient[3]), .Y(n5) );
  MX2X1 U14 ( .A(\u_div/CryTmp[8][3] ), .B(n51), .S0(quotient[8]), .Y(n6) );
  MX2X1 U15 ( .A(\u_div/CryTmp[7][3] ), .B(n53), .S0(quotient[7]), .Y(n7) );
  MX2X1 U16 ( .A(\u_div/CryTmp[6][3] ), .B(n55), .S0(quotient[6]), .Y(n8) );
  MX2X1 U17 ( .A(\u_div/CryTmp[5][3] ), .B(n62), .S0(quotient[5]), .Y(n9) );
  MX2X1 U18 ( .A(\u_div/CryTmp[4][3] ), .B(n63), .S0(quotient[4]), .Y(n10) );
  MX2X1 U19 ( .A(n10), .B(\u_div/SumTmp[3][3] ), .S0(quotient[3]), .Y(n11) );
  MX2X1 U20 ( .A(n6), .B(\u_div/SumTmp[7][3] ), .S0(quotient[7]), .Y(n12) );
  MX2X1 U21 ( .A(n7), .B(\u_div/SumTmp[6][3] ), .S0(quotient[6]), .Y(n13) );
  MX2X1 U22 ( .A(n8), .B(\u_div/SumTmp[5][3] ), .S0(quotient[5]), .Y(n14) );
  MX2X1 U23 ( .A(n9), .B(\u_div/SumTmp[4][3] ), .S0(quotient[4]), .Y(n15) );
  MX2X1 U24 ( .A(n2), .B(\u_div/SumTmp[8][3] ), .S0(quotient[8]), .Y(n16) );
  MX2X1 U25 ( .A(\u_div/PartRem[12][1] ), .B(\u_div/SumTmp[9][3] ), .S0(
        quotient[9]), .Y(n17) );
  MX2X1 U26 ( .A(n12), .B(\u_div/SumTmp[6][4] ), .S0(quotient[6]), .Y(n18) );
  MX2X1 U27 ( .A(n13), .B(\u_div/SumTmp[5][4] ), .S0(quotient[5]), .Y(n19) );
  MX2X1 U28 ( .A(n14), .B(\u_div/SumTmp[4][4] ), .S0(quotient[4]), .Y(n20) );
  MX2X1 U29 ( .A(n15), .B(\u_div/SumTmp[3][4] ), .S0(quotient[3]), .Y(n21) );
  MX2X1 U30 ( .A(n16), .B(\u_div/SumTmp[7][4] ), .S0(quotient[7]), .Y(n22) );
  MX2X1 U31 ( .A(n17), .B(\u_div/SumTmp[8][4] ), .S0(quotient[8]), .Y(n23) );
  MX2X1 U32 ( .A(\u_div/PartRem[13][1] ), .B(\u_div/SumTmp[9][4] ), .S0(
        quotient[9]), .Y(n24) );
  XOR2X1 U33 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/CryTmp[1][3] ), .Y(n25) );
  XOR2X1 U34 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/CryTmp[1][4] ), .Y(n26) );
  XNOR2X1 U35 ( .A(\u_div/PartRem[2][6] ), .B(\u_div/CryTmp[1][6] ), .Y(n27)
         );
  MX2X1 U36 ( .A(\u_div/SumTmp[9][0] ), .B(\u_div/SumTmp[9][0] ), .S0(
        quotient[9]), .Y(n28) );
  MX2X1 U37 ( .A(\u_div/SumTmp[8][0] ), .B(\u_div/SumTmp[8][0] ), .S0(
        quotient[8]), .Y(n29) );
  MX2X1 U38 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[7][0] ), .S0(
        quotient[7]), .Y(n30) );
  MX2X1 U39 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[6][0] ), .S0(
        quotient[6]), .Y(n31) );
  MX2X1 U40 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[5][0] ), .S0(
        quotient[5]), .Y(n32) );
  MX2X1 U41 ( .A(\u_div/SumTmp[4][0] ), .B(\u_div/SumTmp[4][0] ), .S0(
        quotient[4]), .Y(n33) );
  OR2X2 U42 ( .A(\u_div/CryTmp[3][7] ), .B(\u_div/PartRem[4][7] ), .Y(
        quotient[3]) );
  MXI2X1 U43 ( .A(n50), .B(n35), .S0(quotient[4]), .Y(\u_div/PartRem[4][7] )
         );
  OR2X2 U44 ( .A(\u_div/CryTmp[2][7] ), .B(\u_div/PartRem[3][7] ), .Y(
        quotient[2]) );
  MXI2X1 U45 ( .A(n52), .B(n36), .S0(quotient[3]), .Y(\u_div/PartRem[3][7] )
         );
  OR2X2 U46 ( .A(\u_div/CryTmp[1][7] ), .B(\u_div/PartRem[2][7] ), .Y(
        quotient[1]) );
  MXI2X1 U47 ( .A(n54), .B(n37), .S0(quotient[2]), .Y(\u_div/PartRem[2][7] )
         );
  INVX1 U48 ( .A(n50), .Y(\u_div/PartRem[5][6] ) );
  INVX1 U49 ( .A(n52), .Y(\u_div/PartRem[4][6] ) );
  INVX1 U50 ( .A(n54), .Y(\u_div/PartRem[3][6] ) );
  INVX1 U51 ( .A(n56), .Y(\u_div/PartRem[2][6] ) );
  XNOR2X1 U52 ( .A(\u_div/PartRem[6][6] ), .B(\u_div/CryTmp[5][6] ), .Y(n34)
         );
  XNOR2X1 U53 ( .A(\u_div/PartRem[5][6] ), .B(\u_div/CryTmp[4][6] ), .Y(n35)
         );
  XNOR2X1 U54 ( .A(\u_div/PartRem[4][6] ), .B(\u_div/CryTmp[3][6] ), .Y(n36)
         );
  XNOR2X1 U55 ( .A(\u_div/PartRem[3][6] ), .B(\u_div/CryTmp[2][6] ), .Y(n37)
         );
  OR2X2 U56 ( .A(\u_div/CryTmp[4][7] ), .B(\u_div/PartRem[5][7] ), .Y(
        quotient[4]) );
  MXI2X1 U57 ( .A(n49), .B(n34), .S0(quotient[5]), .Y(\u_div/PartRem[5][7] )
         );
  AND2X2 U58 ( .A(\u_div/CryTmp[5][5] ), .B(n18), .Y(\u_div/CryTmp[5][6] ) );
  AND2X2 U59 ( .A(\u_div/CryTmp[4][5] ), .B(n19), .Y(\u_div/CryTmp[4][6] ) );
  AND2X2 U60 ( .A(\u_div/CryTmp[3][5] ), .B(n20), .Y(\u_div/CryTmp[3][6] ) );
  AND2X2 U61 ( .A(\u_div/CryTmp[2][5] ), .B(n21), .Y(\u_div/CryTmp[2][6] ) );
  AND2X2 U62 ( .A(\u_div/CryTmp[1][5] ), .B(\u_div/PartRem[2][5] ), .Y(
        \u_div/CryTmp[1][6] ) );
  INVX1 U63 ( .A(n57), .Y(\u_div/PartRem[2][5] ) );
  MXI2X1 U64 ( .A(n18), .B(\u_div/SumTmp[5][5] ), .S0(quotient[5]), .Y(n50) );
  XOR2X1 U65 ( .A(n18), .B(\u_div/CryTmp[5][5] ), .Y(\u_div/SumTmp[5][5] ) );
  MXI2X1 U66 ( .A(n19), .B(\u_div/SumTmp[4][5] ), .S0(quotient[4]), .Y(n52) );
  XOR2X1 U67 ( .A(n19), .B(\u_div/CryTmp[4][5] ), .Y(\u_div/SumTmp[4][5] ) );
  MXI2X1 U68 ( .A(n20), .B(\u_div/SumTmp[3][5] ), .S0(quotient[3]), .Y(n54) );
  XOR2X1 U69 ( .A(n20), .B(\u_div/CryTmp[3][5] ), .Y(\u_div/SumTmp[3][5] ) );
  MXI2X1 U70 ( .A(n21), .B(\u_div/SumTmp[2][5] ), .S0(quotient[2]), .Y(n56) );
  XOR2X1 U71 ( .A(n21), .B(\u_div/CryTmp[2][5] ), .Y(\u_div/SumTmp[2][5] ) );
  INVX1 U72 ( .A(n49), .Y(\u_div/PartRem[6][6] ) );
  XNOR2X1 U73 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/CryTmp[1][5] ), .Y(n38)
         );
  XNOR2X1 U74 ( .A(\u_div/PartRem[7][6] ), .B(\u_div/CryTmp[6][6] ), .Y(n39)
         );
  OR2X2 U75 ( .A(\u_div/CryTmp[5][7] ), .B(\u_div/PartRem[6][7] ), .Y(
        quotient[5]) );
  MXI2X1 U76 ( .A(n48), .B(n39), .S0(quotient[6]), .Y(\u_div/PartRem[6][7] )
         );
  AND2X2 U77 ( .A(\u_div/CryTmp[6][5] ), .B(n22), .Y(\u_div/CryTmp[6][6] ) );
  OR2X2 U78 ( .A(\u_div/CryTmp[6][4] ), .B(n12), .Y(\u_div/CryTmp[6][5] ) );
  OR2X2 U79 ( .A(\u_div/CryTmp[5][4] ), .B(n13), .Y(\u_div/CryTmp[5][5] ) );
  OR2X2 U80 ( .A(\u_div/CryTmp[4][4] ), .B(n14), .Y(\u_div/CryTmp[4][5] ) );
  OR2X2 U81 ( .A(\u_div/CryTmp[3][4] ), .B(n15), .Y(\u_div/CryTmp[3][5] ) );
  OR2X2 U82 ( .A(\u_div/CryTmp[2][4] ), .B(n11), .Y(\u_div/CryTmp[2][5] ) );
  OR2X2 U83 ( .A(\u_div/CryTmp[1][4] ), .B(\u_div/PartRem[2][4] ), .Y(
        \u_div/CryTmp[1][5] ) );
  MXI2X1 U84 ( .A(n11), .B(\u_div/SumTmp[2][4] ), .S0(quotient[2]), .Y(n57) );
  XNOR2X1 U85 ( .A(n11), .B(\u_div/CryTmp[2][4] ), .Y(\u_div/SumTmp[2][4] ) );
  XNOR2X1 U86 ( .A(n12), .B(\u_div/CryTmp[6][4] ), .Y(\u_div/SumTmp[6][4] ) );
  XNOR2X1 U87 ( .A(n13), .B(\u_div/CryTmp[5][4] ), .Y(\u_div/SumTmp[5][4] ) );
  XNOR2X1 U88 ( .A(n14), .B(\u_div/CryTmp[4][4] ), .Y(\u_div/SumTmp[4][4] ) );
  XNOR2X1 U89 ( .A(n15), .B(\u_div/CryTmp[3][4] ), .Y(\u_div/SumTmp[3][4] ) );
  INVX1 U90 ( .A(n59), .Y(\u_div/PartRem[2][3] ) );
  INVX1 U91 ( .A(n58), .Y(\u_div/PartRem[2][4] ) );
  MXI2X1 U92 ( .A(n22), .B(\u_div/SumTmp[6][5] ), .S0(quotient[6]), .Y(n49) );
  XOR2X1 U93 ( .A(n22), .B(\u_div/CryTmp[6][5] ), .Y(\u_div/SumTmp[6][5] ) );
  INVX1 U94 ( .A(n48), .Y(\u_div/PartRem[7][6] ) );
  XNOR2X1 U95 ( .A(\u_div/PartRem[8][6] ), .B(\u_div/CryTmp[7][6] ), .Y(n40)
         );
  XNOR2X1 U96 ( .A(\u_div/PartRem[9][6] ), .B(\u_div/CryTmp[8][6] ), .Y(n41)
         );
  OR2X2 U97 ( .A(\u_div/CryTmp[6][7] ), .B(\u_div/PartRem[7][7] ), .Y(
        quotient[6]) );
  MXI2X1 U98 ( .A(n47), .B(n40), .S0(quotient[7]), .Y(\u_div/PartRem[7][7] )
         );
  OR2X2 U99 ( .A(\u_div/CryTmp[8][3] ), .B(n2), .Y(\u_div/CryTmp[8][4] ) );
  OR2X2 U100 ( .A(\u_div/CryTmp[7][3] ), .B(n6), .Y(\u_div/CryTmp[7][4] ) );
  OR2X2 U101 ( .A(\u_div/CryTmp[6][3] ), .B(n7), .Y(\u_div/CryTmp[6][4] ) );
  OR2X2 U102 ( .A(\u_div/CryTmp[5][3] ), .B(n8), .Y(\u_div/CryTmp[5][4] ) );
  OR2X2 U103 ( .A(\u_div/CryTmp[4][3] ), .B(n9), .Y(\u_div/CryTmp[4][4] ) );
  OR2X2 U104 ( .A(\u_div/CryTmp[3][3] ), .B(n10), .Y(\u_div/CryTmp[3][4] ) );
  OR2X2 U105 ( .A(\u_div/CryTmp[2][3] ), .B(n5), .Y(\u_div/CryTmp[2][4] ) );
  AND2X2 U106 ( .A(\u_div/CryTmp[8][5] ), .B(n24), .Y(\u_div/CryTmp[8][6] ) );
  AND2X2 U107 ( .A(\u_div/CryTmp[7][5] ), .B(n23), .Y(\u_div/CryTmp[7][6] ) );
  OR2X2 U108 ( .A(\u_div/CryTmp[1][3] ), .B(\u_div/PartRem[2][3] ), .Y(
        \u_div/CryTmp[1][4] ) );
  OR2X2 U109 ( .A(\u_div/CryTmp[8][4] ), .B(n17), .Y(\u_div/CryTmp[8][5] ) );
  OR2X2 U110 ( .A(\u_div/CryTmp[7][4] ), .B(n16), .Y(\u_div/CryTmp[7][5] ) );
  NOR2X1 U111 ( .A(n43), .B(n45), .Y(n42) );
  MX2X1 U112 ( .A(n57), .B(n38), .S0(quotient[1]), .Y(n43) );
  MXI2X1 U113 ( .A(\u_div/CryTmp[2][3] ), .B(n65), .S0(quotient[2]), .Y(n59)
         );
  MXI2X1 U114 ( .A(n5), .B(\u_div/SumTmp[2][3] ), .S0(quotient[2]), .Y(n58) );
  XNOR2X1 U115 ( .A(n5), .B(\u_div/CryTmp[2][3] ), .Y(\u_div/SumTmp[2][3] ) );
  XNOR2X1 U116 ( .A(n16), .B(\u_div/CryTmp[7][4] ), .Y(\u_div/SumTmp[7][4] )
         );
  XNOR2X1 U117 ( .A(n6), .B(\u_div/CryTmp[7][3] ), .Y(\u_div/SumTmp[7][3] ) );
  XNOR2X1 U118 ( .A(n7), .B(\u_div/CryTmp[6][3] ), .Y(\u_div/SumTmp[6][3] ) );
  XNOR2X1 U119 ( .A(n8), .B(\u_div/CryTmp[5][3] ), .Y(\u_div/SumTmp[5][3] ) );
  XNOR2X1 U120 ( .A(n9), .B(\u_div/CryTmp[4][3] ), .Y(\u_div/SumTmp[4][3] ) );
  XNOR2X1 U121 ( .A(n10), .B(\u_div/CryTmp[3][3] ), .Y(\u_div/SumTmp[3][3] )
         );
  MXI2X1 U122 ( .A(n23), .B(\u_div/SumTmp[7][5] ), .S0(quotient[7]), .Y(n48)
         );
  XOR2X1 U123 ( .A(n23), .B(\u_div/CryTmp[7][5] ), .Y(\u_div/SumTmp[7][5] ) );
  INVX1 U124 ( .A(n47), .Y(\u_div/PartRem[8][6] ) );
  INVX1 U125 ( .A(n46), .Y(\u_div/PartRem[9][6] ) );
  OR2X2 U126 ( .A(\u_div/CryTmp[7][7] ), .B(\u_div/PartRem[8][7] ), .Y(
        quotient[7]) );
  MXI2X1 U127 ( .A(n46), .B(n41), .S0(quotient[8]), .Y(\u_div/PartRem[8][7] )
         );
  AND2X2 U128 ( .A(\u_div/CryTmp[9][6] ), .B(\u_div/PartRem[15][1] ), .Y(
        quotient[9]) );
  INVX1 U129 ( .A(n53), .Y(\u_div/CryTmp[7][3] ) );
  MXI2X1 U130 ( .A(n28), .B(n28), .S0(quotient[8]), .Y(n53) );
  INVX1 U131 ( .A(n55), .Y(\u_div/CryTmp[6][3] ) );
  MXI2X1 U132 ( .A(n29), .B(n29), .S0(quotient[7]), .Y(n55) );
  INVX1 U133 ( .A(n62), .Y(\u_div/CryTmp[5][3] ) );
  MXI2X1 U134 ( .A(n30), .B(n30), .S0(quotient[6]), .Y(n62) );
  INVX1 U135 ( .A(n63), .Y(\u_div/CryTmp[4][3] ) );
  MXI2X1 U136 ( .A(n31), .B(n31), .S0(quotient[5]), .Y(n63) );
  INVX1 U137 ( .A(n64), .Y(\u_div/CryTmp[3][3] ) );
  MXI2X1 U138 ( .A(n32), .B(n32), .S0(quotient[4]), .Y(n64) );
  INVX1 U139 ( .A(n65), .Y(\u_div/CryTmp[2][3] ) );
  MXI2X1 U140 ( .A(n33), .B(n33), .S0(quotient[3]), .Y(n65) );
  INVX1 U141 ( .A(n51), .Y(\u_div/CryTmp[8][3] ) );
  MXI2X1 U142 ( .A(a[10]), .B(a[10]), .S0(quotient[9]), .Y(n51) );
  INVX1 U143 ( .A(n60), .Y(\u_div/CryTmp[1][3] ) );
  AND2X2 U144 ( .A(\u_div/CryTmp[9][5] ), .B(\u_div/PartRem[14][1] ), .Y(
        \u_div/CryTmp[9][6] ) );
  OR2X2 U145 ( .A(\u_div/CryTmp[9][4] ), .B(\u_div/PartRem[13][1] ), .Y(
        \u_div/CryTmp[9][5] ) );
  NAND2X1 U146 ( .A(\u_div/PartRem[1][5] ), .B(\u_div/CryTmp[0][5] ), .Y(n45)
         );
  MXI2X1 U147 ( .A(n58), .B(n26), .S0(quotient[1]), .Y(\u_div/PartRem[1][5] )
         );
  NAND2BX1 U148 ( .AN(\u_div/CryTmp[0][4] ), .B(n3), .Y(\u_div/CryTmp[0][5] )
         );
  INVX1 U149 ( .A(a[11]), .Y(n68) );
  XNOR2X1 U150 ( .A(n17), .B(\u_div/CryTmp[8][4] ), .Y(\u_div/SumTmp[8][4] )
         );
  XNOR2X1 U151 ( .A(\u_div/PartRem[13][1] ), .B(\u_div/CryTmp[9][4] ), .Y(
        \u_div/SumTmp[9][4] ) );
  XNOR2X1 U152 ( .A(n2), .B(\u_div/CryTmp[8][3] ), .Y(\u_div/SumTmp[8][3] ) );
  XNOR2X1 U153 ( .A(\u_div/PartRem[12][1] ), .B(a[11]), .Y(
        \u_div/SumTmp[9][3] ) );
  OR2X2 U154 ( .A(a[11]), .B(\u_div/PartRem[12][1] ), .Y(\u_div/CryTmp[9][4] )
         );
  MXI2X1 U155 ( .A(n24), .B(\u_div/SumTmp[8][5] ), .S0(quotient[8]), .Y(n47)
         );
  XOR2X1 U156 ( .A(n24), .B(\u_div/CryTmp[8][5] ), .Y(\u_div/SumTmp[8][5] ) );
  MXI2X1 U157 ( .A(\u_div/PartRem[14][1] ), .B(\u_div/SumTmp[9][5] ), .S0(
        quotient[9]), .Y(n46) );
  XOR2X1 U158 ( .A(\u_div/PartRem[14][1] ), .B(\u_div/CryTmp[9][5] ), .Y(
        \u_div/SumTmp[9][5] ) );
  XNOR2X1 U159 ( .A(\u_div/PartRem[15][1] ), .B(\u_div/CryTmp[9][6] ), .Y(n44)
         );
  OR2X2 U160 ( .A(\u_div/CryTmp[8][7] ), .B(\u_div/PartRem[9][7] ), .Y(
        quotient[8]) );
  MXI2X1 U161 ( .A(n67), .B(n44), .S0(quotient[9]), .Y(\u_div/PartRem[9][7] )
         );
  MX2X1 U162 ( .A(n66), .B(n66), .S0(quotient[2]), .Y(n60) );
  MXI2X1 U163 ( .A(\u_div/SumTmp[3][0] ), .B(\u_div/SumTmp[3][0] ), .S0(
        quotient[3]), .Y(n66) );
  NAND2BX1 U164 ( .AN(\u_div/CryTmp[0][3] ), .B(n1), .Y(\u_div/CryTmp[0][4] )
         );
  MXI2X1 U165 ( .A(n61), .B(n61), .S0(quotient[1]), .Y(\u_div/CryTmp[0][3] )
         );
  INVX1 U166 ( .A(\u_div/PartRem[15][1] ), .Y(n67) );
  MXI2X1 U167 ( .A(\u_div/SumTmp[2][0] ), .B(\u_div/SumTmp[2][0] ), .S0(
        quotient[2]), .Y(n61) );
  NAND2BX1 U168 ( .AN(n42), .B(n4), .Y(quotient[0]) );
endmodule


module Equation_Implementation_DW_div_uns_52 ( a, b, quotient, remainder, 
        divide_by_0 );
  input [18:0] a;
  input [9:0] b;
  output [18:0] quotient;
  output [9:0] remainder;
  output divide_by_0;
  wire   \u_div/SumTmp[2][4] , \u_div/SumTmp[2][5] , \u_div/SumTmp[2][6] ,
         \u_div/SumTmp[2][7] , \u_div/SumTmp[2][8] , \u_div/SumTmp[3][0] ,
         \u_div/SumTmp[3][4] , \u_div/SumTmp[3][5] , \u_div/SumTmp[3][6] ,
         \u_div/SumTmp[3][7] , \u_div/SumTmp[3][8] , \u_div/SumTmp[4][0] ,
         \u_div/SumTmp[4][4] , \u_div/SumTmp[4][5] , \u_div/SumTmp[4][6] ,
         \u_div/SumTmp[4][7] , \u_div/SumTmp[4][8] , \u_div/SumTmp[5][0] ,
         \u_div/SumTmp[5][4] , \u_div/SumTmp[5][5] , \u_div/SumTmp[5][6] ,
         \u_div/SumTmp[5][7] , \u_div/SumTmp[5][8] , \u_div/SumTmp[6][0] ,
         \u_div/SumTmp[6][4] , \u_div/SumTmp[6][5] , \u_div/SumTmp[6][6] ,
         \u_div/SumTmp[6][7] , \u_div/SumTmp[6][8] , \u_div/SumTmp[7][0] ,
         \u_div/SumTmp[7][4] , \u_div/SumTmp[7][5] , \u_div/SumTmp[7][6] ,
         \u_div/SumTmp[7][7] , \u_div/SumTmp[7][8] , \u_div/SumTmp[8][0] ,
         \u_div/SumTmp[8][4] , \u_div/SumTmp[8][5] , \u_div/SumTmp[8][6] ,
         \u_div/SumTmp[8][7] , \u_div/SumTmp[8][8] , \u_div/SumTmp[9][0] ,
         \u_div/SumTmp[9][4] , \u_div/SumTmp[9][5] , \u_div/SumTmp[9][6] ,
         \u_div/SumTmp[9][7] , \u_div/SumTmp[9][8] , \u_div/CryTmp[0][4] ,
         \u_div/CryTmp[0][5] , \u_div/CryTmp[1][4] , \u_div/CryTmp[1][5] ,
         \u_div/CryTmp[1][6] , \u_div/CryTmp[1][7] , \u_div/CryTmp[1][8] ,
         \u_div/CryTmp[1][9] , \u_div/CryTmp[1][10] , \u_div/CryTmp[2][4] ,
         \u_div/CryTmp[2][5] , \u_div/CryTmp[2][6] , \u_div/CryTmp[2][7] ,
         \u_div/CryTmp[2][8] , \u_div/CryTmp[2][9] , \u_div/CryTmp[2][10] ,
         \u_div/CryTmp[3][4] , \u_div/CryTmp[3][5] , \u_div/CryTmp[3][6] ,
         \u_div/CryTmp[3][7] , \u_div/CryTmp[3][8] , \u_div/CryTmp[3][9] ,
         \u_div/CryTmp[3][10] , \u_div/CryTmp[4][4] , \u_div/CryTmp[4][5] ,
         \u_div/CryTmp[4][6] , \u_div/CryTmp[4][7] , \u_div/CryTmp[4][8] ,
         \u_div/CryTmp[4][9] , \u_div/CryTmp[4][10] , \u_div/CryTmp[5][4] ,
         \u_div/CryTmp[5][5] , \u_div/CryTmp[5][6] , \u_div/CryTmp[5][7] ,
         \u_div/CryTmp[5][8] , \u_div/CryTmp[5][9] , \u_div/CryTmp[5][10] ,
         \u_div/CryTmp[6][4] , \u_div/CryTmp[6][5] , \u_div/CryTmp[6][6] ,
         \u_div/CryTmp[6][7] , \u_div/CryTmp[6][8] , \u_div/CryTmp[6][9] ,
         \u_div/CryTmp[6][10] , \u_div/CryTmp[7][4] , \u_div/CryTmp[7][5] ,
         \u_div/CryTmp[7][6] , \u_div/CryTmp[7][7] , \u_div/CryTmp[7][8] ,
         \u_div/CryTmp[7][9] , \u_div/CryTmp[7][10] , \u_div/CryTmp[8][4] ,
         \u_div/CryTmp[8][5] , \u_div/CryTmp[8][6] , \u_div/CryTmp[8][7] ,
         \u_div/CryTmp[8][8] , \u_div/CryTmp[8][9] , \u_div/CryTmp[8][10] ,
         \u_div/CryTmp[9][5] , \u_div/CryTmp[9][6] , \u_div/CryTmp[9][7] ,
         \u_div/CryTmp[9][8] , \u_div/CryTmp[9][9] , \u_div/PartRem[1][5] ,
         \u_div/PartRem[1][6] , \u_div/PartRem[1][7] , \u_div/PartRem[1][8] ,
         \u_div/PartRem[1][9] , \u_div/PartRem[2][4] , \u_div/PartRem[2][5] ,
         \u_div/PartRem[2][6] , \u_div/PartRem[2][7] , \u_div/PartRem[2][8] ,
         \u_div/PartRem[2][9] , \u_div/PartRem[2][10] , \u_div/PartRem[3][9] ,
         \u_div/PartRem[3][10] , \u_div/PartRem[4][9] , \u_div/PartRem[4][10] ,
         \u_div/PartRem[5][9] , \u_div/PartRem[6][9] , \u_div/PartRem[7][9] ,
         \u_div/PartRem[8][9] , \u_div/PartRem[9][9] , \u_div/PartRem[15][1] ,
         \u_div/PartRem[16][1] , \u_div/PartRem[17][1] ,
         \u_div/PartRem[18][1] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99;
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/PartRem[15][1]  = a[15];
  assign \u_div/PartRem[16][1]  = a[16];
  assign \u_div/PartRem[17][1]  = a[17];
  assign \u_div/PartRem[18][1]  = a[18];

  NAND2BX2 U1 ( .AN(\u_div/CryTmp[8][10] ), .B(n69), .Y(quotient[8]) );
  AND2X2 U2 ( .A(\u_div/CryTmp[1][9] ), .B(\u_div/PartRem[2][9] ), .Y(
        \u_div/CryTmp[1][10] ) );
  AND2X2 U3 ( .A(\u_div/CryTmp[2][9] ), .B(\u_div/PartRem[3][9] ), .Y(
        \u_div/CryTmp[2][10] ) );
  AND2X2 U4 ( .A(\u_div/CryTmp[3][9] ), .B(\u_div/PartRem[4][9] ), .Y(
        \u_div/CryTmp[3][10] ) );
  NAND2BX2 U5 ( .AN(\u_div/CryTmp[4][10] ), .B(n61), .Y(quotient[4]) );
  NAND2BX2 U6 ( .AN(\u_div/CryTmp[5][10] ), .B(n63), .Y(quotient[5]) );
  NAND2BX2 U7 ( .AN(\u_div/CryTmp[6][10] ), .B(n65), .Y(quotient[6]) );
  NAND2BX2 U8 ( .AN(\u_div/CryTmp[7][10] ), .B(n67), .Y(quotient[7]) );
  MX2X1 U9 ( .A(a[12]), .B(n99), .S0(quotient[9]), .Y(n1) );
  MX2X1 U10 ( .A(n90), .B(\u_div/CryTmp[1][4] ), .S0(quotient[1]), .Y(n2) );
  AND2X2 U11 ( .A(\u_div/PartRem[1][8] ), .B(n20), .Y(n3) );
  AND2X2 U12 ( .A(\u_div/PartRem[1][6] ), .B(n21), .Y(n4) );
  AND2X2 U13 ( .A(\u_div/PartRem[1][9] ), .B(n3), .Y(n5) );
  MX2X1 U14 ( .A(\u_div/CryTmp[3][4] ), .B(n95), .S0(quotient[3]), .Y(n6) );
  MX2X1 U15 ( .A(\u_div/CryTmp[7][4] ), .B(n97), .S0(quotient[7]), .Y(n7) );
  MX2X1 U16 ( .A(n35), .B(\u_div/SumTmp[3][6] ), .S0(quotient[3]), .Y(n8) );
  MX2X1 U17 ( .A(n29), .B(\u_div/SumTmp[6][6] ), .S0(quotient[6]), .Y(n9) );
  MX2X1 U18 ( .A(n30), .B(\u_div/SumTmp[5][6] ), .S0(quotient[5]), .Y(n10) );
  MX2X1 U19 ( .A(n34), .B(\u_div/SumTmp[7][6] ), .S0(quotient[7]), .Y(n11) );
  MX2X1 U20 ( .A(n36), .B(\u_div/SumTmp[8][6] ), .S0(quotient[8]), .Y(n12) );
  MX2X1 U21 ( .A(a[10]), .B(a[10]), .S0(quotient[9]), .Y(n13) );
  MX2X1 U22 ( .A(n74), .B(n74), .S0(quotient[5]), .Y(n14) );
  MX2X1 U23 ( .A(n55), .B(n55), .S0(quotient[3]), .Y(n15) );
  MX2X1 U24 ( .A(\u_div/CryTmp[8][4] ), .B(n91), .S0(quotient[8]), .Y(n16) );
  MX2X1 U25 ( .A(\u_div/CryTmp[6][4] ), .B(n92), .S0(quotient[6]), .Y(n17) );
  MX2X1 U26 ( .A(\u_div/CryTmp[5][4] ), .B(n93), .S0(quotient[5]), .Y(n18) );
  MX2X1 U27 ( .A(\u_div/CryTmp[4][4] ), .B(n94), .S0(quotient[4]), .Y(n19) );
  AND2X2 U28 ( .A(\u_div/PartRem[1][7] ), .B(n4), .Y(n20) );
  AND2X2 U29 ( .A(\u_div/PartRem[1][5] ), .B(\u_div/CryTmp[0][5] ), .Y(n21) );
  MX2X1 U30 ( .A(n1), .B(\u_div/SumTmp[8][4] ), .S0(quotient[8]), .Y(n22) );
  MX2X1 U31 ( .A(n16), .B(\u_div/SumTmp[7][4] ), .S0(quotient[7]), .Y(n23) );
  MX2X1 U32 ( .A(n7), .B(\u_div/SumTmp[6][4] ), .S0(quotient[6]), .Y(n24) );
  MX2X1 U33 ( .A(n17), .B(\u_div/SumTmp[5][4] ), .S0(quotient[5]), .Y(n25) );
  MX2X1 U34 ( .A(n19), .B(\u_div/SumTmp[3][4] ), .S0(quotient[3]), .Y(n26) );
  MX2X1 U35 ( .A(a[13]), .B(\u_div/SumTmp[9][4] ), .S0(quotient[9]), .Y(n27)
         );
  MX2X1 U36 ( .A(n18), .B(\u_div/SumTmp[4][4] ), .S0(quotient[4]), .Y(n28) );
  MX2X1 U37 ( .A(n22), .B(\u_div/SumTmp[7][5] ), .S0(quotient[7]), .Y(n29) );
  MX2X1 U38 ( .A(n23), .B(\u_div/SumTmp[6][5] ), .S0(quotient[6]), .Y(n30) );
  MX2X1 U39 ( .A(n24), .B(\u_div/SumTmp[5][5] ), .S0(quotient[5]), .Y(n31) );
  MX2X1 U40 ( .A(n31), .B(\u_div/SumTmp[4][6] ), .S0(quotient[4]), .Y(n32) );
  MX2X1 U41 ( .A(n28), .B(\u_div/SumTmp[3][5] ), .S0(quotient[3]), .Y(n33) );
  MX2X1 U42 ( .A(n27), .B(\u_div/SumTmp[8][5] ), .S0(quotient[8]), .Y(n34) );
  MX2X1 U43 ( .A(n25), .B(\u_div/SumTmp[4][5] ), .S0(quotient[4]), .Y(n35) );
  MX2X1 U44 ( .A(a[14]), .B(\u_div/SumTmp[9][5] ), .S0(quotient[9]), .Y(n36)
         );
  MX2X1 U45 ( .A(\u_div/PartRem[15][1] ), .B(\u_div/SumTmp[9][6] ), .S0(
        quotient[9]), .Y(n37) );
  MX2X1 U46 ( .A(n9), .B(\u_div/SumTmp[5][7] ), .S0(quotient[5]), .Y(n38) );
  MX2X1 U47 ( .A(n11), .B(\u_div/SumTmp[6][7] ), .S0(quotient[6]), .Y(n39) );
  MX2X1 U48 ( .A(n10), .B(\u_div/SumTmp[4][7] ), .S0(quotient[4]), .Y(n40) );
  MX2X1 U49 ( .A(n32), .B(\u_div/SumTmp[3][7] ), .S0(quotient[3]), .Y(n41) );
  MX2X1 U50 ( .A(n12), .B(\u_div/SumTmp[7][7] ), .S0(quotient[7]), .Y(n42) );
  MX2X1 U51 ( .A(n37), .B(\u_div/SumTmp[8][7] ), .S0(quotient[8]), .Y(n43) );
  MX2X1 U52 ( .A(\u_div/PartRem[16][1] ), .B(\u_div/SumTmp[9][7] ), .S0(
        quotient[9]), .Y(n44) );
  MX2X1 U53 ( .A(n84), .B(n56), .S0(quotient[1]), .Y(n45) );
  XOR2X1 U54 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/CryTmp[1][4] ), .Y(n46) );
  MX2X1 U55 ( .A(n70), .B(n70), .S0(quotient[8]), .Y(n47) );
  MX2X1 U56 ( .A(n71), .B(n71), .S0(quotient[7]), .Y(n48) );
  MX2X1 U57 ( .A(n72), .B(n72), .S0(quotient[6]), .Y(n49) );
  XNOR2X1 U58 ( .A(\u_div/PartRem[2][7] ), .B(\u_div/CryTmp[1][7] ), .Y(n50)
         );
  XNOR2X1 U59 ( .A(\u_div/PartRem[2][6] ), .B(\u_div/CryTmp[1][6] ), .Y(n51)
         );
  XNOR2X1 U60 ( .A(\u_div/PartRem[2][5] ), .B(\u_div/CryTmp[1][5] ), .Y(n52)
         );
  MX2X1 U61 ( .A(n75), .B(n75), .S0(quotient[4]), .Y(n53) );
  XNOR2X1 U62 ( .A(\u_div/PartRem[2][8] ), .B(\u_div/CryTmp[1][8] ), .Y(n54)
         );
  MX2X1 U63 ( .A(\u_div/SumTmp[4][0] ), .B(\u_div/SumTmp[4][0] ), .S0(
        quotient[4]), .Y(n55) );
  AND2X2 U64 ( .A(\u_div/CryTmp[4][9] ), .B(\u_div/PartRem[5][9] ), .Y(
        \u_div/CryTmp[4][10] ) );
  AND2X2 U65 ( .A(\u_div/CryTmp[5][9] ), .B(\u_div/PartRem[6][9] ), .Y(
        \u_div/CryTmp[5][10] ) );
  AND2X2 U66 ( .A(\u_div/CryTmp[6][9] ), .B(\u_div/PartRem[7][9] ), .Y(
        \u_div/CryTmp[6][10] ) );
  AND2X2 U67 ( .A(\u_div/CryTmp[7][9] ), .B(\u_div/PartRem[8][9] ), .Y(
        \u_div/CryTmp[7][10] ) );
  AND2X2 U68 ( .A(\u_div/CryTmp[8][9] ), .B(\u_div/PartRem[9][9] ), .Y(
        \u_div/CryTmp[8][10] ) );
  INVX1 U69 ( .A(n82), .Y(\u_div/PartRem[4][9] ) );
  XNOR2X1 U70 ( .A(\u_div/PartRem[2][9] ), .B(\u_div/CryTmp[1][9] ), .Y(n56)
         );
  XNOR2X1 U71 ( .A(\u_div/PartRem[5][9] ), .B(\u_div/CryTmp[4][9] ), .Y(n57)
         );
  OR2X2 U72 ( .A(\u_div/CryTmp[3][10] ), .B(\u_div/PartRem[4][10] ), .Y(
        quotient[3]) );
  MXI2X1 U73 ( .A(n81), .B(n57), .S0(quotient[4]), .Y(\u_div/PartRem[4][10] )
         );
  OR2X2 U74 ( .A(\u_div/CryTmp[2][10] ), .B(\u_div/PartRem[3][10] ), .Y(
        quotient[2]) );
  MXI2X1 U75 ( .A(n82), .B(n59), .S0(quotient[3]), .Y(\u_div/PartRem[3][10] )
         );
  OR2X2 U76 ( .A(\u_div/CryTmp[1][10] ), .B(\u_div/PartRem[2][10] ), .Y(
        quotient[1]) );
  MXI2X1 U77 ( .A(n83), .B(n60), .S0(quotient[2]), .Y(\u_div/PartRem[2][10] )
         );
  AND2X2 U78 ( .A(\u_div/CryTmp[4][8] ), .B(n38), .Y(\u_div/CryTmp[4][9] ) );
  AND2X2 U79 ( .A(\u_div/CryTmp[1][8] ), .B(\u_div/PartRem[2][8] ), .Y(
        \u_div/CryTmp[1][9] ) );
  MXI2X1 U80 ( .A(n38), .B(\u_div/SumTmp[4][8] ), .S0(quotient[4]), .Y(n82) );
  XOR2X1 U81 ( .A(n38), .B(\u_div/CryTmp[4][8] ), .Y(\u_div/SumTmp[4][8] ) );
  INVX1 U82 ( .A(n81), .Y(\u_div/PartRem[5][9] ) );
  INVX1 U83 ( .A(n83), .Y(\u_div/PartRem[3][9] ) );
  INVX1 U84 ( .A(n84), .Y(\u_div/PartRem[2][9] ) );
  XNOR2X1 U85 ( .A(\u_div/PartRem[6][9] ), .B(\u_div/CryTmp[5][9] ), .Y(n58)
         );
  XNOR2X1 U86 ( .A(\u_div/PartRem[4][9] ), .B(\u_div/CryTmp[3][9] ), .Y(n59)
         );
  XNOR2X1 U87 ( .A(\u_div/PartRem[3][9] ), .B(\u_div/CryTmp[2][9] ), .Y(n60)
         );
  MX2X1 U88 ( .A(n80), .B(n58), .S0(quotient[5]), .Y(n61) );
  AND2X2 U89 ( .A(\u_div/CryTmp[5][7] ), .B(n9), .Y(\u_div/CryTmp[5][8] ) );
  AND2X2 U90 ( .A(\u_div/CryTmp[5][8] ), .B(n39), .Y(\u_div/CryTmp[5][9] ) );
  AND2X2 U91 ( .A(\u_div/CryTmp[4][7] ), .B(n10), .Y(\u_div/CryTmp[4][8] ) );
  AND2X2 U92 ( .A(\u_div/CryTmp[3][8] ), .B(n40), .Y(\u_div/CryTmp[3][9] ) );
  AND2X2 U93 ( .A(\u_div/CryTmp[2][8] ), .B(n41), .Y(\u_div/CryTmp[2][9] ) );
  AND2X2 U94 ( .A(\u_div/CryTmp[1][7] ), .B(\u_div/PartRem[2][7] ), .Y(
        \u_div/CryTmp[1][8] ) );
  NAND2BX1 U95 ( .AN(n5), .B(n45), .Y(quotient[0]) );
  MXI2X1 U96 ( .A(n39), .B(\u_div/SumTmp[5][8] ), .S0(quotient[5]), .Y(n81) );
  XOR2X1 U97 ( .A(n39), .B(\u_div/CryTmp[5][8] ), .Y(\u_div/SumTmp[5][8] ) );
  MXI2X1 U98 ( .A(n40), .B(\u_div/SumTmp[3][8] ), .S0(quotient[3]), .Y(n83) );
  XOR2X1 U99 ( .A(n40), .B(\u_div/CryTmp[3][8] ), .Y(\u_div/SumTmp[3][8] ) );
  MXI2X1 U100 ( .A(n41), .B(\u_div/SumTmp[2][8] ), .S0(quotient[2]), .Y(n84)
         );
  XOR2X1 U101 ( .A(n41), .B(\u_div/CryTmp[2][8] ), .Y(\u_div/SumTmp[2][8] ) );
  XOR2X1 U102 ( .A(n9), .B(\u_div/CryTmp[5][7] ), .Y(\u_div/SumTmp[5][7] ) );
  XOR2X1 U103 ( .A(n10), .B(\u_div/CryTmp[4][7] ), .Y(\u_div/SumTmp[4][7] ) );
  INVX1 U104 ( .A(n80), .Y(\u_div/PartRem[6][9] ) );
  INVX1 U105 ( .A(n85), .Y(\u_div/PartRem[2][8] ) );
  XNOR2X1 U106 ( .A(\u_div/PartRem[7][9] ), .B(\u_div/CryTmp[6][9] ), .Y(n62)
         );
  MX2X1 U107 ( .A(n79), .B(n62), .S0(quotient[6]), .Y(n63) );
  AND2X2 U108 ( .A(\u_div/CryTmp[6][6] ), .B(n29), .Y(\u_div/CryTmp[6][7] ) );
  AND2X2 U109 ( .A(\u_div/CryTmp[6][7] ), .B(n11), .Y(\u_div/CryTmp[6][8] ) );
  AND2X2 U110 ( .A(\u_div/CryTmp[6][8] ), .B(n42), .Y(\u_div/CryTmp[6][9] ) );
  AND2X2 U111 ( .A(\u_div/CryTmp[5][6] ), .B(n30), .Y(\u_div/CryTmp[5][7] ) );
  AND2X2 U112 ( .A(\u_div/CryTmp[4][6] ), .B(n31), .Y(\u_div/CryTmp[4][7] ) );
  AND2X2 U113 ( .A(\u_div/CryTmp[3][7] ), .B(n32), .Y(\u_div/CryTmp[3][8] ) );
  AND2X2 U114 ( .A(\u_div/CryTmp[2][7] ), .B(n8), .Y(\u_div/CryTmp[2][8] ) );
  AND2X2 U115 ( .A(\u_div/CryTmp[1][6] ), .B(\u_div/PartRem[2][6] ), .Y(
        \u_div/CryTmp[1][7] ) );
  MXI2X1 U116 ( .A(n85), .B(n54), .S0(quotient[1]), .Y(\u_div/PartRem[1][9] )
         );
  MXI2X1 U117 ( .A(n42), .B(\u_div/SumTmp[6][8] ), .S0(quotient[6]), .Y(n80)
         );
  XOR2X1 U118 ( .A(n42), .B(\u_div/CryTmp[6][8] ), .Y(\u_div/SumTmp[6][8] ) );
  MXI2X1 U119 ( .A(n8), .B(\u_div/SumTmp[2][7] ), .S0(quotient[2]), .Y(n85) );
  XOR2X1 U120 ( .A(n8), .B(\u_div/CryTmp[2][7] ), .Y(\u_div/SumTmp[2][7] ) );
  XOR2X1 U121 ( .A(n29), .B(\u_div/CryTmp[6][6] ), .Y(\u_div/SumTmp[6][6] ) );
  XOR2X1 U122 ( .A(n11), .B(\u_div/CryTmp[6][7] ), .Y(\u_div/SumTmp[6][7] ) );
  XOR2X1 U123 ( .A(n30), .B(\u_div/CryTmp[5][6] ), .Y(\u_div/SumTmp[5][6] ) );
  XOR2X1 U124 ( .A(n31), .B(\u_div/CryTmp[4][6] ), .Y(\u_div/SumTmp[4][6] ) );
  XOR2X1 U125 ( .A(n32), .B(\u_div/CryTmp[3][7] ), .Y(\u_div/SumTmp[3][7] ) );
  INVX1 U126 ( .A(n79), .Y(\u_div/PartRem[7][9] ) );
  INVX1 U127 ( .A(n86), .Y(\u_div/PartRem[2][7] ) );
  XNOR2X1 U128 ( .A(\u_div/PartRem[8][9] ), .B(\u_div/CryTmp[7][9] ), .Y(n64)
         );
  MX2X1 U129 ( .A(n78), .B(n64), .S0(quotient[7]), .Y(n65) );
  AND2X2 U130 ( .A(\u_div/CryTmp[8][6] ), .B(n36), .Y(\u_div/CryTmp[8][7] ) );
  AND2X2 U131 ( .A(\u_div/CryTmp[8][7] ), .B(n37), .Y(\u_div/CryTmp[8][8] ) );
  AND2X2 U132 ( .A(\u_div/CryTmp[7][5] ), .B(n22), .Y(\u_div/CryTmp[7][6] ) );
  AND2X2 U133 ( .A(\u_div/CryTmp[7][6] ), .B(n34), .Y(\u_div/CryTmp[7][7] ) );
  AND2X2 U134 ( .A(\u_div/CryTmp[7][7] ), .B(n12), .Y(\u_div/CryTmp[7][8] ) );
  AND2X2 U135 ( .A(\u_div/CryTmp[7][8] ), .B(n43), .Y(\u_div/CryTmp[7][9] ) );
  AND2X2 U136 ( .A(\u_div/CryTmp[6][5] ), .B(n23), .Y(\u_div/CryTmp[6][6] ) );
  AND2X2 U137 ( .A(\u_div/CryTmp[5][5] ), .B(n24), .Y(\u_div/CryTmp[5][6] ) );
  AND2X2 U138 ( .A(\u_div/CryTmp[4][5] ), .B(n25), .Y(\u_div/CryTmp[4][6] ) );
  AND2X2 U139 ( .A(\u_div/CryTmp[3][6] ), .B(n35), .Y(\u_div/CryTmp[3][7] ) );
  AND2X2 U140 ( .A(\u_div/CryTmp[2][6] ), .B(n33), .Y(\u_div/CryTmp[2][7] ) );
  AND2X2 U141 ( .A(\u_div/CryTmp[1][5] ), .B(\u_div/PartRem[2][5] ), .Y(
        \u_div/CryTmp[1][6] ) );
  MXI2X1 U142 ( .A(n86), .B(n50), .S0(quotient[1]), .Y(\u_div/PartRem[1][8] )
         );
  XOR2X1 U143 ( .A(n22), .B(\u_div/CryTmp[7][5] ), .Y(\u_div/SumTmp[7][5] ) );
  XOR2X1 U144 ( .A(n23), .B(\u_div/CryTmp[6][5] ), .Y(\u_div/SumTmp[6][5] ) );
  XOR2X1 U145 ( .A(n24), .B(\u_div/CryTmp[5][5] ), .Y(\u_div/SumTmp[5][5] ) );
  XOR2X1 U146 ( .A(n25), .B(\u_div/CryTmp[4][5] ), .Y(\u_div/SumTmp[4][5] ) );
  INVX1 U147 ( .A(n87), .Y(\u_div/PartRem[2][6] ) );
  MXI2X1 U148 ( .A(n43), .B(\u_div/SumTmp[7][8] ), .S0(quotient[7]), .Y(n79)
         );
  XOR2X1 U149 ( .A(n43), .B(\u_div/CryTmp[7][8] ), .Y(\u_div/SumTmp[7][8] ) );
  MXI2X1 U150 ( .A(n33), .B(\u_div/SumTmp[2][6] ), .S0(quotient[2]), .Y(n86)
         );
  XOR2X1 U151 ( .A(n33), .B(\u_div/CryTmp[2][6] ), .Y(\u_div/SumTmp[2][6] ) );
  XOR2X1 U152 ( .A(n34), .B(\u_div/CryTmp[7][6] ), .Y(\u_div/SumTmp[7][6] ) );
  XOR2X1 U153 ( .A(n12), .B(\u_div/CryTmp[7][7] ), .Y(\u_div/SumTmp[7][7] ) );
  XOR2X1 U154 ( .A(n35), .B(\u_div/CryTmp[3][6] ), .Y(\u_div/SumTmp[3][6] ) );
  INVX1 U155 ( .A(n78), .Y(\u_div/PartRem[8][9] ) );
  XNOR2X1 U156 ( .A(\u_div/PartRem[9][9] ), .B(\u_div/CryTmp[8][9] ), .Y(n66)
         );
  MX2X1 U157 ( .A(n77), .B(n66), .S0(quotient[8]), .Y(n67) );
  AND2X2 U158 ( .A(\u_div/CryTmp[9][9] ), .B(\u_div/PartRem[18][1] ), .Y(
        quotient[9]) );
  INVX1 U159 ( .A(n89), .Y(\u_div/PartRem[2][4] ) );
  AND2X2 U160 ( .A(\u_div/CryTmp[8][5] ), .B(n27), .Y(\u_div/CryTmp[8][6] ) );
  AND2X2 U161 ( .A(\u_div/CryTmp[8][8] ), .B(n44), .Y(\u_div/CryTmp[8][9] ) );
  AND2X2 U162 ( .A(\u_div/CryTmp[3][5] ), .B(n28), .Y(\u_div/CryTmp[3][6] ) );
  AND2X2 U163 ( .A(\u_div/CryTmp[2][5] ), .B(n26), .Y(\u_div/CryTmp[2][6] ) );
  AND2X2 U164 ( .A(\u_div/CryTmp[9][6] ), .B(\u_div/PartRem[15][1] ), .Y(
        \u_div/CryTmp[9][7] ) );
  OR2X2 U165 ( .A(\u_div/CryTmp[8][4] ), .B(n1), .Y(\u_div/CryTmp[8][5] ) );
  OR2X2 U166 ( .A(\u_div/CryTmp[7][4] ), .B(n16), .Y(\u_div/CryTmp[7][5] ) );
  OR2X2 U167 ( .A(\u_div/CryTmp[6][4] ), .B(n7), .Y(\u_div/CryTmp[6][5] ) );
  OR2X2 U168 ( .A(\u_div/CryTmp[5][4] ), .B(n17), .Y(\u_div/CryTmp[5][5] ) );
  OR2X2 U169 ( .A(\u_div/CryTmp[4][4] ), .B(n18), .Y(\u_div/CryTmp[4][5] ) );
  OR2X2 U170 ( .A(\u_div/CryTmp[1][4] ), .B(\u_div/PartRem[2][4] ), .Y(
        \u_div/CryTmp[1][5] ) );
  MXI2X1 U171 ( .A(n87), .B(n51), .S0(quotient[1]), .Y(\u_div/PartRem[1][7] )
         );
  MXI2X1 U172 ( .A(n26), .B(\u_div/SumTmp[2][5] ), .S0(quotient[2]), .Y(n87)
         );
  XOR2X1 U173 ( .A(n26), .B(\u_div/CryTmp[2][5] ), .Y(\u_div/SumTmp[2][5] ) );
  XNOR2X1 U174 ( .A(n1), .B(\u_div/CryTmp[8][4] ), .Y(\u_div/SumTmp[8][4] ) );
  XOR2X1 U175 ( .A(n27), .B(\u_div/CryTmp[8][5] ), .Y(\u_div/SumTmp[8][5] ) );
  XNOR2X1 U176 ( .A(n16), .B(\u_div/CryTmp[7][4] ), .Y(\u_div/SumTmp[7][4] )
         );
  XNOR2X1 U177 ( .A(n7), .B(\u_div/CryTmp[6][4] ), .Y(\u_div/SumTmp[6][4] ) );
  XNOR2X1 U178 ( .A(n17), .B(\u_div/CryTmp[5][4] ), .Y(\u_div/SumTmp[5][4] )
         );
  XNOR2X1 U179 ( .A(n18), .B(\u_div/CryTmp[4][4] ), .Y(\u_div/SumTmp[4][4] )
         );
  XOR2X1 U180 ( .A(n28), .B(\u_div/CryTmp[3][5] ), .Y(\u_div/SumTmp[3][5] ) );
  XOR2X1 U181 ( .A(a[14]), .B(\u_div/CryTmp[9][5] ), .Y(\u_div/SumTmp[9][5] )
         );
  INVX1 U182 ( .A(n88), .Y(\u_div/PartRem[2][5] ) );
  AND2X2 U183 ( .A(\u_div/CryTmp[9][5] ), .B(a[14]), .Y(\u_div/CryTmp[9][6] )
         );
  MXI2X1 U184 ( .A(n44), .B(\u_div/SumTmp[8][8] ), .S0(quotient[8]), .Y(n78)
         );
  XOR2X1 U185 ( .A(n44), .B(\u_div/CryTmp[8][8] ), .Y(\u_div/SumTmp[8][8] ) );
  XOR2X1 U186 ( .A(n36), .B(\u_div/CryTmp[8][6] ), .Y(\u_div/SumTmp[8][6] ) );
  XOR2X1 U187 ( .A(n37), .B(\u_div/CryTmp[8][7] ), .Y(\u_div/SumTmp[8][7] ) );
  XOR2X1 U188 ( .A(\u_div/PartRem[15][1] ), .B(\u_div/CryTmp[9][6] ), .Y(
        \u_div/SumTmp[9][6] ) );
  INVX1 U189 ( .A(n77), .Y(\u_div/PartRem[9][9] ) );
  XNOR2X1 U190 ( .A(\u_div/PartRem[18][1] ), .B(\u_div/CryTmp[9][9] ), .Y(n68)
         );
  MX2X1 U191 ( .A(n98), .B(n68), .S0(quotient[9]), .Y(n69) );
  MXI2X1 U192 ( .A(\u_div/CryTmp[2][4] ), .B(n96), .S0(quotient[2]), .Y(n89)
         );
  INVX1 U193 ( .A(n97), .Y(\u_div/CryTmp[7][4] ) );
  MXI2X1 U194 ( .A(n13), .B(n13), .S0(quotient[8]), .Y(n97) );
  INVX1 U195 ( .A(n92), .Y(\u_div/CryTmp[6][4] ) );
  MXI2X1 U196 ( .A(n47), .B(n47), .S0(quotient[7]), .Y(n92) );
  INVX1 U197 ( .A(n93), .Y(\u_div/CryTmp[5][4] ) );
  MXI2X1 U198 ( .A(n48), .B(n48), .S0(quotient[6]), .Y(n93) );
  INVX1 U199 ( .A(n94), .Y(\u_div/CryTmp[4][4] ) );
  MXI2X1 U200 ( .A(n49), .B(n49), .S0(quotient[5]), .Y(n94) );
  INVX1 U201 ( .A(n91), .Y(\u_div/CryTmp[8][4] ) );
  MXI2X1 U202 ( .A(a[11]), .B(a[11]), .S0(quotient[9]), .Y(n91) );
  INVX1 U203 ( .A(n90), .Y(\u_div/CryTmp[1][4] ) );
  AND2X2 U204 ( .A(\u_div/CryTmp[9][7] ), .B(\u_div/PartRem[16][1] ), .Y(
        \u_div/CryTmp[9][8] ) );
  AND2X2 U205 ( .A(\u_div/CryTmp[9][8] ), .B(\u_div/PartRem[17][1] ), .Y(
        \u_div/CryTmp[9][9] ) );
  OR2X2 U206 ( .A(\u_div/CryTmp[3][4] ), .B(n19), .Y(\u_div/CryTmp[3][5] ) );
  OR2X2 U207 ( .A(\u_div/CryTmp[2][4] ), .B(n6), .Y(\u_div/CryTmp[2][5] ) );
  MXI2X1 U208 ( .A(n88), .B(n52), .S0(quotient[1]), .Y(\u_div/PartRem[1][6] )
         );
  MXI2X1 U209 ( .A(n6), .B(\u_div/SumTmp[2][4] ), .S0(quotient[2]), .Y(n88) );
  XNOR2X1 U210 ( .A(n6), .B(\u_div/CryTmp[2][4] ), .Y(\u_div/SumTmp[2][4] ) );
  XNOR2X1 U211 ( .A(n19), .B(\u_div/CryTmp[3][4] ), .Y(\u_div/SumTmp[3][4] )
         );
  XNOR2X1 U212 ( .A(a[13]), .B(a[12]), .Y(\u_div/SumTmp[9][4] ) );
  OR2X2 U213 ( .A(a[12]), .B(a[13]), .Y(\u_div/CryTmp[9][5] ) );
  MXI2X1 U214 ( .A(\u_div/PartRem[17][1] ), .B(\u_div/SumTmp[9][8] ), .S0(
        quotient[9]), .Y(n77) );
  XOR2X1 U215 ( .A(\u_div/PartRem[17][1] ), .B(\u_div/CryTmp[9][8] ), .Y(
        \u_div/SumTmp[9][8] ) );
  XOR2X1 U216 ( .A(\u_div/PartRem[16][1] ), .B(\u_div/CryTmp[9][7] ), .Y(
        \u_div/SumTmp[9][7] ) );
  MXI2X1 U217 ( .A(n15), .B(n15), .S0(quotient[2]), .Y(n90) );
  INVX1 U218 ( .A(n95), .Y(\u_div/CryTmp[3][4] ) );
  MXI2X1 U219 ( .A(n14), .B(n14), .S0(quotient[4]), .Y(n95) );
  INVX1 U220 ( .A(n96), .Y(\u_div/CryTmp[2][4] ) );
  MXI2X1 U221 ( .A(n53), .B(n53), .S0(quotient[3]), .Y(n96) );
  MXI2X1 U222 ( .A(n89), .B(n46), .S0(quotient[1]), .Y(\u_div/PartRem[1][5] )
         );
  NAND2BX1 U223 ( .AN(\u_div/CryTmp[0][4] ), .B(n2), .Y(\u_div/CryTmp[0][5] )
         );
  INVX1 U224 ( .A(a[12]), .Y(n99) );
  MX2X1 U225 ( .A(\u_div/SumTmp[9][0] ), .B(\u_div/SumTmp[9][0] ), .S0(
        quotient[9]), .Y(n70) );
  MX2X1 U226 ( .A(\u_div/SumTmp[8][0] ), .B(\u_div/SumTmp[8][0] ), .S0(
        quotient[8]), .Y(n71) );
  MX2X1 U227 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[7][0] ), .S0(
        quotient[7]), .Y(n72) );
  MX2X1 U228 ( .A(n73), .B(n73), .S0(quotient[1]), .Y(\u_div/CryTmp[0][4] ) );
  MX2X1 U229 ( .A(n76), .B(n76), .S0(quotient[2]), .Y(n73) );
  MX2X1 U230 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[6][0] ), .S0(
        quotient[6]), .Y(n74) );
  MX2X1 U231 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[5][0] ), .S0(
        quotient[5]), .Y(n75) );
  INVX1 U232 ( .A(\u_div/PartRem[18][1] ), .Y(n98) );
  MX2X1 U233 ( .A(\u_div/SumTmp[3][0] ), .B(\u_div/SumTmp[3][0] ), .S0(
        quotient[3]), .Y(n76) );
endmodule


module Equation_Implementation ( Im_block, Ready, W_block, clk, ena_in, params, 
        rst, block_done, block_out, M2 );
  input [31:0] Im_block;
  input [31:0] W_block;
  input [46:0] params;
  output [31:0] block_out;
  output [19:0] M2;
  input Ready, clk, ena_in, rst;
  output block_done;
  wire   sums_done, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N214, N215, N216, N217, N218, N219, N220, N238, N239,
         N240, N241, N242, N243, N244, N245, N250, N251, N253, N255, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306,
         N307, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N394, N395, N396, N397, N398, N399, N400, N401,
         N402, N403, N404, N405, eq345_done, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N509, N510, N511, N512, N513, N514, N515,
         N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526,
         N527, N528, N529, N530, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, N568, N569, N570, N571, N572, eq12_done, N635,
         N636, N637, N638, N639, N640, N641, N642, N643, N644, N645, N646,
         N647, N648, N649, N650, N651, N652, N653, N654, N655, N656, N657,
         N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, N668,
         N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679,
         N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, N690,
         N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701,
         N702, N703, N704, N705, N706, N707, N708, N709, N710, N711, N712,
         N713, N714, N715, N716, N717, N718, N719, N720, N721, N722, N723,
         N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734,
         N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745,
         N746, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N871, N918,
         N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929,
         N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940,
         N941, N942, N943, N958, N959, N960, N961, N962, N963, N964, N965,
         N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011,
         N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021,
         N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1075,
         N1076, N1156, n268, n270, n271, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, N390, N389,
         N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378,
         N377, N376, N375, N374, N373, N372, N371, N370, N366, N365, N364,
         N363, N362, N361, N360, N359, N345, N344, N343, N342, N341, N340,
         N339, N338, N337, N336, N335, N334, N295, N294, N293, N292, N291,
         N290, N289, N288, N287, N286, N285, N284, N283, N279, N278, N277,
         N276, N275, N274, N273, N272, N590, N589, N588, N587, N586, N585,
         N584, N583, N582, N999, N998, N997, N996, N995, N994, N993, N992,
         N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981,
         N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970,
         N969, N968, N967, N966, N1001, N1000, N178, N177, N176, N175, N174,
         N173, N172, N171, N170, N149, N148, N147, N146, N145, N144, N143,
         N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N1159,
         N1158, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908,
         N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897,
         N896, N895, N894, N893, N892, N891, N890, N889, N756, N755, N754,
         N753, N752, N751, N750, N749, N748, N806, N805, N804, N803, N802,
         N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791,
         N789, N788, N786, N785, N784, N783, N782, N781, N780, N779, N778,
         N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767,
         N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N630,
         N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N597,
         N596, N595, N594, N593, \mult_134_2/n38 , \mult_134_2/n37 ,
         \mult_134_2/n36 , \mult_134_2/n35 , \mult_134_2/n34 ,
         \mult_134_2/n33 , \sub_1_root_sub_0_root_add_81_6/carry[8] ,
         \sub_1_root_sub_0_root_add_81_6/carry[7] ,
         \sub_1_root_sub_0_root_add_81_6/carry[6] ,
         \sub_1_root_sub_0_root_add_81_6/carry[5] ,
         \sub_1_root_sub_0_root_add_81_6/carry[4] ,
         \sub_1_root_sub_0_root_add_81_6/carry[3] ,
         \sub_1_root_sub_0_root_add_81_6/carry[2] , \sub_136_2/carry[10] ,
         \sub_136_2/carry[7] , \sub_136_2/carry[6] , \sub_136_2/carry[5] ,
         \sub_136_2/carry[3] , \sub_136_2/carry[2] ,
         \sub_2_root_sub_0_root_sub_81_2/carry[8] ,
         \sub_2_root_sub_0_root_sub_81_2/carry[7] ,
         \sub_2_root_sub_0_root_sub_81_2/carry[6] ,
         \sub_2_root_sub_0_root_sub_81_2/carry[5] ,
         \sub_2_root_sub_0_root_sub_81_2/carry[4] ,
         \sub_2_root_sub_0_root_sub_81_2/carry[3] ,
         \sub_2_root_sub_0_root_sub_81_2/carry[2] ,
         \sub_2_root_sub_0_root_sub_81_2/carry[1] , \mult_136/n6 ,
         \mult_136/n5 , \mult_136/n4 , \mult_136/n3 , \mult_136/n2 ,
         \mult_134/n6 , \mult_134/n5 , \mult_134/n4 , \mult_134/n3 ,
         \mult_134/n2 , \mult_134/n1 , n1, n2, n3, n4, n5, n7, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214;
  wire   [2:0] i;
  wire   [11:0] sum4;
  wire   [2:0] endOfRow;
  wire   [11:0] sum5;
  wire   [11:0] sum3;
  wire   [9:0] Mu;
  wire   [9:0] Sigma;
  wire   [8:0] G;
  wire   [9:0] pow;
  wire   [9:0] alpha;
  wire   [9:0] beta;
  wire   [2:0] i_res;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165;
  assign M2[19] = 1'b0;
  assign M2[18] = 1'b0;
  assign M2[17] = 1'b0;
  assign M2[16] = 1'b0;
  assign M2[15] = 1'b0;
  assign M2[14] = 1'b0;
  assign M2[13] = 1'b0;
  assign M2[12] = 1'b0;
  assign M2[11] = 1'b0;
  assign M2[10] = 1'b0;
  assign M2[9] = 1'b0;
  assign M2[8] = 1'b0;
  assign M2[7] = 1'b0;
  assign M2[6] = 1'b0;
  assign M2[5] = 1'b0;
  assign M2[4] = 1'b0;
  assign M2[3] = 1'b0;
  assign N583 = params[22];
  assign N582 = params[21];
  assign N749 = params[36];
  assign N748 = params[35];

  NOR3X4 U251 ( .A(n422), .B(n417), .C(n421), .Y(n402) );
  NOR3X4 U287 ( .A(i[1]), .B(i[2]), .C(i[0]), .Y(n429) );
  NOR3X4 U331 ( .A(i[0]), .B(i[1]), .C(n211), .Y(n454) );
  Power2 pow2 ( .Mu(Mu), .pow({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, pow[7:5], SYNOPSYS_UNCONNECTED__2, pow[3:1], 
        N796}) );
  Equation_Implementation_DW_div_uns_5 div_111 ( .a(sum5), .b(params[10:8]), 
        .quotient({SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, N572, N571, N570, N569, N568, N567, N566, 
        N565, N564}) );
  Equation_Implementation_DW01_sub_0 sub_0_root_sub_81_3 ( .A({N271, N270, 
        N269, N268, N267, N266, N265, N264, N263, N262, N261, N260}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, N245, N244, N243, N242, N241, N240, N239, N238}), 
        .CI(1'b0), .DIFF({N332, N331, N330, N329, N328, N327, N326, N325, N324, 
        N323, N322, N321}) );
  Equation_Implementation_DW01_add_141 add_68 ( .A(sum3), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N366, N365, N364, N363, N362, N361, N360, N359}), .CI(1'b0), 
        .SUM({N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, 
        N111}) );
  Equation_Implementation_DW01_add_142 r594 ( .A(sum5), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N220, N219, N218, N217, N216, N215, N214, N382}), .CI(1'b0), 
        .SUM({N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, 
        N260}) );
  Equation_Implementation_DW01_inc_0 r580 ( .A({1'b0, params[7:0]}), .SUM({
        N130, N129, N128, N127, N126, N125, N124, N123, N500}) );
  Equation_Implementation_DW01_sub_6 sub_3_root_sub_0_root_add_81_6 ( .A(sum5), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N245, N244, N243, N242, N241, N240, N239, 
        N238}), .CI(1'b0), .DIFF({N381, N380, N379, N378, N377, N376, N375, 
        N374, N373, N372, N371, N370}) );
  Equation_Implementation_DW01_add_148 add_0_root_sub_0_root_add_81_6 ( .A({
        N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370}), .B({n5, n5, n5, N390, N389, N388, N387, N386, N385, N384, N383, N382}), 
        .CI(1'b0), .SUM({N405, N404, N403, N402, N401, N400, N399, N398, N397, 
        N396, N395, N394}) );
  Equation_Implementation_DW01_add_147 add_1_root_sub_0_root_add_81_4 ( .A(
        sum5), .B({1'b0, 1'b0, 1'b0, 1'b0, N245, N244, N243, N242, N241, N240, 
        N239, N238}), .CI(1'b0), .SUM({N345, N344, N343, N342, N341, N340, 
        N339, N338, N337, N336, N335, N334}) );
  Equation_Implementation_DW01_sub_4 sub_0_root_sub_0_root_add_81_4 ( .A({N345, 
        N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N220, N219, N218, N217, N216, N215, N214, 
        N382}), .CI(1'b0), .DIFF({N357, N356, N355, N354, N353, N352, N351, 
        N350, N349, N348, N347, N346}) );
  Equation_Implementation_DW01_sub_9 sub_1_root_sub_0_root_sub_81_2 ( .A({N271, 
        N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N366, N365, N364, N363, N362, N361, N360, 
        N359}), .CI(1'b0), .DIFF({N295, N294, N293, N292, N291, N290, N289, 
        N288, N287, N286, N285, N284}) );
  Equation_Implementation_DW01_add_150 add_0_root_sub_0_root_sub_81_2 ( .A({
        N283, N283, N283, N283, N279, N278, N277, N276, N275, N274, N273, N272}), .B({N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284}), .CI(1'b0), .SUM({N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, 
        N297, N296}) );
  Equation_Implementation_DW01_add_152 add_134 ( .A({N590, N589, N588, N587, 
        N586, N585, N584, N583, N582, 1'b0}), .B({N736, N735, N734, N733, N732, 
        N731, N730, N729, N728, N727}), .CI(1'b0), .SUM({N746, N745, N744, 
        N743, N742, N741, N740, N739, N738, N737}) );
  Equation_Implementation_DW_mult_uns_5 mult_158_6 ( .a(alpha), .b({n183, n185, 
        n187, n189, n191, n193, n195, n197}), .product({N983, N982, N981, N980, 
        N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, 
        N967, N966}) );
  Equation_Implementation_DW_mult_uns_4 mult_158_8 ( .a(beta), .b({N965, N964, 
        N963, N962, N961, N960, N959, N958}), .product({N1001, N1000, N999, 
        N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, 
        N986, N985, N984}) );
  Equation_Implementation_DW01_add_143 add_158_2 ( .A({1'b0, N983, N982, N981, 
        N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, 
        N968, N967, N966}), .B({1'b0, N1001, N1000, N999, N998, N997, N996, 
        N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984}), .CI(1'b0), .SUM({N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, 
        N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, 
        N1002}) );
  Equation_Implementation_DW01_inc_1 r582 ( .A({1'b0, params[7:0]}), .SUM({
        N140, N139, N138, N137, N136, N135, N134, N133, 
        SYNOPSYS_UNCONNECTED__6}) );
  Equation_Implementation_DW01_sub_3 sub_72 ( .A({1'b0, N140, N139, N138, N137, 
        N136, N135, N134, N133}), .B({1'b0, N366, N365, N364, N363, N362, N361, 
        N360, N359}), .CI(1'b0), .DIFF({N149, N148, N147, N146, N145, N144, 
        N143, N142, N141}) );
  Equation_Implementation_DW01_add_146 add_72_3 ( .A(sum4), .B({N149, N149, 
        N149, N149, N148, N147, N146, N145, N144, N143, N142, N141}), .CI(1'b0), .SUM({N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150}) );
  Equation_Implementation_DW01_sub_2 sub_72_2 ( .A({1'b0, N366, N365, N364, 
        N363, N362, N361, N360, N359}), .B({1'b0, N140, N139, N138, N137, N136, 
        N135, N134, N133}), .CI(1'b0), .DIFF({N178, N177, N176, N175, N174, 
        N173, N172, N171, N170}) );
  Equation_Implementation_DW01_add_145 add_72_5 ( .A(sum4), .B({N178, N178, 
        N178, N178, N177, N176, N175, N174, N173, N172, N171, N170}), .CI(1'b0), .SUM({N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179}) );
  Equation_Implementation_DW_mult_uns_7 mult_158_2 ( .a(params[34:28]), .b({
        n183, n185, n187, n189, n191, n193, n195, n197}), .product({N903, N902, 
        N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, 
        N889}) );
  Equation_Implementation_DW_mult_uns_6 mult_158_4 ( .a({params[40:37], N749, 
        N748}), .b({N965, N964, N963, N962, N961, N960, N959, N958}), 
        .product({N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, 
        N907, N906, N905, N904}) );
  Equation_Implementation_DW01_add_144 add_158 ( .A({1'b0, N903, N902, N901, 
        N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889}), .B({1'b0, 1'b0, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, 
        N907, N906, N905, N904}), .CI(1'b0), .SUM({N933, N932, N931, N930, 
        N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918}) );
  Equation_Implementation_DW01_add_151 add_136 ( .A({N756, N755, N754, N753, 
        N752, N751, N750, N749, N748, 1'b0}), .B({N848, N847, N846, N845, N844, 
        N843, N842, N841, N840, N839}), .CI(1'b0), .SUM({N858, N857, N856, 
        N855, N854, N853, N852, N851, N850, N849}) );
  Equation_Implementation_DW_mult_uns_12 mult_134_4 ( .a({N694, N693, N692, 
        N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, 
        N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, 
        N667, N666, N665, N664, N663}), .b({1'b1, 1'b1, pow[7:5], 1'b0, 
        pow[3:1], n48}), .product({SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, N726, N725, N724, N723, N722, N721, N720, 
        N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, 
        N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, 
        N695}) );
  Equation_Implementation_DW01_sub_8 sub_136 ( .A({1'b0, params[46:41]}), .B({
        1'b0, params[40:37], N749, N748}), .CI(1'b0), .DIFF({N763, N762, N761, 
        N760, N759, N758, N757}) );
  Equation_Implementation_DW_mult_uns_10 mult_136_2 ( .a({N763, N763, N763, 
        N763, N763, N763, N763, N763, N763, N763, N763, N763, N763, N763, N763, 
        N763, N763, N763, N763, N763, N763, N763, N763, N763, N763, N763, N762, 
        N761, N760, N759, N758, N757}), .b(Sigma), .product({
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, N795, N794, N793, 
        N792, N791, SYNOPSYS_UNCONNECTED__27, N789, N788, 
        SYNOPSYS_UNCONNECTED__28, N786, N785, N784, N783, N782, N781, N780, 
        N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, 
        N767, N766, N765, N764}) );
  Equation_Implementation_DW_mult_uns_9 mult_136_3 ( .a({N795, N794, n38, N792, 
        N791, n45, N789, N788, n40, N786, N785, n43, N783, N782, n41, N780, 
        N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, 
        N767, N766, N765, N764}), .b({N806, N806, N806, N806, N806, N806, N806, 
        N806, N806, N806, N806, N806, N806, N806, N806, N806, N806, N806, N806, 
        N806, N806, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, 
        n48}), .product({SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, N838, N837, N836, 
        N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, 
        N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, 
        N811, N810, N809, N808, N807}) );
  Equation_Implementation_DW01_sub_1 sub_134 ( .A({1'b0, params[34:28]}), .B({
        1'b0, params[27:23], N583, N582}), .CI(1'b0), .DIFF({N630, N597, N596, 
        N595, N594, N593, N601, N600}) );
  Equation_Implementation_DW_mult_uns_3 mult_109 ( .a(sum3), .b({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0}), .product({N499, N498, 
        N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, 
        N485, N484, N483, N482, N481, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63}) );
  Equation_Implementation_DW_mult_uns_2 mult_110_2 ( .a({sum4, 1'b0}), .b({
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0}), 
        .product({N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, 
        N543, N542, N541, N540, N539, N538, N537, N536, N535, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67}) );
  Equation_Implementation_DW_mult_uns_0 mult_134_3 ( .a({n12, n12, n12, n12, 
        n12, n12, n12, n12, n12, n12, n12, n12, n12, n12, n12, n12, n12, n12, 
        n12, n12, n12, N609, N608, N607, N606, N605, N604, N603, N602, N601, 
        N600, 1'b0}), .b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 
        1'b0}), .product({SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, N662, N661, N660, 
        N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, 
        N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, 
        N635, SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81}) );
  Equation_Implementation_DW_mult_uns_8 mult_109_2 ( .a(params[10:8]), .b({
        N130, N129, N128, N127, N126, N125, N124, N123, N500}), .product({N520, 
        N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509}) );
  ADDFX2 \mult_134_2/U49  ( .A(N594), .B(N601), .CI(\mult_134_2/n38 ), .CO(
        \mult_134_2/n37 ), .S(N603) );
  ADDFX2 \mult_134_2/U48  ( .A(N595), .B(N593), .CI(\mult_134_2/n37 ), .CO(
        \mult_134_2/n36 ), .S(N604) );
  ADDFX2 \mult_134_2/U47  ( .A(N596), .B(N594), .CI(\mult_134_2/n36 ), .CO(
        \mult_134_2/n35 ), .S(N605) );
  ADDFX2 \mult_134_2/U46  ( .A(N597), .B(N595), .CI(\mult_134_2/n35 ), .CO(
        \mult_134_2/n34 ), .S(N606) );
  ADDFX2 \mult_134_2/U45  ( .A(N596), .B(n12), .CI(\mult_134_2/n34 ), .CO(
        \mult_134_2/n33 ), .S(N607) );
  ADDFX2 \mult_134_2/U44  ( .A(N597), .B(n12), .CI(\mult_134_2/n33 ), .CO(N609), .S(N608) );
  ADDHXL \mult_136/U7  ( .A(N748), .B(params[37]), .CO(\mult_136/n6 ), .S(N750) );
  ADDFX2 \mult_136/U6  ( .A(params[38]), .B(N749), .CI(\mult_136/n6 ), .CO(
        \mult_136/n5 ), .S(N751) );
  ADDFX2 \mult_136/U5  ( .A(params[39]), .B(params[37]), .CI(\mult_136/n5 ), 
        .CO(\mult_136/n4 ), .S(N752) );
  ADDFX2 \mult_136/U4  ( .A(params[40]), .B(params[38]), .CI(\mult_136/n4 ), 
        .CO(\mult_136/n3 ), .S(N753) );
  ADDHXL \mult_136/U3  ( .A(params[39]), .B(\mult_136/n3 ), .CO(\mult_136/n2 ), 
        .S(N754) );
  ADDHXL \mult_136/U2  ( .A(params[40]), .B(\mult_136/n2 ), .CO(N756), .S(N755) );
  ADDHXL \mult_134/U7  ( .A(N582), .B(params[23]), .CO(\mult_134/n6 ), .S(N584) );
  ADDFX2 \mult_134/U6  ( .A(params[24]), .B(N583), .CI(\mult_134/n6 ), .CO(
        \mult_134/n5 ), .S(N585) );
  ADDFX2 \mult_134/U5  ( .A(params[25]), .B(params[23]), .CI(\mult_134/n5 ), 
        .CO(\mult_134/n4 ), .S(N586) );
  ADDFX2 \mult_134/U4  ( .A(params[26]), .B(params[24]), .CI(\mult_134/n4 ), 
        .CO(\mult_134/n3 ), .S(N587) );
  ADDFX2 \mult_134/U3  ( .A(params[27]), .B(params[25]), .CI(\mult_134/n3 ), 
        .CO(\mult_134/n2 ), .S(N588) );
  ADDHXL \mult_134/U2  ( .A(params[26]), .B(\mult_134/n2 ), .CO(\mult_134/n1 ), 
        .S(N589) );
  Equation_Implementation_DW_div_uns_13 div_134 ( .a({N662, N661, N660, N659, 
        N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, 
        N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, 
        1'b0, 1'b0, 1'b0, 1'b0}), .b(Sigma), .quotient({N694, N693, N692, N691, 
        N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, 
        N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, 
        N666, N665, N664, N663}) );
  Equation_Implementation_DW_div_uns_19 div_134_2 ( .a({N726, N725, N724, N723, 
        N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, 
        N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, 
        N698, N697, N696, N695}), .b({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0, 1'b0}), .quotient({SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, N736, N735, N734, N733, N732, N731, N730, 
        N729, N728, N727}) );
  Equation_Implementation_DW_div_uns_24 div_136 ( .a({N838, N837, N836, N835, 
        N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, 
        N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, 
        N810, N809, N808, N807}), .b({1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .quotient({SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, N848, N847, N846, 
        N845, N844, N843, N842, N841, N840, N839}) );
  Equation_Implementation_DW_div_uns_29 div_109 ( .a({N499, N498, N497, N496, 
        N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, 
        N483, N482, N481, 1'b0, 1'b0, 1'b0}), .b({N520, N519, N518, N517, N516, 
        N515, N514, N513, N512, N511, N510, N509}), .quotient({
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, N530, N529, N528, 
        N527, N526, N525, N524, N523, N522, N521}) );
  Equation_Implementation_DW_div_uns_34 div_110 ( .a({N553, N552, N551, N550, 
        N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, 
        N537, N536, N535, 1'b0, 1'b0, 1'b0, 1'b0}), .b({N520, N519, N518, N517, 
        N516, N515, N514, N513, N512, N511, N510, N509}), .quotient({
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, N563, N562, N561, N560, N559, N558, N557, 
        N556, N555, N554}) );
  Equation_Implementation_DW_div_uns_46 div_158 ( .a({N933, N932, N931, N930, 
        N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918}), .b({1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .quotient({
        SYNOPSYS_UNCONNECTED__151, SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, N943, N942, N941, 
        N940, N939, N938, N937, N936, N935, N934}) );
  Equation_Implementation_DW_div_uns_52 div_158_2 ( .a({N1020, N1019, N1018, 
        N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, 
        N1007, N1006, N1005, N1004, N1003, N1002}), .b({1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0}), .quotient({
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, SYNOPSYS_UNCONNECTED__160, 
        SYNOPSYS_UNCONNECTED__161, SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, N1030, N1029, N1028, N1027, N1026, N1025, 
        N1024, N1023, N1022, N1021}) );
  DFFHQX1 eq345_done_reg ( .D(n518), .CK(clk), .Q(eq345_done) );
  DFFHQX1 \block_out_reg[31]  ( .D(n516), .CK(clk), .Q(block_out[31]) );
  DFFHQX1 \block_out_reg[30]  ( .D(n515), .CK(clk), .Q(block_out[30]) );
  DFFHQX1 \block_out_reg[29]  ( .D(n514), .CK(clk), .Q(block_out[29]) );
  DFFHQX1 \block_out_reg[28]  ( .D(n513), .CK(clk), .Q(block_out[28]) );
  DFFHQX1 \block_out_reg[27]  ( .D(n512), .CK(clk), .Q(block_out[27]) );
  DFFHQX1 \block_out_reg[26]  ( .D(n511), .CK(clk), .Q(block_out[26]) );
  DFFHQX1 \block_out_reg[25]  ( .D(n510), .CK(clk), .Q(block_out[25]) );
  DFFHQX1 \block_out_reg[24]  ( .D(n509), .CK(clk), .Q(block_out[24]) );
  DFFHQX1 \block_out_reg[15]  ( .D(n500), .CK(clk), .Q(block_out[15]) );
  DFFHQX1 \block_out_reg[14]  ( .D(n499), .CK(clk), .Q(block_out[14]) );
  DFFHQX1 \block_out_reg[13]  ( .D(n498), .CK(clk), .Q(block_out[13]) );
  DFFHQX1 \block_out_reg[12]  ( .D(n497), .CK(clk), .Q(block_out[12]) );
  DFFHQX1 \block_out_reg[11]  ( .D(n496), .CK(clk), .Q(block_out[11]) );
  DFFHQX1 \block_out_reg[10]  ( .D(n495), .CK(clk), .Q(block_out[10]) );
  DFFHQX1 \block_out_reg[9]  ( .D(n494), .CK(clk), .Q(block_out[9]) );
  DFFHQX1 \block_out_reg[8]  ( .D(n493), .CK(clk), .Q(block_out[8]) );
  DFFHQX1 \block_out_reg[23]  ( .D(n508), .CK(clk), .Q(block_out[23]) );
  DFFHQX1 \block_out_reg[22]  ( .D(n507), .CK(clk), .Q(block_out[22]) );
  DFFHQX1 \block_out_reg[21]  ( .D(n506), .CK(clk), .Q(block_out[21]) );
  DFFHQX1 \block_out_reg[20]  ( .D(n505), .CK(clk), .Q(block_out[20]) );
  DFFHQX1 \block_out_reg[19]  ( .D(n504), .CK(clk), .Q(block_out[19]) );
  DFFHQX1 \block_out_reg[18]  ( .D(n503), .CK(clk), .Q(block_out[18]) );
  DFFHQX1 \block_out_reg[17]  ( .D(n502), .CK(clk), .Q(block_out[17]) );
  DFFHQX1 \block_out_reg[16]  ( .D(n501), .CK(clk), .Q(block_out[16]) );
  DFFHQX1 \block_out_reg[7]  ( .D(n492), .CK(clk), .Q(block_out[7]) );
  DFFHQX1 \block_out_reg[6]  ( .D(n491), .CK(clk), .Q(block_out[6]) );
  DFFHQX1 \block_out_reg[5]  ( .D(n490), .CK(clk), .Q(block_out[5]) );
  DFFHQX1 \block_out_reg[4]  ( .D(n489), .CK(clk), .Q(block_out[4]) );
  DFFHQX1 \block_out_reg[3]  ( .D(n488), .CK(clk), .Q(block_out[3]) );
  DFFHQX1 \block_out_reg[2]  ( .D(n487), .CK(clk), .Q(block_out[2]) );
  DFFHQX1 \block_out_reg[1]  ( .D(n486), .CK(clk), .Q(block_out[1]) );
  DFFHQX1 \block_out_reg[0]  ( .D(n485), .CK(clk), .Q(block_out[0]) );
  DFFHQX1 sums_done_reg ( .D(n519), .CK(clk), .Q(sums_done) );
  DFFHQX1 eq12_done_reg ( .D(n517), .CK(clk), .Q(eq12_done) );
  EDFFX1 \G_reg[8]  ( .D(N572), .E(n36), .CK(clk), .Q(G[8]) );
  DFFHQX1 \M2_reg[0]  ( .D(params[8]), .CK(clk), .Q(M2[0]) );
  DFFHQX1 \M2_reg[2]  ( .D(params[10]), .CK(clk), .Q(M2[2]) );
  DFFHQX1 \M2_reg[1]  ( .D(params[9]), .CK(clk), .Q(M2[1]) );
  EDFFX1 \G_reg[7]  ( .D(N571), .E(n37), .CK(clk), .Q(G[7]) );
  DFFHQX1 block_done_reg ( .D(n549), .CK(clk), .Q(block_done) );
  EDFFX1 \G_reg[6]  ( .D(N570), .E(n36), .CK(clk), .Q(G[6]) );
  EDFFX1 \G_reg[0]  ( .D(N564), .E(n37), .CK(clk), .Q(G[0]) );
  EDFFX1 \G_reg[3]  ( .D(N567), .E(n37), .CK(clk), .Q(G[3]), .QN(n4) );
  EDFFX1 \G_reg[5]  ( .D(N569), .E(n37), .CK(clk), .QN(n3) );
  EDFFX1 \G_reg[2]  ( .D(N566), .E(n37), .CK(clk), .Q(G[2]) );
  EDFFX1 \G_reg[1]  ( .D(N565), .E(n37), .CK(clk), .Q(G[1]), .QN(n7) );
  EDFFX1 \G_reg[4]  ( .D(N568), .E(n36), .CK(clk), .Q(G[4]) );
  DFFHQX1 \endOfRow_reg[2]  ( .D(n534), .CK(clk), .Q(endOfRow[2]) );
  DFFHQX1 \endOfRow_reg[0]  ( .D(n521), .CK(clk), .Q(endOfRow[0]) );
  DFFHQX1 \endOfRow_reg[1]  ( .D(n520), .CK(clk), .Q(endOfRow[1]) );
  EDFFX1 \beta_reg[9]  ( .D(N858), .E(n14), .CK(clk), .Q(beta[9]) );
  EDFFX1 \beta_reg[8]  ( .D(N857), .E(n14), .CK(clk), .Q(beta[8]) );
  EDFFX1 \beta_reg[7]  ( .D(N856), .E(n14), .CK(clk), .Q(beta[7]) );
  EDFFX1 \alpha_reg[9]  ( .D(N746), .E(n14), .CK(clk), .Q(alpha[9]) );
  EDFFX1 \alpha_reg[8]  ( .D(N745), .E(n14), .CK(clk), .Q(alpha[8]) );
  EDFFX1 \alpha_reg[7]  ( .D(N744), .E(n14), .CK(clk), .Q(alpha[7]) );
  EDFFX1 \beta_reg[6]  ( .D(N855), .E(n14), .CK(clk), .Q(beta[6]) );
  EDFFX1 \beta_reg[5]  ( .D(N854), .E(n14), .CK(clk), .Q(beta[5]) );
  EDFFX1 \beta_reg[4]  ( .D(N853), .E(n14), .CK(clk), .Q(beta[4]) );
  EDFFX1 \beta_reg[3]  ( .D(N852), .E(n14), .CK(clk), .Q(beta[3]) );
  EDFFX1 \alpha_reg[6]  ( .D(N743), .E(n14), .CK(clk), .Q(alpha[6]) );
  EDFFX1 \alpha_reg[5]  ( .D(N742), .E(n14), .CK(clk), .Q(alpha[5]) );
  EDFFX1 \alpha_reg[4]  ( .D(N741), .E(n14), .CK(clk), .Q(alpha[4]) );
  EDFFX1 \alpha_reg[3]  ( .D(N740), .E(n14), .CK(clk), .Q(alpha[3]) );
  EDFFX1 \beta_reg[2]  ( .D(N851), .E(n14), .CK(clk), .Q(beta[2]) );
  EDFFX1 \beta_reg[1]  ( .D(N850), .E(n14), .CK(clk), .Q(beta[1]) );
  EDFFX1 \beta_reg[0]  ( .D(N849), .E(n14), .CK(clk), .Q(beta[0]) );
  EDFFX1 \alpha_reg[2]  ( .D(N739), .E(n14), .CK(clk), .Q(alpha[2]) );
  EDFFX1 \alpha_reg[1]  ( .D(N738), .E(n14), .CK(clk), .Q(alpha[1]) );
  EDFFX1 \alpha_reg[0]  ( .D(N737), .E(n14), .CK(clk), .Q(alpha[0]) );
  EDFFX1 \i_res_reg[0]  ( .D(n178), .E(n291), .CK(clk), .Q(i_res[0]), .QN(n271) );
  EDFFX1 \i_res_reg[1]  ( .D(N1075), .E(n291), .CK(clk), .Q(i_res[1]), .QN(
        n270) );
  EDFFX2 \i_res_reg[2]  ( .D(N1076), .E(n291), .CK(clk), .Q(i_res[2]), .QN(
        n268) );
  EDFFTRX1 \sum3_reg[10]  ( .RN(n18), .D(N121), .E(n24), .CK(clk), .Q(sum3[10]) );
  EDFFTRX1 \sum3_reg[11]  ( .RN(n18), .D(N122), .E(n24), .CK(clk), .Q(sum3[11]) );
  EDFFTRX1 \sum3_reg[9]  ( .RN(n18), .D(N120), .E(n24), .CK(clk), .Q(sum3[9])
         );
  EDFFTRX1 \sum3_reg[5]  ( .RN(n18), .D(N116), .E(n24), .CK(clk), .Q(sum3[5])
         );
  EDFFTRX1 \sum3_reg[6]  ( .RN(n18), .D(N117), .E(n24), .CK(clk), .Q(sum3[6])
         );
  EDFFTRX1 \sum3_reg[7]  ( .RN(n18), .D(N118), .E(n24), .CK(clk), .Q(sum3[7])
         );
  EDFFTRX1 \sum3_reg[8]  ( .RN(n18), .D(N119), .E(n24), .CK(clk), .Q(sum3[8])
         );
  EDFFTRX1 \sum3_reg[3]  ( .RN(n18), .D(N114), .E(n24), .CK(clk), .Q(sum3[3])
         );
  EDFFTRX1 \sum3_reg[4]  ( .RN(n18), .D(N115), .E(n24), .CK(clk), .Q(sum3[4])
         );
  EDFFTRX1 \sum3_reg[2]  ( .RN(n18), .D(N113), .E(n24), .CK(clk), .Q(sum3[2])
         );
  EDFFTRX2 \sum3_reg[0]  ( .RN(n18), .D(N111), .E(n24), .CK(clk), .Q(sum3[0])
         );
  DFFHQX1 \sum4_reg[10]  ( .D(n536), .CK(clk), .Q(sum4[10]) );
  EDFFX1 \Mu_reg[7]  ( .D(N528), .E(n37), .CK(clk), .Q(Mu[7]) );
  EDFFX1 \Mu_reg[9]  ( .D(N530), .E(n36), .CK(clk), .Q(Mu[9]) );
  EDFFX1 \Mu_reg[8]  ( .D(N529), .E(n36), .CK(clk), .Q(Mu[8]) );
  EDFFX1 \Mu_reg[3]  ( .D(N524), .E(n37), .CK(clk), .Q(Mu[3]) );
  EDFFX2 \Mu_reg[2]  ( .D(N523), .E(n37), .CK(clk), .Q(Mu[2]) );
  EDFFX1 \Mu_reg[0]  ( .D(N521), .E(n37), .CK(clk), .Q(Mu[0]) );
  EDFFX1 \Mu_reg[6]  ( .D(N527), .E(n37), .CK(clk), .Q(Mu[6]) );
  EDFFX1 \Mu_reg[5]  ( .D(N526), .E(n37), .CK(clk), .Q(Mu[5]) );
  EDFFX1 \Mu_reg[1]  ( .D(N522), .E(n37), .CK(clk), .Q(Mu[1]) );
  EDFFX1 \Mu_reg[4]  ( .D(N525), .E(n37), .CK(clk), .Q(Mu[4]) );
  EDFFX1 \Sigma_reg[4]  ( .D(N558), .E(n36), .CK(clk), .Q(Sigma[4]) );
  EDFFX1 \Sigma_reg[3]  ( .D(N557), .E(n36), .CK(clk), .Q(Sigma[3]) );
  EDFFX1 \Sigma_reg[1]  ( .D(N555), .E(n36), .CK(clk), .Q(Sigma[1]) );
  EDFFX1 \Sigma_reg[2]  ( .D(N556), .E(n36), .CK(clk), .Q(Sigma[2]) );
  EDFFX1 \Sigma_reg[5]  ( .D(N559), .E(n36), .CK(clk), .Q(Sigma[5]) );
  EDFFX1 \Sigma_reg[8]  ( .D(N562), .E(n36), .CK(clk), .Q(Sigma[8]) );
  EDFFX1 \Sigma_reg[6]  ( .D(N560), .E(n36), .CK(clk), .Q(Sigma[6]) );
  EDFFX1 \Sigma_reg[9]  ( .D(N563), .E(n36), .CK(clk), .Q(Sigma[9]) );
  EDFFX1 \Sigma_reg[0]  ( .D(N554), .E(n36), .CK(clk), .Q(Sigma[0]) );
  EDFFX1 \Sigma_reg[7]  ( .D(N561), .E(n36), .CK(clk), .Q(Sigma[7]) );
  DFFHQX2 \sum4_reg[0]  ( .D(n546), .CK(clk), .Q(sum4[0]) );
  DFFHQX2 \i_reg[1]  ( .D(n547), .CK(clk), .Q(i[1]) );
  DFFHQX2 \i_reg[2]  ( .D(n175), .CK(clk), .Q(i[2]) );
  DFFHQX2 \sum5_reg[10]  ( .D(n523), .CK(clk), .Q(sum5[10]) );
  DFFHQX2 \sum5_reg[9]  ( .D(n524), .CK(clk), .Q(sum5[9]) );
  DFFHQX2 \sum5_reg[8]  ( .D(n525), .CK(clk), .Q(sum5[8]) );
  DFFHQX2 \sum4_reg[1]  ( .D(n545), .CK(clk), .Q(sum4[1]) );
  DFFHQX2 \sum5_reg[0]  ( .D(n533), .CK(clk), .Q(sum5[0]) );
  DFFHQX2 \i_reg[0]  ( .D(n548), .CK(clk), .Q(i[0]) );
  DFFHQX2 \sum4_reg[4]  ( .D(n542), .CK(clk), .Q(sum4[4]) );
  DFFHQX2 \sum4_reg[3]  ( .D(n543), .CK(clk), .Q(sum4[3]) );
  DFFHQX2 \sum4_reg[9]  ( .D(n537), .CK(clk), .Q(sum4[9]) );
  DFFHQX2 \sum4_reg[8]  ( .D(n538), .CK(clk), .Q(sum4[8]) );
  DFFHQX2 \sum4_reg[2]  ( .D(n544), .CK(clk), .Q(sum4[2]) );
  DFFHQX2 \sum5_reg[1]  ( .D(n532), .CK(clk), .Q(sum5[1]) );
  DFFHQX2 \sum5_reg[2]  ( .D(n531), .CK(clk), .Q(sum5[2]) );
  DFFHQX2 \sum5_reg[3]  ( .D(n530), .CK(clk), .Q(sum5[3]) );
  DFFHQX2 \sum5_reg[4]  ( .D(n529), .CK(clk), .Q(sum5[4]) );
  DFFHQX2 \sum5_reg[5]  ( .D(n528), .CK(clk), .Q(sum5[5]) );
  DFFHQX2 \sum5_reg[6]  ( .D(n527), .CK(clk), .Q(sum5[6]) );
  DFFHQX2 \sum5_reg[7]  ( .D(n526), .CK(clk), .Q(sum5[7]) );
  DFFHQX2 \sum4_reg[7]  ( .D(n539), .CK(clk), .Q(sum4[7]) );
  DFFHQX2 \sum4_reg[6]  ( .D(n540), .CK(clk), .Q(sum4[6]) );
  DFFHQX2 \sum4_reg[5]  ( .D(n541), .CK(clk), .Q(sum4[5]) );
  DFFHQX2 \sum4_reg[11]  ( .D(n535), .CK(clk), .Q(sum4[11]) );
  DFFHQX2 \sum5_reg[11]  ( .D(n522), .CK(clk), .Q(sum5[11]) );
  EDFFTRX2 \sum3_reg[1]  ( .RN(n18), .D(N112), .E(n24), .CK(clk), .Q(sum3[1])
         );
  OR2X2 U11 ( .A(n206), .B(n176), .Y(n1) );
  INVX1 U12 ( .A(pow[2]), .Y(n52) );
  NAND2X2 U13 ( .A(n471), .B(n472), .Y(n2) );
  CMPR22X1 U14 ( .A(N600), .B(N593), .CO(\mult_134_2/n38 ), .S(N602) );
  NOR3XL U20 ( .A(i[0]), .B(i[2]), .C(n210), .Y(n431) );
  NOR3XL U25 ( .A(i[1]), .B(i[2]), .C(n209), .Y(n430) );
  CLKINVX3 U28 ( .A(\sub_136_2/carry[5] ), .Y(N800) );
  AOI22XL U29 ( .A0(N303), .A1(n28), .B0(sum5[7]), .B1(n46), .Y(n317) );
  AOI22XL U32 ( .A0(N302), .A1(n28), .B0(sum5[6]), .B1(n46), .Y(n319) );
  AOI22XL U33 ( .A0(N301), .A1(n28), .B0(sum5[5]), .B1(n46), .Y(n321) );
  AOI22XL U34 ( .A0(N300), .A1(n28), .B0(sum5[4]), .B1(n46), .Y(n323) );
  AOI22XL U35 ( .A0(N299), .A1(n28), .B0(sum5[3]), .B1(n46), .Y(n325) );
  AOI22XL U36 ( .A0(N298), .A1(n28), .B0(sum5[2]), .B1(n46), .Y(n327) );
  AOI22XL U37 ( .A0(N297), .A1(n28), .B0(sum5[1]), .B1(n46), .Y(n329) );
  AOI22XL U38 ( .A0(N307), .A1(n28), .B0(sum5[11]), .B1(n46), .Y(n304) );
  BUFX3 U39 ( .A(n284), .Y(n22) );
  BUFX3 U40 ( .A(n286), .Y(n23) );
  BUFX3 U41 ( .A(n290), .Y(n21) );
  BUFX3 U42 ( .A(n288), .Y(n19) );
  BUFX3 U43 ( .A(n356), .Y(n17) );
  XNOR2X1 U44 ( .A(params[11]), .B(n209), .Y(n421) );
  AOI21X1 U45 ( .A0(n440), .A1(n441), .B0(n339), .Y(N215) );
  AOI21X1 U46 ( .A0(n438), .A1(n439), .B0(n339), .Y(N216) );
  INVX1 U47 ( .A(n49), .Y(n48) );
  INVX1 U48 ( .A(\sub_136_2/carry[10] ), .Y(N806) );
  CLKINVX3 U49 ( .A(n1), .Y(n47) );
  CLKINVX3 U50 ( .A(n1), .Y(n46) );
  INVX1 U51 ( .A(N796), .Y(n49) );
  INVX1 U52 ( .A(n335), .Y(n172) );
  BUFX3 U53 ( .A(n307), .Y(n30) );
  AND4X2 U54 ( .A(n176), .B(n333), .C(n334), .D(n335), .Y(n307) );
  CLKINVX3 U55 ( .A(n294), .Y(n37) );
  INVX1 U56 ( .A(pow[1]), .Y(n53) );
  INVX1 U57 ( .A(pow[3]), .Y(n54) );
  INVXL U58 ( .A(pow[5]), .Y(n51) );
  INVX1 U59 ( .A(n39), .Y(n38) );
  INVX1 U60 ( .A(N793), .Y(n39) );
  INVX1 U61 ( .A(n42), .Y(n41) );
  INVX1 U62 ( .A(N781), .Y(n42) );
  INVX1 U63 ( .A(n44), .Y(n43) );
  INVX1 U64 ( .A(N784), .Y(n44) );
  INVX1 U65 ( .A(n44), .Y(n40) );
  INVX1 U66 ( .A(n44), .Y(n45) );
  NAND2X1 U67 ( .A(N251), .B(N250), .Y(n335) );
  BUFX3 U68 ( .A(n308), .Y(n31) );
  NOR3X1 U69 ( .A(n25), .B(n172), .C(n333), .Y(n308) );
  INVX1 U70 ( .A(n116), .Y(n149) );
  INVX1 U71 ( .A(n114), .Y(n148) );
  NAND2X1 U72 ( .A(N255), .B(N251), .Y(n333) );
  INVX1 U73 ( .A(n87), .Y(N255) );
  INVX1 U74 ( .A(n86), .Y(n113) );
  BUFX3 U75 ( .A(n309), .Y(n28) );
  NOR2X1 U76 ( .A(n335), .B(n25), .Y(n309) );
  INVX1 U77 ( .A(n422), .Y(n173) );
  NAND2X1 U78 ( .A(N253), .B(N250), .Y(n334) );
  INVX1 U79 ( .A(n122), .Y(N253) );
  INVX1 U80 ( .A(n121), .Y(n151) );
  BUFX3 U81 ( .A(n306), .Y(n29) );
  NOR3X1 U82 ( .A(n25), .B(n172), .C(n334), .Y(n306) );
  INVX1 U83 ( .A(n81), .Y(n110) );
  INVX1 U84 ( .A(n79), .Y(n108) );
  INVX1 U85 ( .A(\sub_2_root_sub_0_root_sub_81_2/carry[8] ), .Y(N283) );
  BUFX3 U86 ( .A(n341), .Y(n26) );
  NOR2X1 U87 ( .A(n25), .B(N131), .Y(n341) );
  BUFX3 U88 ( .A(n342), .Y(n27) );
  AND2X2 U89 ( .A(N131), .B(n176), .Y(n342) );
  INVX1 U90 ( .A(n296), .Y(n174) );
  CLKINVX3 U91 ( .A(n25), .Y(n176) );
  CLKINVX3 U92 ( .A(n294), .Y(n36) );
  BUFX3 U93 ( .A(N630), .Y(n12) );
  INVX1 U94 ( .A(params[8]), .Y(n50) );
  NOR2X1 U95 ( .A(n171), .B(n2), .Y(n275) );
  INVX1 U96 ( .A(n480), .Y(n171) );
  AOI22X1 U97 ( .A0(N1021), .A1(n13), .B0(N934), .B1(N871), .Y(n480) );
  NOR2BX1 U98 ( .AN(n479), .B(n2), .Y(n277) );
  AOI22X1 U99 ( .A0(N1022), .A1(n13), .B0(N935), .B1(N871), .Y(n479) );
  NOR2BX1 U100 ( .AN(n478), .B(n2), .Y(n278) );
  AOI22X1 U101 ( .A0(N1023), .A1(n13), .B0(N936), .B1(N871), .Y(n478) );
  NOR2BX1 U102 ( .AN(n477), .B(n2), .Y(n279) );
  AOI22X1 U103 ( .A0(N1024), .A1(n13), .B0(N937), .B1(N871), .Y(n477) );
  NOR2BX1 U104 ( .AN(n476), .B(n2), .Y(n280) );
  AOI22X1 U105 ( .A0(N1025), .A1(n13), .B0(N938), .B1(N871), .Y(n476) );
  NOR2BX1 U106 ( .AN(n475), .B(n2), .Y(n281) );
  AOI22X1 U107 ( .A0(N1026), .A1(n13), .B0(N939), .B1(N871), .Y(n475) );
  NOR2BX1 U108 ( .AN(n474), .B(n2), .Y(n282) );
  AOI22X1 U109 ( .A0(N1027), .A1(n13), .B0(N940), .B1(N871), .Y(n474) );
  NOR2BX1 U110 ( .AN(n473), .B(n2), .Y(n283) );
  AOI22X1 U111 ( .A0(N1028), .A1(n13), .B0(N941), .B1(N871), .Y(n473) );
  AOI22X1 U112 ( .A0(N1029), .A1(n13), .B0(N942), .B1(N871), .Y(n472) );
  AOI22X1 U113 ( .A0(N1030), .A1(n13), .B0(N943), .B1(N871), .Y(n471) );
  INVX1 U114 ( .A(n123), .Y(n147) );
  INVX1 U115 ( .A(N365), .Y(n141) );
  INVX1 U116 ( .A(N238), .Y(n146) );
  NOR2BX2 U117 ( .AN(n423), .B(n421), .Y(n400) );
  AND2X2 U118 ( .A(n423), .B(n421), .Y(n401) );
  INVX1 U119 ( .A(N244), .Y(n143) );
  INVX1 U120 ( .A(n118), .Y(n150) );
  XOR2X1 U121 ( .A(n426), .B(n425), .Y(n422) );
  INVX1 U122 ( .A(N240), .Y(n145) );
  AND3X2 U123 ( .A(n422), .B(n417), .C(n424), .Y(n423) );
  AND4X2 U124 ( .A(n173), .B(n424), .C(n421), .D(n417), .Y(n399) );
  INVX1 U125 ( .A(n88), .Y(n106) );
  INVX1 U126 ( .A(N382), .Y(n105) );
  INVX1 U127 ( .A(N241), .Y(n144) );
  INVX1 U128 ( .A(n83), .Y(n112) );
  INVX1 U129 ( .A(N215), .Y(n109) );
  INVX1 U130 ( .A(N360), .Y(n140) );
  ADDFX2 U131 ( .A(N239), .B(n140), .CI(
        \sub_2_root_sub_0_root_sub_81_2/carry[1] ), .CO(
        \sub_2_root_sub_0_root_sub_81_2/carry[2] ), .S(N273) );
  INVX1 U132 ( .A(N360), .Y(n107) );
  ADDFX2 U133 ( .A(N245), .B(n142), .CI(
        \sub_2_root_sub_0_root_sub_81_2/carry[7] ), .CO(
        \sub_2_root_sub_0_root_sub_81_2/carry[8] ), .S(N279) );
  ADDFX2 U134 ( .A(N243), .B(n457), .CI(
        \sub_2_root_sub_0_root_sub_81_2/carry[5] ), .CO(
        \sub_2_root_sub_0_root_sub_81_2/carry[6] ), .S(N277) );
  ADDFX2 U135 ( .A(N240), .B(n469), .CI(
        \sub_2_root_sub_0_root_sub_81_2/carry[2] ), .CO(
        \sub_2_root_sub_0_root_sub_81_2/carry[3] ), .S(N274) );
  ADDFX2 U136 ( .A(N241), .B(n74), .CI(
        \sub_2_root_sub_0_root_sub_81_2/carry[3] ), .CO(
        \sub_2_root_sub_0_root_sub_81_2/carry[4] ), .S(N275) );
  ADDFX2 U137 ( .A(N242), .B(n459), .CI(
        \sub_2_root_sub_0_root_sub_81_2/carry[4] ), .CO(
        \sub_2_root_sub_0_root_sub_81_2/carry[5] ), .S(N276) );
  ADDFX2 U138 ( .A(N244), .B(n455), .CI(
        \sub_2_root_sub_0_root_sub_81_2/carry[6] ), .CO(
        \sub_2_root_sub_0_root_sub_81_2/carry[7] ), .S(N278) );
  INVX1 U139 ( .A(n73), .Y(n78) );
  INVX1 U140 ( .A(N130), .Y(n77) );
  INVX1 U141 ( .A(N216), .Y(n111) );
  NOR2X1 U142 ( .A(N366), .B(\sub_1_root_sub_0_root_add_81_6/carry[8] ), .Y(n5) );
  ADDFX2 U143 ( .A(N365), .B(n59), .CI(
        \sub_1_root_sub_0_root_add_81_6/carry[7] ), .CO(
        \sub_1_root_sub_0_root_add_81_6/carry[8] ), .S(N389) );
  INVX1 U144 ( .A(N220), .Y(n59) );
  INVX1 U145 ( .A(N362), .Y(n74) );
  ADDFX2 U146 ( .A(N364), .B(n58), .CI(
        \sub_1_root_sub_0_root_add_81_6/carry[6] ), .CO(
        \sub_1_root_sub_0_root_add_81_6/carry[7] ), .S(N388) );
  INVX1 U147 ( .A(N219), .Y(n58) );
  ADDFX2 U148 ( .A(N359), .B(n55), .CI(n105), .CO(
        \sub_1_root_sub_0_root_add_81_6/carry[2] ), .S(N383) );
  INVX1 U149 ( .A(N214), .Y(n55) );
  ADDFX2 U150 ( .A(N362), .B(n56), .CI(
        \sub_1_root_sub_0_root_add_81_6/carry[4] ), .CO(
        \sub_1_root_sub_0_root_add_81_6/carry[5] ), .S(N386) );
  INVX1 U151 ( .A(N217), .Y(n56) );
  ADDFX2 U152 ( .A(N363), .B(n57), .CI(
        \sub_1_root_sub_0_root_add_81_6/carry[5] ), .CO(
        \sub_1_root_sub_0_root_add_81_6/carry[6] ), .S(N387) );
  INVX1 U153 ( .A(N218), .Y(n57) );
  ADDFX2 U154 ( .A(N360), .B(n109), .CI(
        \sub_1_root_sub_0_root_add_81_6/carry[2] ), .CO(
        \sub_1_root_sub_0_root_add_81_6/carry[3] ), .S(N384) );
  ADDFX2 U155 ( .A(N361), .B(n111), .CI(
        \sub_1_root_sub_0_root_add_81_6/carry[3] ), .CO(
        \sub_1_root_sub_0_root_add_81_6/carry[4] ), .S(N385) );
  BUFX3 U156 ( .A(n166), .Y(n13) );
  INVX1 U157 ( .A(N366), .Y(n142) );
  INVX1 U158 ( .A(N128), .Y(n76) );
  INVX1 U159 ( .A(N126), .Y(n75) );
  AOI21X1 U160 ( .A0(n339), .A1(n176), .B0(n206), .Y(n296) );
  AOI21X1 U161 ( .A0(n209), .A1(n176), .B0(n47), .Y(n354) );
  BUFX3 U162 ( .A(n303), .Y(n25) );
  NAND2X1 U163 ( .A(n24), .B(n18), .Y(n303) );
  NOR2X2 U164 ( .A(n362), .B(n363), .Y(N1156) );
  BUFX3 U165 ( .A(n285), .Y(n34) );
  NAND2X1 U166 ( .A(n23), .B(N1156), .Y(n285) );
  BUFX3 U167 ( .A(n287), .Y(n33) );
  NAND2X1 U168 ( .A(n19), .B(N1156), .Y(n287) );
  BUFX3 U169 ( .A(n289), .Y(n32) );
  NAND2X1 U170 ( .A(n21), .B(N1156), .Y(n289) );
  BUFX3 U171 ( .A(n276), .Y(n35) );
  NAND2X1 U172 ( .A(N1156), .B(n22), .Y(n276) );
  INVX1 U173 ( .A(N1158), .Y(n178) );
  XNOR2X1 U174 ( .A(N1159), .B(n178), .Y(N1075) );
  CLKINVX3 U175 ( .A(n18), .Y(n206) );
  OAI21XL U176 ( .A0(n24), .A1(n206), .B0(n294), .Y(n519) );
  NAND2X1 U177 ( .A(n18), .B(n363), .Y(n291) );
  BUFX4 U178 ( .A(n208), .Y(n14) );
  INVX1 U179 ( .A(n292), .Y(n208) );
  NAND2X1 U180 ( .A(n294), .B(n292), .Y(n518) );
  NOR3X1 U181 ( .A(i_res[1]), .B(i_res[2]), .C(n271), .Y(n284) );
  NOR3X1 U182 ( .A(i_res[0]), .B(i_res[2]), .C(n270), .Y(n286) );
  NOR3X1 U183 ( .A(n270), .B(i_res[2]), .C(n271), .Y(n288) );
  OAI2BB2X1 U184 ( .B0(n275), .B1(n35), .A0N(block_out[0]), .A1N(n35), .Y(n485) );
  OAI2BB2X1 U185 ( .B0(n275), .B1(n34), .A0N(block_out[8]), .A1N(n34), .Y(n493) );
  OAI2BB2X1 U186 ( .B0(n275), .B1(n33), .A0N(block_out[16]), .A1N(n33), .Y(
        n501) );
  OAI2BB2X1 U187 ( .B0(n275), .B1(n32), .A0N(block_out[24]), .A1N(n32), .Y(
        n509) );
  INVX1 U188 ( .A(n394), .Y(n197) );
  AOI221X1 U189 ( .A0(n19), .A1(Im_block[16]), .B0(n21), .B1(Im_block[24]), 
        .C0(n205), .Y(n394) );
  INVX1 U190 ( .A(n395), .Y(n205) );
  AOI22X1 U191 ( .A0(Im_block[0]), .A1(n22), .B0(Im_block[8]), .B1(n23), .Y(
        n395) );
  INVX1 U192 ( .A(n392), .Y(n195) );
  AOI221X1 U193 ( .A0(n19), .A1(Im_block[17]), .B0(n21), .B1(Im_block[25]), 
        .C0(n204), .Y(n392) );
  INVX1 U194 ( .A(n393), .Y(n204) );
  AOI22X1 U195 ( .A0(Im_block[1]), .A1(n22), .B0(Im_block[9]), .B1(n23), .Y(
        n393) );
  INVX1 U196 ( .A(n388), .Y(n191) );
  AOI221X1 U197 ( .A0(n19), .A1(Im_block[19]), .B0(n21), .B1(Im_block[27]), 
        .C0(n202), .Y(n388) );
  INVX1 U198 ( .A(n389), .Y(n202) );
  AOI22X1 U199 ( .A0(Im_block[3]), .A1(n22), .B0(Im_block[11]), .B1(n23), .Y(
        n389) );
  INVX1 U200 ( .A(n390), .Y(n193) );
  AOI221X1 U201 ( .A0(n19), .A1(Im_block[18]), .B0(n21), .B1(Im_block[26]), 
        .C0(n203), .Y(n390) );
  INVX1 U202 ( .A(n391), .Y(n203) );
  AOI22X1 U203 ( .A0(Im_block[2]), .A1(n22), .B0(Im_block[10]), .B1(n23), .Y(
        n391) );
  INVX1 U204 ( .A(n386), .Y(n189) );
  AOI221X1 U205 ( .A0(n19), .A1(Im_block[20]), .B0(n21), .B1(Im_block[28]), 
        .C0(n201), .Y(n386) );
  INVX1 U206 ( .A(n387), .Y(n201) );
  AOI22X1 U207 ( .A0(Im_block[4]), .A1(n22), .B0(Im_block[12]), .B1(n23), .Y(
        n387) );
  NAND2X1 U208 ( .A(n378), .B(n379), .Y(N958) );
  AOI22X1 U209 ( .A0(W_block[0]), .A1(n22), .B0(W_block[8]), .B1(n23), .Y(n379) );
  AOI22X1 U210 ( .A0(W_block[16]), .A1(n19), .B0(W_block[24]), .B1(n21), .Y(
        n378) );
  NAND2X1 U211 ( .A(n376), .B(n377), .Y(N959) );
  AOI22X1 U212 ( .A0(W_block[1]), .A1(n22), .B0(W_block[9]), .B1(n23), .Y(n377) );
  AOI22X1 U213 ( .A0(W_block[17]), .A1(n19), .B0(W_block[25]), .B1(n21), .Y(
        n376) );
  NAND2X1 U214 ( .A(n372), .B(n373), .Y(N961) );
  AOI22X1 U215 ( .A0(W_block[3]), .A1(n22), .B0(W_block[11]), .B1(n23), .Y(
        n373) );
  AOI22X1 U216 ( .A0(W_block[19]), .A1(n19), .B0(W_block[27]), .B1(n21), .Y(
        n372) );
  NAND2X1 U217 ( .A(n374), .B(n375), .Y(N960) );
  AOI22X1 U218 ( .A0(W_block[2]), .A1(n22), .B0(W_block[10]), .B1(n23), .Y(
        n375) );
  AOI22X1 U219 ( .A0(W_block[18]), .A1(n19), .B0(W_block[26]), .B1(n21), .Y(
        n374) );
  NAND2X1 U220 ( .A(n370), .B(n371), .Y(N962) );
  AOI22X1 U221 ( .A0(W_block[4]), .A1(n22), .B0(W_block[12]), .B1(n23), .Y(
        n371) );
  AOI22X1 U222 ( .A0(W_block[20]), .A1(n19), .B0(W_block[28]), .B1(n21), .Y(
        n370) );
  NAND2X1 U223 ( .A(n368), .B(n369), .Y(N963) );
  AOI22X1 U224 ( .A0(W_block[5]), .A1(n22), .B0(W_block[13]), .B1(n23), .Y(
        n369) );
  AOI22X1 U225 ( .A0(W_block[21]), .A1(n19), .B0(W_block[29]), .B1(n21), .Y(
        n368) );
  NAND2X1 U226 ( .A(n366), .B(n367), .Y(N964) );
  AOI22X1 U227 ( .A0(W_block[6]), .A1(n22), .B0(W_block[14]), .B1(n23), .Y(
        n367) );
  AOI22X1 U228 ( .A0(W_block[22]), .A1(n19), .B0(W_block[30]), .B1(n21), .Y(
        n366) );
  NOR3X1 U229 ( .A(i_res[0]), .B(i_res[1]), .C(n268), .Y(n290) );
  INVX1 U230 ( .A(n380), .Y(n183) );
  AOI221X1 U231 ( .A0(n19), .A1(Im_block[23]), .B0(n21), .B1(Im_block[31]), 
        .C0(n198), .Y(n380) );
  INVX1 U232 ( .A(n381), .Y(n198) );
  AOI22X1 U233 ( .A0(Im_block[7]), .A1(n22), .B0(Im_block[15]), .B1(n23), .Y(
        n381) );
  INVX1 U234 ( .A(n384), .Y(n187) );
  AOI221X1 U235 ( .A0(n19), .A1(Im_block[21]), .B0(n21), .B1(Im_block[29]), 
        .C0(n200), .Y(n384) );
  INVX1 U236 ( .A(n385), .Y(n200) );
  AOI22X1 U237 ( .A0(Im_block[5]), .A1(n22), .B0(Im_block[13]), .B1(n23), .Y(
        n385) );
  INVX1 U238 ( .A(n382), .Y(n185) );
  AOI221X1 U239 ( .A0(n19), .A1(Im_block[22]), .B0(n21), .B1(Im_block[30]), 
        .C0(n199), .Y(n382) );
  INVX1 U240 ( .A(n383), .Y(n199) );
  AOI22X1 U241 ( .A0(Im_block[6]), .A1(n22), .B0(Im_block[14]), .B1(n23), .Y(
        n383) );
  NAND2X1 U242 ( .A(n364), .B(n365), .Y(N965) );
  AOI22X1 U243 ( .A0(W_block[7]), .A1(n22), .B0(W_block[15]), .B1(n23), .Y(
        n365) );
  AOI22X1 U244 ( .A0(W_block[23]), .A1(n19), .B0(W_block[31]), .B1(n21), .Y(
        n364) );
  OAI2BB2X1 U245 ( .B0(n277), .B1(n35), .A0N(block_out[1]), .A1N(n35), .Y(n486) );
  OAI2BB2X1 U246 ( .B0(n277), .B1(n34), .A0N(block_out[9]), .A1N(n34), .Y(n494) );
  OAI2BB2X1 U247 ( .B0(n277), .B1(n33), .A0N(block_out[17]), .A1N(n33), .Y(
        n502) );
  OAI2BB2X1 U248 ( .B0(n277), .B1(n32), .A0N(block_out[25]), .A1N(n32), .Y(
        n510) );
  OAI2BB2X1 U249 ( .B0(n278), .B1(n35), .A0N(block_out[2]), .A1N(n35), .Y(n487) );
  OAI2BB2X1 U250 ( .B0(n278), .B1(n34), .A0N(block_out[10]), .A1N(n34), .Y(
        n495) );
  OAI2BB2X1 U252 ( .B0(n278), .B1(n33), .A0N(block_out[18]), .A1N(n33), .Y(
        n503) );
  OAI2BB2X1 U253 ( .B0(n278), .B1(n32), .A0N(block_out[26]), .A1N(n32), .Y(
        n511) );
  OAI2BB2X1 U254 ( .B0(n279), .B1(n35), .A0N(block_out[3]), .A1N(n35), .Y(n488) );
  OAI2BB2X1 U255 ( .B0(n279), .B1(n34), .A0N(block_out[11]), .A1N(n34), .Y(
        n496) );
  OAI2BB2X1 U256 ( .B0(n279), .B1(n33), .A0N(block_out[19]), .A1N(n33), .Y(
        n504) );
  OAI2BB2X1 U257 ( .B0(n279), .B1(n32), .A0N(block_out[27]), .A1N(n32), .Y(
        n512) );
  OAI2BB2X1 U258 ( .B0(n280), .B1(n35), .A0N(block_out[4]), .A1N(n35), .Y(n489) );
  OAI2BB2X1 U259 ( .B0(n280), .B1(n34), .A0N(block_out[12]), .A1N(n34), .Y(
        n497) );
  OAI2BB2X1 U260 ( .B0(n280), .B1(n33), .A0N(block_out[20]), .A1N(n33), .Y(
        n505) );
  OAI2BB2X1 U261 ( .B0(n280), .B1(n32), .A0N(block_out[28]), .A1N(n32), .Y(
        n513) );
  OAI2BB2X1 U262 ( .B0(n281), .B1(n35), .A0N(block_out[5]), .A1N(n35), .Y(n490) );
  OAI2BB2X1 U263 ( .B0(n281), .B1(n34), .A0N(block_out[13]), .A1N(n34), .Y(
        n498) );
  OAI2BB2X1 U264 ( .B0(n281), .B1(n33), .A0N(block_out[21]), .A1N(n33), .Y(
        n506) );
  OAI2BB2X1 U265 ( .B0(n281), .B1(n32), .A0N(block_out[29]), .A1N(n32), .Y(
        n514) );
  OAI2BB2X1 U266 ( .B0(n282), .B1(n35), .A0N(block_out[6]), .A1N(n35), .Y(n491) );
  OAI2BB2X1 U267 ( .B0(n282), .B1(n34), .A0N(block_out[14]), .A1N(n34), .Y(
        n499) );
  OAI2BB2X1 U268 ( .B0(n282), .B1(n33), .A0N(block_out[22]), .A1N(n33), .Y(
        n507) );
  OAI2BB2X1 U269 ( .B0(n282), .B1(n32), .A0N(block_out[30]), .A1N(n32), .Y(
        n515) );
  OAI2BB2X1 U270 ( .B0(n283), .B1(n35), .A0N(block_out[7]), .A1N(n35), .Y(n492) );
  OAI2BB2X1 U271 ( .B0(n283), .B1(n34), .A0N(block_out[15]), .A1N(n34), .Y(
        n500) );
  OAI2BB2X1 U272 ( .B0(n283), .B1(n33), .A0N(block_out[23]), .A1N(n33), .Y(
        n508) );
  OAI2BB2X1 U273 ( .B0(n283), .B1(n32), .A0N(block_out[31]), .A1N(n32), .Y(
        n516) );
  AOI21X2 U274 ( .A0(n415), .A1(n416), .B0(n398), .Y(N238) );
  AOI22X1 U275 ( .A0(n399), .A1(Im_block[0]), .B0(n400), .B1(Im_block[8]), .Y(
        n416) );
  AOI22X1 U276 ( .A0(n401), .A1(Im_block[16]), .B0(n402), .B1(Im_block[24]), 
        .Y(n415) );
  AOI22X1 U277 ( .A0(i[1]), .A1(params[12]), .B0(n425), .B1(n426), .Y(n424) );
  XOR2X1 U278 ( .A(i[2]), .B(n424), .Y(n417) );
  INVX1 U279 ( .A(i[1]), .Y(n210) );
  XNOR2X1 U280 ( .A(params[12]), .B(n210), .Y(n425) );
  NAND2X1 U281 ( .A(n304), .B(n305), .Y(n522) );
  AOI222X1 U282 ( .A0(N332), .A1(n29), .B0(N405), .B1(n30), .C0(N357), .C1(n31), .Y(n305) );
  NAND2X1 U283 ( .A(n311), .B(n312), .Y(n523) );
  AOI22X1 U284 ( .A0(N306), .A1(n28), .B0(sum5[10]), .B1(n46), .Y(n311) );
  AOI222X1 U285 ( .A0(N331), .A1(n29), .B0(N404), .B1(n30), .C0(N356), .C1(n31), .Y(n312) );
  NAND2X1 U286 ( .A(n313), .B(n314), .Y(n524) );
  AOI22X1 U288 ( .A0(N305), .A1(n28), .B0(sum5[9]), .B1(n46), .Y(n313) );
  AOI222X1 U289 ( .A0(N330), .A1(n29), .B0(N403), .B1(n30), .C0(N355), .C1(n31), .Y(n314) );
  NAND2X1 U290 ( .A(n315), .B(n316), .Y(n525) );
  AOI22X1 U291 ( .A0(N304), .A1(n28), .B0(sum5[8]), .B1(n46), .Y(n315) );
  AOI222X1 U292 ( .A0(N329), .A1(n29), .B0(N402), .B1(n30), .C0(N354), .C1(n31), .Y(n316) );
  NAND2X1 U293 ( .A(n317), .B(n318), .Y(n526) );
  AOI222X1 U294 ( .A0(N328), .A1(n29), .B0(N401), .B1(n30), .C0(N353), .C1(n31), .Y(n318) );
  NAND2X1 U295 ( .A(n319), .B(n320), .Y(n527) );
  AOI222X1 U296 ( .A0(N327), .A1(n29), .B0(N400), .B1(n30), .C0(N352), .C1(n31), .Y(n320) );
  NAND2X1 U297 ( .A(n321), .B(n322), .Y(n528) );
  AOI222X1 U298 ( .A0(N326), .A1(n29), .B0(N399), .B1(n30), .C0(N351), .C1(n31), .Y(n322) );
  NAND2X1 U299 ( .A(n323), .B(n324), .Y(n529) );
  AOI222X1 U300 ( .A0(N325), .A1(n29), .B0(N398), .B1(n30), .C0(N350), .C1(n31), .Y(n324) );
  NAND2X1 U301 ( .A(n325), .B(n326), .Y(n530) );
  AOI222X1 U302 ( .A0(N324), .A1(n29), .B0(N397), .B1(n30), .C0(N349), .C1(n31), .Y(n326) );
  NAND2X1 U303 ( .A(n327), .B(n328), .Y(n531) );
  AOI222X1 U304 ( .A0(N323), .A1(n29), .B0(N396), .B1(n30), .C0(N348), .C1(n31), .Y(n328) );
  NAND2X1 U305 ( .A(n329), .B(n330), .Y(n532) );
  AOI222X1 U306 ( .A0(N322), .A1(n29), .B0(N395), .B1(n30), .C0(N347), .C1(n31), .Y(n330) );
  NAND2X1 U307 ( .A(n331), .B(n332), .Y(n533) );
  AOI22X1 U308 ( .A0(N296), .A1(n28), .B0(sum5[0]), .B1(n46), .Y(n331) );
  AOI222X1 U309 ( .A0(N321), .A1(n29), .B0(N394), .B1(n30), .C0(N346), .C1(n31), .Y(n332) );
  OAI211X4 U310 ( .A0(params[10]), .A1(n417), .B0(n418), .C0(n419), .Y(n398)
         );
  NAND3X1 U311 ( .A(n180), .B(n181), .C(n422), .Y(n418) );
  NAND4X1 U312 ( .A(n420), .B(n421), .C(n180), .D(n50), .Y(n419) );
  NAND2X1 U313 ( .A(n173), .B(params[9]), .Y(n420) );
  AOI21X2 U314 ( .A0(n411), .A1(n412), .B0(n398), .Y(N240) );
  AOI22X1 U315 ( .A0(n399), .A1(Im_block[2]), .B0(n400), .B1(Im_block[10]), 
        .Y(n412) );
  AOI22X1 U316 ( .A0(n401), .A1(Im_block[18]), .B0(n402), .B1(Im_block[26]), 
        .Y(n411) );
  AOI21X2 U317 ( .A0(n413), .A1(n414), .B0(n398), .Y(N239) );
  AOI22X1 U318 ( .A0(n399), .A1(Im_block[1]), .B0(n400), .B1(Im_block[9]), .Y(
        n414) );
  AOI22X1 U319 ( .A0(n401), .A1(Im_block[17]), .B0(n402), .B1(Im_block[25]), 
        .Y(n413) );
  CLKINVX3 U320 ( .A(i[0]), .Y(n209) );
  AND2X2 U321 ( .A(params[11]), .B(i[0]), .Y(n426) );
  AOI21X2 U322 ( .A0(n444), .A1(n445), .B0(n339), .Y(N382) );
  AOI22X1 U323 ( .A0(n16), .A1(Im_block[16]), .B0(Im_block[24]), .B1(n17), .Y(
        n444) );
  AOI22X1 U324 ( .A0(n429), .A1(Im_block[0]), .B0(n15), .B1(Im_block[8]), .Y(
        n445) );
  AOI21X2 U325 ( .A0(n407), .A1(n408), .B0(n398), .Y(N242) );
  AOI22X1 U326 ( .A0(n399), .A1(Im_block[4]), .B0(n400), .B1(Im_block[12]), 
        .Y(n408) );
  AOI22X1 U327 ( .A0(n401), .A1(Im_block[20]), .B0(n402), .B1(Im_block[28]), 
        .Y(n407) );
  AOI21X2 U328 ( .A0(n409), .A1(n410), .B0(n398), .Y(N241) );
  AOI22X1 U329 ( .A0(n399), .A1(Im_block[3]), .B0(n400), .B1(Im_block[11]), 
        .Y(n410) );
  AOI22X1 U330 ( .A0(n401), .A1(Im_block[19]), .B0(n402), .B1(Im_block[27]), 
        .Y(n409) );
  INVX1 U332 ( .A(params[10]), .Y(n180) );
  INVX1 U333 ( .A(params[9]), .Y(n181) );
  AOI21X2 U334 ( .A0(n403), .A1(n404), .B0(n398), .Y(N244) );
  AOI22X1 U335 ( .A0(n399), .A1(Im_block[6]), .B0(n400), .B1(Im_block[14]), 
        .Y(n404) );
  AOI22X1 U336 ( .A0(n401), .A1(Im_block[22]), .B0(n402), .B1(Im_block[30]), 
        .Y(n403) );
  AOI21X2 U337 ( .A0(n405), .A1(n406), .B0(n398), .Y(N243) );
  AOI22X1 U338 ( .A0(n399), .A1(Im_block[5]), .B0(n400), .B1(Im_block[13]), 
        .Y(n406) );
  AOI22X1 U339 ( .A0(n401), .A1(Im_block[21]), .B0(n402), .B1(Im_block[29]), 
        .Y(n405) );
  AOI22X1 U340 ( .A0(n16), .A1(Im_block[18]), .B0(Im_block[26]), .B1(n17), .Y(
        n440) );
  AOI22X1 U341 ( .A0(n429), .A1(Im_block[2]), .B0(n15), .B1(Im_block[10]), .Y(
        n441) );
  BUFX3 U342 ( .A(n430), .Y(n15) );
  CLKINVX3 U343 ( .A(n483), .Y(N359) );
  AOI221X1 U344 ( .A0(Im_block[0]), .A1(n15), .B0(Im_block[8]), .B1(n16), .C0(
        n196), .Y(n483) );
  INVX1 U345 ( .A(n484), .Y(n196) );
  AOI22X1 U346 ( .A0(Im_block[16]), .A1(n17), .B0(n454), .B1(Im_block[24]), 
        .Y(n484) );
  INVX1 U347 ( .A(i[2]), .Y(n211) );
  NOR3X1 U348 ( .A(n210), .B(i[2]), .C(n209), .Y(n356) );
  BUFX3 U349 ( .A(n431), .Y(n16) );
  CLKINVX3 U350 ( .A(n481), .Y(N360) );
  AOI221X1 U351 ( .A0(Im_block[1]), .A1(n15), .B0(Im_block[9]), .B1(n16), .C0(
        n194), .Y(n481) );
  INVX1 U352 ( .A(n482), .Y(n194) );
  AOI22X1 U353 ( .A0(Im_block[17]), .A1(n17), .B0(n454), .B1(Im_block[25]), 
        .Y(n482) );
  CLKINVX3 U354 ( .A(n469), .Y(N361) );
  AOI221X1 U355 ( .A0(Im_block[2]), .A1(n15), .B0(Im_block[10]), .B1(n16), 
        .C0(n192), .Y(n469) );
  INVX1 U356 ( .A(n470), .Y(n192) );
  AOI22X1 U357 ( .A0(Im_block[18]), .A1(n17), .B0(n454), .B1(Im_block[26]), 
        .Y(n470) );
  AOI21X2 U358 ( .A0(n396), .A1(n397), .B0(n398), .Y(N245) );
  AOI22X1 U359 ( .A0(n399), .A1(Im_block[7]), .B0(n400), .B1(Im_block[15]), 
        .Y(n397) );
  AOI22X1 U360 ( .A0(n401), .A1(Im_block[23]), .B0(n402), .B1(Im_block[31]), 
        .Y(n396) );
  CLKINVX3 U361 ( .A(n459), .Y(N363) );
  AOI221X1 U362 ( .A0(Im_block[4]), .A1(n15), .B0(Im_block[12]), .B1(n16), 
        .C0(n188), .Y(n459) );
  INVX1 U363 ( .A(n460), .Y(n188) );
  AOI22X1 U364 ( .A0(Im_block[20]), .A1(n17), .B0(n454), .B1(Im_block[28]), 
        .Y(n460) );
  AND3X2 U365 ( .A(n446), .B(n447), .C(n448), .Y(n339) );
  XNOR2X1 U366 ( .A(endOfRow[0]), .B(i[0]), .Y(n447) );
  XNOR2X1 U367 ( .A(endOfRow[1]), .B(i[1]), .Y(n446) );
  XNOR2X1 U368 ( .A(endOfRow[2]), .B(i[2]), .Y(n448) );
  AOI22X1 U369 ( .A0(n16), .A1(Im_block[19]), .B0(Im_block[27]), .B1(n17), .Y(
        n438) );
  AOI22X1 U370 ( .A0(n429), .A1(Im_block[3]), .B0(n15), .B1(Im_block[11]), .Y(
        n439) );
  AOI21X2 U371 ( .A0(n442), .A1(n443), .B0(n339), .Y(N214) );
  AOI22X1 U372 ( .A0(n16), .A1(Im_block[17]), .B0(Im_block[25]), .B1(n17), .Y(
        n442) );
  AOI22X1 U373 ( .A0(n429), .A1(Im_block[1]), .B0(n15), .B1(Im_block[9]), .Y(
        n443) );
  AOI21X2 U374 ( .A0(n436), .A1(n437), .B0(n339), .Y(N217) );
  AOI22X1 U375 ( .A0(n16), .A1(Im_block[20]), .B0(Im_block[28]), .B1(n17), .Y(
        n436) );
  AOI22X1 U376 ( .A0(n429), .A1(Im_block[4]), .B0(n15), .B1(Im_block[12]), .Y(
        n437) );
  OAI2BB1X1 U377 ( .A0N(sum4[0]), .A1N(n47), .B0(n353), .Y(n546) );
  AOI22X1 U378 ( .A0(N179), .A1(n26), .B0(N150), .B1(n27), .Y(n353) );
  OAI2BB1X1 U379 ( .A0N(sum4[1]), .A1N(n47), .B0(n352), .Y(n545) );
  AOI22X1 U380 ( .A0(N180), .A1(n26), .B0(N151), .B1(n27), .Y(n352) );
  OAI2BB1X1 U381 ( .A0N(sum4[2]), .A1N(n47), .B0(n351), .Y(n544) );
  AOI22X1 U382 ( .A0(N181), .A1(n26), .B0(N152), .B1(n27), .Y(n351) );
  OAI2BB1X1 U383 ( .A0N(sum4[3]), .A1N(n47), .B0(n350), .Y(n543) );
  AOI22X1 U384 ( .A0(N182), .A1(n26), .B0(N153), .B1(n27), .Y(n350) );
  OAI2BB1X1 U385 ( .A0N(sum4[4]), .A1N(n47), .B0(n349), .Y(n542) );
  AOI22X1 U386 ( .A0(N183), .A1(n26), .B0(N154), .B1(n27), .Y(n349) );
  OAI2BB1X1 U387 ( .A0N(sum4[5]), .A1N(n47), .B0(n348), .Y(n541) );
  AOI22X1 U388 ( .A0(N184), .A1(n26), .B0(N155), .B1(n27), .Y(n348) );
  OAI2BB1X1 U389 ( .A0N(sum4[6]), .A1N(n47), .B0(n347), .Y(n540) );
  AOI22X1 U390 ( .A0(N185), .A1(n26), .B0(N156), .B1(n27), .Y(n347) );
  OAI2BB1X1 U391 ( .A0N(sum4[7]), .A1N(n47), .B0(n346), .Y(n539) );
  AOI22X1 U392 ( .A0(N186), .A1(n26), .B0(N157), .B1(n27), .Y(n346) );
  OAI2BB1X1 U393 ( .A0N(sum4[8]), .A1N(n47), .B0(n345), .Y(n538) );
  AOI22X1 U394 ( .A0(N187), .A1(n26), .B0(N158), .B1(n27), .Y(n345) );
  OAI2BB1X1 U395 ( .A0N(sum4[9]), .A1N(n47), .B0(n344), .Y(n537) );
  AOI22X1 U396 ( .A0(N188), .A1(n26), .B0(N159), .B1(n27), .Y(n344) );
  OAI2BB1X1 U397 ( .A0N(sum4[10]), .A1N(n47), .B0(n343), .Y(n536) );
  AOI22X1 U398 ( .A0(N189), .A1(n26), .B0(N160), .B1(n27), .Y(n343) );
  OAI2BB1X1 U399 ( .A0N(sum4[11]), .A1N(n47), .B0(n340), .Y(n535) );
  AOI22X1 U400 ( .A0(N190), .A1(n26), .B0(N161), .B1(n27), .Y(n340) );
  CLKINVX3 U401 ( .A(n461), .Y(N362) );
  AOI221X1 U402 ( .A0(Im_block[3]), .A1(n15), .B0(Im_block[11]), .B1(n16), 
        .C0(n190), .Y(n461) );
  INVX1 U403 ( .A(n462), .Y(n190) );
  AOI22X1 U404 ( .A0(Im_block[19]), .A1(n17), .B0(n454), .B1(Im_block[27]), 
        .Y(n462) );
  AOI21X2 U405 ( .A0(n434), .A1(n435), .B0(n339), .Y(N218) );
  AOI22X1 U406 ( .A0(n16), .A1(Im_block[21]), .B0(Im_block[29]), .B1(n17), .Y(
        n434) );
  AOI22X1 U407 ( .A0(n429), .A1(Im_block[5]), .B0(n15), .B1(Im_block[13]), .Y(
        n435) );
  AOI21X2 U408 ( .A0(n432), .A1(n433), .B0(n339), .Y(N219) );
  AOI22X1 U409 ( .A0(n16), .A1(Im_block[22]), .B0(Im_block[30]), .B1(n17), .Y(
        n432) );
  AOI22X1 U410 ( .A0(n429), .A1(Im_block[6]), .B0(n15), .B1(Im_block[14]), .Y(
        n433) );
  CLKINVX3 U411 ( .A(n455), .Y(N365) );
  AOI221X1 U412 ( .A0(Im_block[6]), .A1(n15), .B0(Im_block[14]), .B1(n16), 
        .C0(n184), .Y(n455) );
  INVX1 U413 ( .A(n456), .Y(n184) );
  AOI22X1 U414 ( .A0(Im_block[22]), .A1(n17), .B0(n454), .B1(Im_block[30]), 
        .Y(n456) );
  CLKINVX3 U415 ( .A(n457), .Y(N364) );
  AOI221X1 U416 ( .A0(Im_block[5]), .A1(n15), .B0(Im_block[13]), .B1(n16), 
        .C0(n186), .Y(n457) );
  INVX1 U417 ( .A(n458), .Y(n186) );
  AOI22X1 U418 ( .A0(Im_block[21]), .A1(n17), .B0(n454), .B1(Im_block[29]), 
        .Y(n458) );
  CLKINVX3 U419 ( .A(n166), .Y(N871) );
  INVX1 U420 ( .A(params[20]), .Y(n170) );
  AOI21X2 U421 ( .A0(n427), .A1(n428), .B0(n339), .Y(N220) );
  AOI22X1 U422 ( .A0(n16), .A1(Im_block[23]), .B0(Im_block[31]), .B1(n17), .Y(
        n427) );
  AOI22X1 U423 ( .A0(n429), .A1(Im_block[7]), .B0(n15), .B1(Im_block[15]), .Y(
        n428) );
  CLKINVX3 U424 ( .A(n452), .Y(N366) );
  AOI221X1 U425 ( .A0(Im_block[7]), .A1(n15), .B0(Im_block[15]), .B1(n16), 
        .C0(n182), .Y(n452) );
  INVX1 U426 ( .A(n453), .Y(n182) );
  AOI22X1 U427 ( .A0(Im_block[23]), .A1(n17), .B0(n454), .B1(Im_block[31]), 
        .Y(n453) );
  AOI21X1 U428 ( .A0(params[14]), .A1(n7), .B0(params[13]), .Y(n156) );
  INVX1 U429 ( .A(params[14]), .Y(n167) );
  INVX1 U430 ( .A(params[16]), .Y(n168) );
  INVX1 U431 ( .A(params[19]), .Y(n169) );
  OAI21XL U432 ( .A0(n301), .A1(n212), .B0(n302), .Y(n521) );
  AOI2BB1X1 U433 ( .A0N(n25), .A1N(params[11]), .B0(n296), .Y(n301) );
  OAI211X1 U434 ( .A0(n206), .A1(n212), .B0(n174), .C0(params[11]), .Y(n302)
         );
  INVX1 U435 ( .A(endOfRow[0]), .Y(n212) );
  INVX1 U436 ( .A(n355), .Y(n175) );
  AOI22X1 U437 ( .A0(n176), .A1(n17), .B0(n357), .B1(i[2]), .Y(n355) );
  OAI21XL U438 ( .A0(n25), .A1(i[1]), .B0(n354), .Y(n357) );
  NAND2X1 U439 ( .A(params[10]), .B(n211), .Y(n359) );
  OAI21XL U440 ( .A0(n336), .A1(n214), .B0(n337), .Y(n534) );
  AOI21X1 U441 ( .A0(n338), .A1(n176), .B0(n296), .Y(n336) );
  NAND4BXL U442 ( .AN(n338), .B(n176), .C(n174), .D(n214), .Y(n337) );
  AOI22X1 U443 ( .A0(endOfRow[1]), .A1(params[12]), .B0(n300), .B1(n299), .Y(
        n338) );
  BUFX3 U444 ( .A(n295), .Y(n24) );
  AOI31X1 U445 ( .A0(n358), .A1(n50), .A2(n359), .B0(n177), .Y(n295) );
  AOI21X1 U446 ( .A0(n210), .A1(params[9]), .B0(n209), .Y(n358) );
  OAI32X1 U447 ( .A0(n25), .A1(i[1]), .A2(n209), .B0(n354), .B1(n210), .Y(n547) );
  INVX1 U448 ( .A(n360), .Y(n177) );
  AOI32X1 U449 ( .A0(n359), .A1(n181), .A2(i[1]), .B0(i[2]), .B1(n180), .Y(
        n360) );
  OAI221XL U450 ( .A0(i[0]), .A1(n25), .B0(n209), .B1(n1), .C0(n18), .Y(n548)
         );
  NOR2X1 U451 ( .A(n180), .B(i_res[2]), .Y(n450) );
  OAI22X1 U452 ( .A0(n213), .A1(n174), .B0(n296), .B1(n297), .Y(n520) );
  AOI22X1 U453 ( .A0(n176), .A1(n298), .B0(params[12]), .B1(n206), .Y(n297) );
  XOR2X1 U454 ( .A(n299), .B(n300), .Y(n298) );
  OAI31X1 U455 ( .A0(n449), .A1(params[8]), .A2(n450), .B0(n451), .Y(n362) );
  OAI21XL U456 ( .A0(i_res[1]), .A1(n181), .B0(i_res[0]), .Y(n449) );
  AOI32X1 U457 ( .A0(n179), .A1(n181), .A2(i_res[1]), .B0(i_res[2]), .B1(n180), 
        .Y(n451) );
  INVX1 U458 ( .A(n450), .Y(n179) );
  AND2X2 U459 ( .A(i_res[0]), .B(N1156), .Y(N1158) );
  AND2X2 U460 ( .A(i_res[1]), .B(N1156), .Y(N1159) );
  XOR2X1 U461 ( .A(n10), .B(n11), .Y(N1076) );
  NAND2X1 U462 ( .A(N1156), .B(i_res[2]), .Y(n10) );
  NAND2X1 U463 ( .A(N1159), .B(N1158), .Y(n11) );
  NAND3X1 U464 ( .A(Ready), .B(n18), .C(eq12_done), .Y(n363) );
  BUFX4 U465 ( .A(n293), .Y(n18) );
  NOR2X1 U466 ( .A(block_done), .B(rst), .Y(n293) );
  NOR2X1 U467 ( .A(ena_in), .B(n361), .Y(n549) );
  AOI21X1 U468 ( .A0(n207), .A1(n362), .B0(n206), .Y(n361) );
  INVX1 U469 ( .A(n363), .Y(n207) );
  NAND2X1 U470 ( .A(sums_done), .B(n18), .Y(n294) );
  NAND2X1 U471 ( .A(eq345_done), .B(n18), .Y(n292) );
  XNOR2X1 U472 ( .A(n213), .B(params[12]), .Y(n300) );
  AND2X2 U473 ( .A(params[11]), .B(endOfRow[0]), .Y(n299) );
  INVX1 U474 ( .A(endOfRow[1]), .Y(n213) );
  OAI2BB1X1 U475 ( .A0N(n18), .A1N(eq12_done), .B0(n292), .Y(n517) );
  INVX1 U476 ( .A(endOfRow[2]), .Y(n214) );
  XNOR2X1 U477 ( .A(\sub_1_root_sub_0_root_add_81_6/carry[8] ), .B(N366), .Y(
        N390) );
  OR2X1 U478 ( .A(n483), .B(N238), .Y(
        \sub_2_root_sub_0_root_sub_81_2/carry[1] ) );
  XNOR2X1 U479 ( .A(N238), .B(n483), .Y(N272) );
  INVX1 U480 ( .A(\sub_136_2/carry[10] ), .Y(N805) );
  INVX1 U481 ( .A(\sub_136_2/carry[10] ), .Y(N804) );
  OR2X1 U482 ( .A(n52), .B(\sub_136_2/carry[7] ), .Y(\sub_136_2/carry[10] ) );
  XNOR2X1 U483 ( .A(\sub_136_2/carry[7] ), .B(n52), .Y(N803) );
  OR2X1 U484 ( .A(n49), .B(\sub_136_2/carry[6] ), .Y(\sub_136_2/carry[7] ) );
  XNOR2X1 U485 ( .A(\sub_136_2/carry[6] ), .B(n49), .Y(N802) );
  OR2X1 U486 ( .A(n51), .B(\sub_136_2/carry[5] ), .Y(\sub_136_2/carry[6] ) );
  XNOR2X1 U487 ( .A(\sub_136_2/carry[5] ), .B(n51), .Y(N801) );
  OR2X1 U488 ( .A(n54), .B(\sub_136_2/carry[3] ), .Y(\sub_136_2/carry[5] ) );
  XNOR2X1 U489 ( .A(\sub_136_2/carry[3] ), .B(n54), .Y(N799) );
  AND2X1 U490 ( .A(\sub_136_2/carry[2] ), .B(n52), .Y(\sub_136_2/carry[3] ) );
  XOR2X1 U491 ( .A(n52), .B(\sub_136_2/carry[2] ), .Y(N798) );
  AND2X1 U492 ( .A(n49), .B(n53), .Y(\sub_136_2/carry[2] ) );
  XOR2X1 U493 ( .A(n53), .B(n49), .Y(N797) );
  XOR2X1 U494 ( .A(\mult_134/n1 ), .B(params[27]), .Y(N590) );
  NAND2BX1 U495 ( .AN(N363), .B(N127), .Y(n60) );
  OAI222XL U496 ( .A0(n76), .A1(n60), .B0(N364), .B1(n60), .C0(N364), .C1(n76), 
        .Y(n61) );
  OAI222XL U497 ( .A0(N129), .A1(n61), .B0(n141), .B1(n61), .C0(N129), .C1(
        n141), .Y(n72) );
  NOR2BX1 U498 ( .AN(N363), .B(N127), .Y(n62) );
  OAI22X1 U499 ( .A0(n62), .A1(n76), .B0(N364), .B1(n62), .Y(n70) );
  NAND2BX1 U500 ( .AN(N125), .B(N361), .Y(n63) );
  AOI22X1 U501 ( .A0(n63), .A1(n74), .B0(n63), .B1(N126), .Y(n68) );
  AOI2BB1X1 U502 ( .A0N(n481), .A1N(N124), .B0(N359), .Y(n64) );
  AOI22X1 U503 ( .A0(N124), .A1(n107), .B0(n64), .B1(N123), .Y(n67) );
  NOR2BX1 U504 ( .AN(N125), .B(N361), .Y(n65) );
  AOI22X1 U505 ( .A0(n65), .A1(n74), .B0(N126), .B1(n65), .Y(n66) );
  OAI221XL U506 ( .A0(N362), .A1(n75), .B0(n68), .B1(n67), .C0(n66), .Y(n69)
         );
  OAI211X1 U507 ( .A0(N129), .A1(n455), .B0(n70), .C0(n69), .Y(n71) );
  AOI22X1 U508 ( .A0(n77), .A1(N366), .B0(n72), .B1(n71), .Y(n73) );
  OAI21XL U509 ( .A0(N366), .A1(n77), .B0(n78), .Y(N131) );
  NAND2X1 U510 ( .A(N220), .B(n452), .Y(n102) );
  NAND2BX1 U511 ( .AN(N217), .B(N363), .Y(n84) );
  NAND2BX1 U512 ( .AN(N363), .B(N217), .Y(n96) );
  NAND2X1 U513 ( .A(n84), .B(n96), .Y(n98) );
  NAND2X1 U514 ( .A(N359), .B(n105), .Y(n80) );
  NOR2X1 U515 ( .A(n109), .B(N361), .Y(n93) );
  NAND2X1 U516 ( .A(N361), .B(n109), .Y(n82) );
  NAND2BX1 U517 ( .AN(n93), .B(n82), .Y(n90) );
  OAI21XL U518 ( .A0(n80), .A1(n107), .B0(N214), .Y(n79) );
  AOI211X1 U519 ( .A0(n80), .A1(n107), .B0(n90), .C0(n108), .Y(n81) );
  NAND2X1 U520 ( .A(N362), .B(n111), .Y(n91) );
  NOR2X1 U521 ( .A(n111), .B(N362), .Y(n94) );
  AOI31X1 U522 ( .A0(n110), .A1(n82), .A2(n91), .B0(n94), .Y(n83) );
  NAND2BX1 U523 ( .AN(N218), .B(N364), .Y(n100) );
  OAI211X1 U524 ( .A0(n98), .A1(n112), .B0(n100), .C0(n84), .Y(n85) );
  NAND2BX1 U525 ( .AN(N364), .B(N218), .Y(n95) );
  XNOR2X1 U526 ( .A(N365), .B(N219), .Y(n99) );
  AOI32X1 U527 ( .A0(n85), .A1(n95), .A2(n99), .B0(N365), .B1(n58), .Y(n86) );
  NOR2X1 U528 ( .A(n142), .B(N220), .Y(n104) );
  AOI21X1 U529 ( .A0(n102), .A1(n113), .B0(n104), .Y(n87) );
  NOR2X1 U530 ( .A(n105), .B(N359), .Y(n88) );
  AOI21X1 U531 ( .A0(n88), .A1(n107), .B0(N214), .Y(n89) );
  AOI211X1 U532 ( .A0(N360), .A1(n106), .B0(n90), .C0(n89), .Y(n92) );
  OAI31X1 U533 ( .A0(n94), .A1(n93), .A2(n92), .B0(n91), .Y(n97) );
  OAI211X1 U534 ( .A0(n98), .A1(n97), .B0(n96), .C0(n95), .Y(n101) );
  AOI32X1 U535 ( .A0(n101), .A1(n100), .A2(n99), .B0(N219), .B1(n141), .Y(n103) );
  OAI21XL U536 ( .A0(n104), .A1(n103), .B0(n102), .Y(N250) );
  NAND2X1 U537 ( .A(N245), .B(n142), .Y(n137) );
  NAND2BX1 U538 ( .AN(N242), .B(N363), .Y(n119) );
  NAND2BX1 U539 ( .AN(N363), .B(N242), .Y(n131) );
  NAND2X1 U540 ( .A(n119), .B(n131), .Y(n133) );
  NAND2X1 U541 ( .A(N359), .B(n146), .Y(n115) );
  NOR2X1 U542 ( .A(n145), .B(N361), .Y(n128) );
  NAND2X1 U543 ( .A(N361), .B(n145), .Y(n117) );
  NAND2BX1 U544 ( .AN(n128), .B(n117), .Y(n125) );
  OAI21XL U545 ( .A0(n115), .A1(n140), .B0(N239), .Y(n114) );
  AOI211X1 U546 ( .A0(n115), .A1(n140), .B0(n125), .C0(n148), .Y(n116) );
  NAND2X1 U547 ( .A(N362), .B(n144), .Y(n126) );
  NOR2X1 U548 ( .A(n144), .B(N362), .Y(n129) );
  AOI31X1 U549 ( .A0(n149), .A1(n117), .A2(n126), .B0(n129), .Y(n118) );
  NAND2BX1 U550 ( .AN(N243), .B(N364), .Y(n135) );
  OAI211X1 U551 ( .A0(n133), .A1(n150), .B0(n135), .C0(n119), .Y(n120) );
  NAND2BX1 U552 ( .AN(N364), .B(N243), .Y(n130) );
  XNOR2X1 U553 ( .A(N365), .B(N244), .Y(n134) );
  AOI32X1 U554 ( .A0(n120), .A1(n130), .A2(n134), .B0(N365), .B1(n143), .Y(
        n121) );
  NOR2X1 U555 ( .A(n142), .B(N245), .Y(n139) );
  AOI21X1 U556 ( .A0(n137), .A1(n151), .B0(n139), .Y(n122) );
  NOR2X1 U557 ( .A(n146), .B(N359), .Y(n123) );
  AOI21X1 U558 ( .A0(n123), .A1(n140), .B0(N239), .Y(n124) );
  AOI211X1 U559 ( .A0(N360), .A1(n147), .B0(n125), .C0(n124), .Y(n127) );
  OAI31X1 U560 ( .A0(n129), .A1(n128), .A2(n127), .B0(n126), .Y(n132) );
  OAI211X1 U561 ( .A0(n133), .A1(n132), .B0(n131), .C0(n130), .Y(n136) );
  AOI32X1 U562 ( .A0(n136), .A1(n135), .A2(n134), .B0(N244), .B1(n141), .Y(
        n138) );
  OAI21XL U563 ( .A0(n139), .A1(n138), .B0(n137), .Y(N251) );
  NAND2BX1 U564 ( .AN(params[17]), .B(G[4]), .Y(n152) );
  OAI222XL U565 ( .A0(n3), .A1(n152), .B0(params[18]), .B1(n152), .C0(
        params[18]), .C1(n3), .Y(n153) );
  OAI222XL U566 ( .A0(G[6]), .A1(n153), .B0(n169), .B1(n153), .C0(G[6]), .C1(
        n169), .Y(n164) );
  NOR2BX1 U567 ( .AN(params[17]), .B(G[4]), .Y(n154) );
  OAI22X1 U568 ( .A0(n154), .A1(n3), .B0(params[18]), .B1(n154), .Y(n162) );
  NAND2BX1 U569 ( .AN(G[2]), .B(params[15]), .Y(n155) );
  AOI22X1 U570 ( .A0(n155), .A1(n168), .B0(n155), .B1(G[3]), .Y(n160) );
  AOI22X1 U571 ( .A0(G[1]), .A1(n167), .B0(n156), .B1(G[0]), .Y(n159) );
  NOR2BX1 U572 ( .AN(G[2]), .B(params[15]), .Y(n157) );
  AOI22X1 U573 ( .A0(n157), .A1(n168), .B0(G[3]), .B1(n157), .Y(n158) );
  OAI221XL U574 ( .A0(params[16]), .A1(n4), .B0(n160), .B1(n159), .C0(n158), 
        .Y(n161) );
  OAI211X1 U575 ( .A0(G[6]), .A1(n169), .B0(n162), .C0(n161), .Y(n163) );
  AOI2BB2X1 U576 ( .B0(n164), .B1(n163), .A0N(n170), .A1N(G[7]), .Y(n165) );
  AOI211X1 U577 ( .A0(G[7]), .A1(n170), .B0(n165), .C0(G[8]), .Y(n166) );
endmodule


module Control_And_Registers_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [19:0] A;
  input [19:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175;

  INVX1 U59 ( .A(B[3]), .Y(n121) );
  INVX1 U60 ( .A(B[6]), .Y(n120) );
  INVX1 U61 ( .A(B[9]), .Y(n119) );
  INVX1 U62 ( .A(B[13]), .Y(n122) );
  INVX1 U63 ( .A(B[15]), .Y(n123) );
  INVX1 U64 ( .A(B[18]), .Y(n125) );
  INVX1 U65 ( .A(n150), .Y(n118) );
  INVX1 U66 ( .A(B[1]), .Y(n117) );
  INVX1 U67 ( .A(n139), .Y(n124) );
  INVX1 U68 ( .A(A[12]), .Y(n129) );
  INVX1 U69 ( .A(A[8]), .Y(n131) );
  INVX1 U70 ( .A(A[17]), .Y(n127) );
  INVX1 U71 ( .A(A[5]), .Y(n132) );
  INVX1 U72 ( .A(A[14]), .Y(n128) );
  INVX1 U73 ( .A(A[10]), .Y(n130) );
  INVX1 U74 ( .A(A[19]), .Y(n126) );
  INVX1 U75 ( .A(A[3]), .Y(n133) );
  OAI221XL U76 ( .A0(B[19]), .A1(n134), .B0(B[19]), .B1(n126), .C0(n135), .Y(
        GE_LT_GT_LE) );
  AOI2BB1X1 U77 ( .A0N(n126), .A1N(n134), .B0(n136), .Y(n135) );
  AOI21X1 U78 ( .A0(n137), .A1(n138), .B0(n124), .Y(n136) );
  OAI22X1 U79 ( .A0(n140), .A1(B[19]), .B0(n140), .B1(n126), .Y(n139) );
  OAI21XL U80 ( .A0(A[18]), .A1(n125), .B0(n141), .Y(n140) );
  OAI22X1 U81 ( .A0(n142), .A1(n127), .B0(B[17]), .B1(n142), .Y(n141) );
  NOR2BX1 U82 ( .AN(B[16]), .B(A[16]), .Y(n142) );
  OAI211X1 U83 ( .A0(A[15]), .A1(n123), .B0(n143), .C0(n144), .Y(n138) );
  OAI221XL U84 ( .A0(B[10]), .A1(n145), .B0(B[10]), .B1(n130), .C0(n146), .Y(
        n144) );
  AOI2BB1X1 U85 ( .A0N(n130), .A1N(n145), .B0(n147), .Y(n146) );
  AOI21X1 U86 ( .A0(n148), .A1(n149), .B0(n118), .Y(n147) );
  OAI22X1 U87 ( .A0(n151), .A1(B[10]), .B0(n151), .B1(n130), .Y(n150) );
  OAI21XL U88 ( .A0(A[9]), .A1(n119), .B0(n152), .Y(n151) );
  OAI22X1 U89 ( .A0(n153), .A1(n131), .B0(B[8]), .B1(n153), .Y(n152) );
  NOR2BX1 U90 ( .AN(B[7]), .B(A[7]), .Y(n153) );
  OAI211X1 U91 ( .A0(A[6]), .A1(n120), .B0(n154), .C0(n155), .Y(n149) );
  OAI221XL U92 ( .A0(B[3]), .A1(n133), .B0(n156), .B1(n157), .C0(n158), .Y(
        n155) );
  AOI22X1 U93 ( .A0(n159), .A1(n121), .B0(A[3]), .B1(n159), .Y(n158) );
  NOR2BX1 U94 ( .AN(A[2]), .B(B[2]), .Y(n159) );
  AOI22X1 U95 ( .A0(A[1]), .A1(n117), .B0(n160), .B1(A[0]), .Y(n157) );
  AOI2BB1X1 U96 ( .A0N(n117), .A1N(A[1]), .B0(B[0]), .Y(n160) );
  AOI22X1 U97 ( .A0(n161), .A1(n121), .B0(n161), .B1(A[3]), .Y(n156) );
  NAND2BX1 U98 ( .AN(A[2]), .B(B[2]), .Y(n161) );
  OAI22X1 U99 ( .A0(n162), .A1(n132), .B0(B[5]), .B1(n162), .Y(n154) );
  NOR2BX1 U100 ( .AN(B[4]), .B(A[4]), .Y(n162) );
  OAI222XL U101 ( .A0(A[6]), .A1(n163), .B0(n120), .B1(n163), .C0(A[6]), .C1(
        n120), .Y(n148) );
  OAI222XL U102 ( .A0(n132), .A1(n164), .B0(B[5]), .B1(n164), .C0(B[5]), .C1(
        n132), .Y(n163) );
  NAND2BX1 U103 ( .AN(B[4]), .B(A[4]), .Y(n164) );
  OAI222XL U104 ( .A0(A[9]), .A1(n165), .B0(n165), .B1(n119), .C0(A[9]), .C1(
        n119), .Y(n145) );
  OAI222XL U105 ( .A0(n166), .A1(n131), .B0(B[8]), .B1(n166), .C0(B[8]), .C1(
        n131), .Y(n165) );
  NAND2BX1 U106 ( .AN(B[7]), .B(A[7]), .Y(n166) );
  OAI22X1 U107 ( .A0(n167), .A1(n128), .B0(B[14]), .B1(n167), .Y(n143) );
  OAI21XL U108 ( .A0(A[13]), .A1(n122), .B0(n168), .Y(n167) );
  OAI22X1 U109 ( .A0(n169), .A1(n129), .B0(B[12]), .B1(n169), .Y(n168) );
  NOR2BX1 U110 ( .AN(B[11]), .B(A[11]), .Y(n169) );
  OAI222XL U111 ( .A0(A[15]), .A1(n170), .B0(n123), .B1(n170), .C0(A[15]), 
        .C1(n123), .Y(n137) );
  OAI222XL U112 ( .A0(B[14]), .A1(n128), .B0(B[14]), .B1(n171), .C0(n128), 
        .C1(n171), .Y(n170) );
  OAI222XL U113 ( .A0(A[13]), .A1(n172), .B0(n122), .B1(n172), .C0(A[13]), 
        .C1(n122), .Y(n171) );
  OAI222XL U114 ( .A0(n129), .A1(n173), .B0(B[12]), .B1(n173), .C0(B[12]), 
        .C1(n129), .Y(n172) );
  NAND2BX1 U115 ( .AN(B[11]), .B(A[11]), .Y(n173) );
  OAI222XL U116 ( .A0(A[18]), .A1(n174), .B0(n174), .B1(n125), .C0(A[18]), 
        .C1(n125), .Y(n134) );
  OAI222XL U117 ( .A0(n175), .A1(n127), .B0(B[17]), .B1(n175), .C0(B[17]), 
        .C1(n127), .Y(n174) );
  NAND2BX1 U118 ( .AN(B[16]), .B(A[16]), .Y(n175) );
endmodule


module Control_And_Registers_DW01_add_15 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR3X2 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .Y(SUM[9]) );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module Control_And_Registers_DW01_inc_0 ( A, SUM );
  input [19:0] A;
  output [19:0] SUM;

  wire   [19:2] carry;

  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  CMPR22X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(SUM[19]), .S(SUM[18]) );
  CMPR22X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  CMPR22X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  CMPR22X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  CMPR22X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  CMPR22X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  CMPR22X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  CMPR22X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVXL U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module Control_And_Registers_DW01_inc_1 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[12]), .B(A[12]), .Y(SUM[12]) );
endmodule


module Control_And_Registers_DW_mult_uns_2 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n130,
         n131, n132, n134, n135, n136, n137, n139, n140, n141, n142, n143,
         n145, n146, n147, n148, n149, n150, n152, n153, n154, n155, n156,
         n157, n158, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329;

  ADDFX2 U3 ( .A(n30), .B(n38), .CI(n3), .CO(n2), .S(product[18]) );
  ADDFX2 U4 ( .A(n39), .B(n47), .CI(n4), .CO(n3), .S(product[17]) );
  ADDFX2 U5 ( .A(n48), .B(n58), .CI(n5), .CO(n4), .S(product[16]) );
  ADDFX2 U6 ( .A(n59), .B(n68), .CI(n6), .CO(n5), .S(product[15]) );
  ADDFX2 U7 ( .A(n69), .B(n78), .CI(n7), .CO(n6), .S(product[14]) );
  ADDFX2 U8 ( .A(n79), .B(n86), .CI(n8), .CO(n7), .S(product[13]) );
  ADDFX2 U9 ( .A(n87), .B(n94), .CI(n9), .CO(n8), .S(product[12]) );
  ADDFX2 U10 ( .A(n95), .B(n101), .CI(n10), .CO(n9), .S(product[11]) );
  ADDFX2 U11 ( .A(n102), .B(n108), .CI(n11), .CO(n10), .S(product[10]) );
  ADDFX2 U12 ( .A(n109), .B(n113), .CI(n12), .CO(n11), .S(product[9]) );
  ADDFX2 U13 ( .A(n114), .B(n117), .CI(n13), .CO(n12), .S(product[8]) );
  ADDFX2 U14 ( .A(n118), .B(n121), .CI(n14), .CO(n13), .S(product[7]) );
  ADDFX2 U15 ( .A(n122), .B(n124), .CI(n15), .CO(n14), .S(product[6]) );
  ADDFX2 U16 ( .A(n126), .B(n127), .CI(n16), .CO(n15), .S(product[5]) );
  ADDFX2 U17 ( .A(n128), .B(n209), .CI(n17), .CO(n16), .S(product[4]) );
  ADDHXL U18 ( .A(n211), .B(n18), .CO(n17), .S(product[3]) );
  ADDHXL U19 ( .A(a[1]), .B(n212), .CO(n18), .S(product[2]) );
  CMPR42X1 U29 ( .A(n40), .B(n44), .C(n33), .D(n41), .ICI(n37), .S(n30), .ICO(
        n28), .CO(n29) );
  CMPR42X1 U30 ( .A(n152), .B(n130), .C(n43), .D(n145), .ICI(n36), .S(n33), 
        .ICO(n31), .CO(n32) );
  CMPR42X1 U31 ( .A(n134), .B(a[9]), .C(n160), .D(n168), .ICI(n139), .S(n36), 
        .ICO(n34), .CO(n35) );
  CMPR42X1 U32 ( .A(n49), .B(n45), .C(n42), .D(n50), .ICI(n46), .S(n39), .ICO(
        n37), .CO(n38) );
  CMPR42X1 U33 ( .A(n140), .B(n153), .C(n55), .D(n52), .ICI(n53), .S(n42), 
        .ICO(n40), .CO(n41) );
  CMPR42X1 U34 ( .A(n131), .B(n146), .C(n135), .D(n169), .ICI(n161), .S(n45), 
        .ICO(n43), .CO(n44) );
  CMPR42X1 U35 ( .A(n60), .B(n54), .C(n51), .D(n61), .ICI(n57), .S(n48), .ICO(
        n46), .CO(n47) );
  CMPR42X1 U36 ( .A(n154), .B(n162), .C(n63), .D(n65), .ICI(n56), .S(n51), 
        .ICO(n49), .CO(n50) );
  CMPR42X1 U37 ( .A(n132), .B(n177), .C(n147), .D(n141), .ICI(n170), .S(n54), 
        .ICO(n52), .CO(n53) );
  ADDHXL U38 ( .A(a[8]), .B(n136), .CO(n55), .S(n56) );
  CMPR42X1 U39 ( .A(n70), .B(n66), .C(n62), .D(n71), .ICI(n67), .S(n59), .ICO(
        n57), .CO(n58) );
  CMPR42X1 U40 ( .A(n155), .B(n163), .C(n73), .D(n75), .ICI(n64), .S(n62), 
        .ICO(n60), .CO(n61) );
  ADDFX2 U41 ( .A(n148), .B(n178), .CI(n171), .CO(n63), .S(n64) );
  ADDHXL U42 ( .A(n142), .B(n137), .CO(n65), .S(n66) );
  CMPR42X1 U43 ( .A(n76), .B(n74), .C(n72), .D(n81), .ICI(n77), .S(n69), .ICO(
        n67), .CO(n68) );
  CMPR42X1 U44 ( .A(n179), .B(n156), .C(n80), .D(n172), .ICI(n83), .S(n72), 
        .ICO(n70), .CO(n71) );
  ADDFX2 U45 ( .A(n185), .B(n164), .CI(n143), .CO(n73), .S(n74) );
  ADDHXL U46 ( .A(a[7]), .B(n149), .CO(n75), .S(n76) );
  CMPR42X1 U47 ( .A(n84), .B(n91), .C(n82), .D(n89), .ICI(n85), .S(n79), .ICO(
        n77), .CO(n78) );
  CMPR42X1 U48 ( .A(n180), .B(n165), .C(n150), .D(n173), .ICI(n88), .S(n82), 
        .ICO(n80), .CO(n81) );
  ADDHXL U49 ( .A(n157), .B(n186), .CO(n83), .S(n84) );
  CMPR42X1 U50 ( .A(n96), .B(n98), .C(n90), .D(n92), .ICI(n93), .S(n87), .ICO(
        n85), .CO(n86) );
  CMPR42X1 U51 ( .A(n158), .B(n192), .C(n181), .D(n174), .ICI(n187), .S(n90), 
        .ICO(n88), .CO(n89) );
  ADDHXL U52 ( .A(a[6]), .B(n166), .CO(n91), .S(n92) );
  CMPR42X1 U53 ( .A(n103), .B(n105), .C(n99), .D(n97), .ICI(n100), .S(n95), 
        .ICO(n93), .CO(n94) );
  ADDFX2 U54 ( .A(n182), .B(n193), .CI(n188), .CO(n96), .S(n97) );
  ADDHXL U55 ( .A(n175), .B(n167), .CO(n98), .S(n99) );
  CMPR42X1 U56 ( .A(n110), .B(n194), .C(n106), .D(n104), .ICI(n107), .S(n102), 
        .ICO(n100), .CO(n101) );
  ADDFX2 U57 ( .A(n176), .B(n198), .CI(n189), .CO(n103), .S(n104) );
  ADDHXL U58 ( .A(a[5]), .B(n183), .CO(n105), .S(n106) );
  CMPR42X1 U59 ( .A(n195), .B(n199), .C(n111), .D(n115), .ICI(n112), .S(n109), 
        .ICO(n107), .CO(n108) );
  ADDHXL U60 ( .A(n190), .B(n184), .CO(n110), .S(n111) );
  CMPR42X1 U61 ( .A(n191), .B(n203), .C(n119), .D(n200), .ICI(n116), .S(n114), 
        .ICO(n112), .CO(n113) );
  ADDHXL U62 ( .A(a[4]), .B(n196), .CO(n115), .S(n116) );
  ADDFX2 U63 ( .A(n123), .B(n201), .CI(n120), .CO(n117), .S(n118) );
  ADDHXL U64 ( .A(n204), .B(n197), .CO(n119), .S(n120) );
  ADDFX2 U65 ( .A(n202), .B(n205), .CI(n125), .CO(n121), .S(n122) );
  ADDHXL U66 ( .A(a[3]), .B(n207), .CO(n123), .S(n124) );
  ADDHXL U67 ( .A(n208), .B(n206), .CO(n125), .S(n126) );
  ADDHXL U68 ( .A(a[2]), .B(n210), .CO(n127), .S(n128) );
  CLKINVX3 U180 ( .A(n288), .Y(n291) );
  INVX1 U181 ( .A(n288), .Y(n292) );
  CLKINVX3 U182 ( .A(product[0]), .Y(n278) );
  CLKINVX3 U183 ( .A(n280), .Y(n282) );
  INVX1 U184 ( .A(n284), .Y(n287) );
  CLKINVX3 U185 ( .A(n293), .Y(n295) );
  CLKINVX3 U186 ( .A(n284), .Y(n286) );
  CLKINVX3 U187 ( .A(n296), .Y(n298) );
  CLKINVX3 U188 ( .A(n299), .Y(n301) );
  INVX1 U189 ( .A(n290), .Y(n288) );
  INVX1 U190 ( .A(n280), .Y(n283) );
  INVX1 U191 ( .A(product[0]), .Y(n279) );
  CLKINVX3 U192 ( .A(n302), .Y(n304) );
  INVX1 U193 ( .A(n277), .Y(product[0]) );
  INVX1 U194 ( .A(b[0]), .Y(n277) );
  INVX1 U195 ( .A(n281), .Y(n280) );
  INVX1 U196 ( .A(b[1]), .Y(n281) );
  INVX1 U197 ( .A(n285), .Y(n284) );
  INVX1 U198 ( .A(b[2]), .Y(n285) );
  INVX1 U199 ( .A(b[3]), .Y(n290) );
  INVX1 U200 ( .A(n297), .Y(n296) );
  INVX1 U201 ( .A(b[5]), .Y(n297) );
  INVX1 U202 ( .A(n300), .Y(n299) );
  INVX1 U203 ( .A(b[6]), .Y(n300) );
  INVX1 U204 ( .A(n294), .Y(n293) );
  INVX1 U205 ( .A(b[4]), .Y(n294) );
  INVX1 U206 ( .A(n303), .Y(n302) );
  INVX1 U207 ( .A(b[7]), .Y(n303) );
  CLKINVX3 U208 ( .A(b[8]), .Y(n312) );
  CLKINVX3 U209 ( .A(b[10]), .Y(n310) );
  CLKINVX3 U210 ( .A(b[11]), .Y(n309) );
  CLKINVX3 U211 ( .A(b[9]), .Y(n311) );
  CLKINVX3 U212 ( .A(b[12]), .Y(n308) );
  INVX1 U213 ( .A(b[13]), .Y(n307) );
  INVX1 U214 ( .A(b[14]), .Y(n306) );
  INVX1 U215 ( .A(b[15]), .Y(n305) );
  INVX1 U216 ( .A(n290), .Y(n289) );
  XOR2X1 U217 ( .A(n313), .B(n314), .Y(product[19]) );
  XOR2X1 U218 ( .A(n315), .B(n29), .Y(n314) );
  XOR2X1 U219 ( .A(n316), .B(n317), .Y(n315) );
  XOR2X1 U220 ( .A(n318), .B(n319), .Y(n317) );
  XOR2X1 U221 ( .A(n320), .B(n321), .Y(n319) );
  XNOR2X1 U222 ( .A(n28), .B(n2), .Y(n321) );
  NAND2X1 U223 ( .A(b[11]), .B(n302), .Y(n320) );
  XOR2X1 U224 ( .A(n322), .B(n323), .Y(n318) );
  NAND2X1 U225 ( .A(b[13]), .B(n296), .Y(n323) );
  NAND2X1 U226 ( .A(b[12]), .B(n299), .Y(n322) );
  XOR2X1 U227 ( .A(n324), .B(n325), .Y(n316) );
  XOR2X1 U228 ( .A(n326), .B(n327), .Y(n325) );
  NAND2X1 U229 ( .A(b[14]), .B(n293), .Y(n327) );
  NAND2X1 U230 ( .A(b[15]), .B(n289), .Y(n326) );
  XOR2X1 U231 ( .A(n328), .B(n34), .Y(n324) );
  NAND2X1 U232 ( .A(b[10]), .B(b[8]), .Y(n328) );
  XOR2X1 U233 ( .A(n329), .B(n31), .Y(n313) );
  XNOR2X1 U234 ( .A(n35), .B(n32), .Y(n329) );
  NOR2X1 U235 ( .A(n278), .B(n282), .Y(n212) );
  NOR2X1 U236 ( .A(n278), .B(n286), .Y(n211) );
  NOR2X1 U237 ( .A(n282), .B(n287), .Y(n210) );
  NOR2X1 U238 ( .A(n291), .B(n278), .Y(n209) );
  NOR2X1 U239 ( .A(n291), .B(n283), .Y(n208) );
  NOR2X1 U240 ( .A(n291), .B(n287), .Y(n207) );
  NOR2X1 U241 ( .A(n295), .B(n279), .Y(n206) );
  NOR2X1 U242 ( .A(n295), .B(n283), .Y(n205) );
  NOR2X1 U243 ( .A(n295), .B(n286), .Y(n204) );
  NOR2X1 U244 ( .A(n291), .B(n295), .Y(n203) );
  NOR2X1 U245 ( .A(n298), .B(n279), .Y(n202) );
  NOR2X1 U246 ( .A(n298), .B(n282), .Y(n201) );
  NOR2X1 U247 ( .A(n298), .B(n286), .Y(n200) );
  NOR2X1 U248 ( .A(n291), .B(n298), .Y(n199) );
  NOR2X1 U249 ( .A(n295), .B(n298), .Y(n198) );
  NOR2X1 U250 ( .A(n301), .B(n278), .Y(n197) );
  NOR2X1 U251 ( .A(n301), .B(n282), .Y(n196) );
  NOR2X1 U252 ( .A(n301), .B(n286), .Y(n195) );
  NOR2X1 U253 ( .A(n291), .B(n301), .Y(n194) );
  NOR2X1 U254 ( .A(n295), .B(n301), .Y(n193) );
  NOR2X1 U255 ( .A(n301), .B(n298), .Y(n192) );
  NOR2X1 U256 ( .A(n304), .B(n278), .Y(n191) );
  NOR2X1 U257 ( .A(n304), .B(n282), .Y(n190) );
  NOR2X1 U258 ( .A(n304), .B(n286), .Y(n189) );
  NOR2X1 U259 ( .A(n291), .B(n304), .Y(n188) );
  NOR2X1 U260 ( .A(n295), .B(n304), .Y(n187) );
  NOR2X1 U261 ( .A(n304), .B(n298), .Y(n186) );
  NOR2X1 U262 ( .A(n304), .B(n301), .Y(n185) );
  NOR2X1 U263 ( .A(n312), .B(n278), .Y(n184) );
  NOR2X1 U264 ( .A(n312), .B(n282), .Y(n183) );
  NOR2X1 U265 ( .A(n312), .B(n286), .Y(n182) );
  NOR2X1 U266 ( .A(n312), .B(n292), .Y(n181) );
  NOR2X1 U267 ( .A(n312), .B(n295), .Y(n180) );
  NOR2X1 U268 ( .A(n312), .B(n298), .Y(n179) );
  NOR2X1 U269 ( .A(n312), .B(n301), .Y(n178) );
  NOR2X1 U270 ( .A(n312), .B(n304), .Y(n177) );
  NOR2X1 U271 ( .A(n278), .B(n311), .Y(n176) );
  NOR2X1 U272 ( .A(n282), .B(n311), .Y(n175) );
  NOR2X1 U273 ( .A(n286), .B(n311), .Y(n174) );
  NOR2X1 U274 ( .A(n291), .B(n311), .Y(n173) );
  NOR2X1 U275 ( .A(n295), .B(n311), .Y(n172) );
  NOR2X1 U276 ( .A(n298), .B(n311), .Y(n171) );
  NOR2X1 U277 ( .A(n301), .B(n311), .Y(n170) );
  NOR2X1 U278 ( .A(n304), .B(n311), .Y(n169) );
  NOR2X1 U279 ( .A(n312), .B(n311), .Y(n168) );
  NOR2X1 U280 ( .A(n310), .B(n278), .Y(n167) );
  NOR2X1 U281 ( .A(n310), .B(n282), .Y(n166) );
  NOR2X1 U282 ( .A(n310), .B(n286), .Y(n165) );
  NOR2X1 U283 ( .A(n310), .B(n292), .Y(n164) );
  NOR2X1 U284 ( .A(n310), .B(n295), .Y(n163) );
  NOR2X1 U285 ( .A(n310), .B(n298), .Y(n162) );
  NOR2X1 U286 ( .A(n310), .B(n301), .Y(n161) );
  NOR2X1 U287 ( .A(n310), .B(n304), .Y(n160) );
  NOR2X1 U288 ( .A(n309), .B(n278), .Y(n158) );
  NOR2X1 U289 ( .A(n309), .B(n282), .Y(n157) );
  NOR2X1 U290 ( .A(n309), .B(n286), .Y(n156) );
  NOR2X1 U291 ( .A(n291), .B(n309), .Y(n155) );
  NOR2X1 U292 ( .A(n295), .B(n309), .Y(n154) );
  NOR2X1 U293 ( .A(n309), .B(n298), .Y(n153) );
  NOR2X1 U294 ( .A(n309), .B(n301), .Y(n152) );
  NOR2X1 U295 ( .A(n308), .B(n278), .Y(n150) );
  NOR2X1 U296 ( .A(n308), .B(n282), .Y(n149) );
  NOR2X1 U297 ( .A(n308), .B(n286), .Y(n148) );
  NOR2X1 U298 ( .A(n291), .B(n308), .Y(n147) );
  NOR2X1 U299 ( .A(n295), .B(n308), .Y(n146) );
  NOR2X1 U300 ( .A(n308), .B(n298), .Y(n145) );
  NOR2X1 U301 ( .A(n307), .B(n278), .Y(n143) );
  NOR2X1 U302 ( .A(n307), .B(n282), .Y(n142) );
  NOR2X1 U303 ( .A(n307), .B(n286), .Y(n141) );
  NOR2X1 U304 ( .A(n291), .B(n307), .Y(n140) );
  NOR2X1 U305 ( .A(n295), .B(n307), .Y(n139) );
  NOR2X1 U306 ( .A(n306), .B(n278), .Y(n137) );
  NOR2X1 U307 ( .A(n306), .B(n282), .Y(n136) );
  NOR2X1 U308 ( .A(n306), .B(n286), .Y(n135) );
  NOR2X1 U309 ( .A(n291), .B(n306), .Y(n134) );
  NOR2X1 U310 ( .A(n305), .B(n278), .Y(n132) );
  NOR2X1 U311 ( .A(n305), .B(n282), .Y(n131) );
  NOR2X1 U312 ( .A(n305), .B(n286), .Y(n130) );
endmodule


module Control_And_Registers_DW_mult_uns_1 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n130,
         n131, n132, n134, n135, n136, n137, n139, n140, n141, n142, n143,
         n145, n146, n147, n148, n149, n150, n152, n153, n154, n155, n156,
         n157, n158, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334;

  ADDFX2 U3 ( .A(n30), .B(n38), .CI(n3), .CO(n2), .S(product[18]) );
  ADDFX2 U4 ( .A(n39), .B(n47), .CI(n4), .CO(n3), .S(product[17]) );
  ADDFX2 U5 ( .A(n48), .B(n58), .CI(n5), .CO(n4), .S(product[16]) );
  ADDFX2 U6 ( .A(n59), .B(n68), .CI(n6), .CO(n5), .S(product[15]) );
  ADDFX2 U7 ( .A(n69), .B(n78), .CI(n7), .CO(n6), .S(product[14]) );
  ADDFX2 U8 ( .A(n79), .B(n86), .CI(n8), .CO(n7), .S(product[13]) );
  ADDFX2 U9 ( .A(n87), .B(n94), .CI(n9), .CO(n8), .S(product[12]) );
  ADDFX2 U10 ( .A(n95), .B(n101), .CI(n10), .CO(n9), .S(product[11]) );
  ADDFX2 U11 ( .A(n102), .B(n108), .CI(n11), .CO(n10), .S(product[10]) );
  ADDFX2 U12 ( .A(n109), .B(n113), .CI(n12), .CO(n11), .S(product[9]) );
  ADDFX2 U13 ( .A(n114), .B(n117), .CI(n13), .CO(n12), .S(product[8]) );
  ADDFX2 U14 ( .A(n118), .B(n121), .CI(n14), .CO(n13), .S(product[7]) );
  ADDFX2 U15 ( .A(n122), .B(n124), .CI(n15), .CO(n14), .S(product[6]) );
  ADDFX2 U16 ( .A(n126), .B(n127), .CI(n16), .CO(n15), .S(product[5]) );
  ADDFX2 U17 ( .A(n128), .B(n209), .CI(n17), .CO(n16), .S(product[4]) );
  ADDHXL U18 ( .A(n211), .B(n18), .CO(n17), .S(product[3]) );
  ADDHXL U19 ( .A(n281), .B(n212), .CO(n18), .S(product[2]) );
  CMPR42X1 U29 ( .A(n40), .B(n44), .C(n33), .D(n41), .ICI(n37), .S(n30), .ICO(
        n28), .CO(n29) );
  CMPR42X1 U30 ( .A(n152), .B(n130), .C(n43), .D(n145), .ICI(n36), .S(n33), 
        .ICO(n31), .CO(n32) );
  CMPR42X1 U31 ( .A(n134), .B(a[9]), .C(n160), .D(n168), .ICI(n139), .S(n36), 
        .ICO(n34), .CO(n35) );
  CMPR42X1 U32 ( .A(n49), .B(n45), .C(n42), .D(n50), .ICI(n46), .S(n39), .ICO(
        n37), .CO(n38) );
  CMPR42X1 U33 ( .A(n140), .B(n153), .C(n55), .D(n52), .ICI(n53), .S(n42), 
        .ICO(n40), .CO(n41) );
  CMPR42X1 U34 ( .A(n131), .B(n146), .C(n135), .D(n169), .ICI(n161), .S(n45), 
        .ICO(n43), .CO(n44) );
  CMPR42X1 U35 ( .A(n60), .B(n54), .C(n51), .D(n61), .ICI(n57), .S(n48), .ICO(
        n46), .CO(n47) );
  CMPR42X1 U36 ( .A(n154), .B(n162), .C(n63), .D(n65), .ICI(n56), .S(n51), 
        .ICO(n49), .CO(n50) );
  CMPR42X1 U37 ( .A(n132), .B(n177), .C(n147), .D(n141), .ICI(n170), .S(n54), 
        .ICO(n52), .CO(n53) );
  ADDHXL U38 ( .A(a[8]), .B(n136), .CO(n55), .S(n56) );
  CMPR42X1 U39 ( .A(n70), .B(n66), .C(n62), .D(n71), .ICI(n67), .S(n59), .ICO(
        n57), .CO(n58) );
  CMPR42X1 U40 ( .A(n155), .B(n163), .C(n73), .D(n75), .ICI(n64), .S(n62), 
        .ICO(n60), .CO(n61) );
  ADDFX2 U41 ( .A(n148), .B(n178), .CI(n171), .CO(n63), .S(n64) );
  ADDHXL U42 ( .A(n142), .B(n137), .CO(n65), .S(n66) );
  CMPR42X1 U43 ( .A(n76), .B(n74), .C(n72), .D(n81), .ICI(n77), .S(n69), .ICO(
        n67), .CO(n68) );
  CMPR42X1 U44 ( .A(n179), .B(n156), .C(n80), .D(n172), .ICI(n83), .S(n72), 
        .ICO(n70), .CO(n71) );
  ADDFX2 U45 ( .A(n185), .B(n164), .CI(n143), .CO(n73), .S(n74) );
  ADDHXL U46 ( .A(n306), .B(n149), .CO(n75), .S(n76) );
  CMPR42X1 U47 ( .A(n84), .B(n91), .C(n82), .D(n89), .ICI(n85), .S(n79), .ICO(
        n77), .CO(n78) );
  CMPR42X1 U48 ( .A(n180), .B(n165), .C(n150), .D(n173), .ICI(n88), .S(n82), 
        .ICO(n80), .CO(n81) );
  ADDHXL U49 ( .A(n157), .B(n186), .CO(n83), .S(n84) );
  CMPR42X1 U50 ( .A(n96), .B(n98), .C(n90), .D(n92), .ICI(n93), .S(n87), .ICO(
        n85), .CO(n86) );
  CMPR42X1 U51 ( .A(n158), .B(n192), .C(n181), .D(n174), .ICI(n187), .S(n90), 
        .ICO(n88), .CO(n89) );
  ADDHXL U52 ( .A(n302), .B(n166), .CO(n91), .S(n92) );
  CMPR42X1 U53 ( .A(n103), .B(n105), .C(n99), .D(n97), .ICI(n100), .S(n95), 
        .ICO(n93), .CO(n94) );
  ADDFX2 U54 ( .A(n182), .B(n193), .CI(n188), .CO(n96), .S(n97) );
  ADDHXL U55 ( .A(n175), .B(n167), .CO(n98), .S(n99) );
  CMPR42X1 U56 ( .A(n110), .B(n194), .C(n106), .D(n104), .ICI(n107), .S(n102), 
        .ICO(n100), .CO(n101) );
  ADDFX2 U57 ( .A(n176), .B(n198), .CI(n189), .CO(n103), .S(n104) );
  ADDHXL U58 ( .A(n298), .B(n183), .CO(n105), .S(n106) );
  CMPR42X1 U59 ( .A(n195), .B(n199), .C(n111), .D(n115), .ICI(n112), .S(n109), 
        .ICO(n107), .CO(n108) );
  ADDHXL U60 ( .A(n190), .B(n184), .CO(n110), .S(n111) );
  CMPR42X1 U61 ( .A(n191), .B(n203), .C(n119), .D(n200), .ICI(n116), .S(n114), 
        .ICO(n112), .CO(n113) );
  ADDHXL U62 ( .A(n295), .B(n196), .CO(n115), .S(n116) );
  ADDFX2 U63 ( .A(n123), .B(n201), .CI(n120), .CO(n117), .S(n118) );
  ADDHXL U64 ( .A(n204), .B(n197), .CO(n119), .S(n120) );
  ADDFX2 U65 ( .A(n202), .B(n205), .CI(n125), .CO(n121), .S(n122) );
  ADDHXL U66 ( .A(n291), .B(n207), .CO(n123), .S(n124) );
  ADDHXL U67 ( .A(n208), .B(n206), .CO(n125), .S(n126) );
  ADDHXL U68 ( .A(n286), .B(n210), .CO(n127), .S(n128) );
  CLKINVX3 U180 ( .A(n280), .Y(n283) );
  INVX1 U181 ( .A(n285), .Y(n289) );
  CLKINVX3 U182 ( .A(n295), .Y(n297) );
  CLKINVX3 U183 ( .A(n285), .Y(n288) );
  CLKINVX3 U184 ( .A(n290), .Y(n293) );
  CLKINVX3 U185 ( .A(n298), .Y(n301) );
  CLKINVX3 U186 ( .A(n302), .Y(n305) );
  INVX1 U187 ( .A(n280), .Y(n284) );
  CLKINVX3 U188 ( .A(n306), .Y(n309) );
  INVX1 U189 ( .A(n290), .Y(n294) );
  INVX1 U190 ( .A(n287), .Y(n286) );
  INVX1 U191 ( .A(n282), .Y(n281) );
  CLKINVX3 U192 ( .A(product[0]), .Y(n278) );
  INVX1 U193 ( .A(n282), .Y(n280) );
  INVX1 U194 ( .A(n287), .Y(n285) );
  INVX1 U195 ( .A(n292), .Y(n290) );
  INVX1 U196 ( .A(n296), .Y(n295) );
  INVX1 U197 ( .A(n300), .Y(n298) );
  INVX1 U198 ( .A(n304), .Y(n302) );
  INVX1 U199 ( .A(product[0]), .Y(n279) );
  INVX1 U200 ( .A(n308), .Y(n306) );
  INVX1 U201 ( .A(n292), .Y(n291) );
  INVX1 U202 ( .A(n300), .Y(n299) );
  INVX1 U203 ( .A(n277), .Y(product[0]) );
  INVX1 U204 ( .A(a[0]), .Y(n277) );
  INVX1 U205 ( .A(a[1]), .Y(n282) );
  INVX1 U206 ( .A(a[2]), .Y(n287) );
  INVX1 U207 ( .A(a[3]), .Y(n292) );
  INVX1 U208 ( .A(a[5]), .Y(n300) );
  INVX1 U209 ( .A(a[6]), .Y(n304) );
  INVX1 U210 ( .A(a[4]), .Y(n296) );
  INVX1 U211 ( .A(a[7]), .Y(n308) );
  INVX1 U212 ( .A(n308), .Y(n307) );
  CLKINVX3 U213 ( .A(a[8]), .Y(n317) );
  CLKINVX3 U214 ( .A(a[10]), .Y(n315) );
  CLKINVX3 U215 ( .A(a[11]), .Y(n314) );
  CLKINVX3 U216 ( .A(a[9]), .Y(n316) );
  CLKINVX3 U217 ( .A(a[12]), .Y(n313) );
  INVX1 U218 ( .A(a[13]), .Y(n312) );
  INVX1 U219 ( .A(a[14]), .Y(n311) );
  INVX1 U220 ( .A(a[15]), .Y(n310) );
  NAND2BX1 U221 ( .AN(n296), .B(a[14]), .Y(n332) );
  INVX1 U222 ( .A(n304), .Y(n303) );
  XOR2X1 U223 ( .A(n318), .B(n319), .Y(product[19]) );
  XOR2X1 U224 ( .A(n320), .B(n29), .Y(n319) );
  XOR2X1 U225 ( .A(n321), .B(n322), .Y(n320) );
  XOR2X1 U226 ( .A(n323), .B(n324), .Y(n322) );
  XOR2X1 U227 ( .A(n325), .B(n326), .Y(n324) );
  XNOR2X1 U228 ( .A(n28), .B(n2), .Y(n326) );
  NAND2X1 U229 ( .A(n307), .B(a[11]), .Y(n325) );
  XOR2X1 U230 ( .A(n327), .B(n328), .Y(n323) );
  NAND2X1 U231 ( .A(n299), .B(a[13]), .Y(n328) );
  NAND2X1 U232 ( .A(n303), .B(a[12]), .Y(n327) );
  XOR2X1 U233 ( .A(n329), .B(n330), .Y(n321) );
  XOR2X1 U234 ( .A(n331), .B(n332), .Y(n330) );
  NAND2X1 U235 ( .A(n291), .B(a[15]), .Y(n331) );
  XOR2X1 U236 ( .A(n333), .B(n34), .Y(n329) );
  NAND2X1 U237 ( .A(a[8]), .B(a[10]), .Y(n333) );
  XOR2X1 U238 ( .A(n334), .B(n31), .Y(n318) );
  XNOR2X1 U239 ( .A(n35), .B(n32), .Y(n334) );
  NOR2X1 U240 ( .A(n278), .B(n283), .Y(n212) );
  NOR2X1 U241 ( .A(n278), .B(n288), .Y(n211) );
  NOR2X1 U242 ( .A(n283), .B(n289), .Y(n210) );
  NOR2X1 U243 ( .A(n293), .B(n278), .Y(n209) );
  NOR2X1 U244 ( .A(n293), .B(n284), .Y(n208) );
  NOR2X1 U245 ( .A(n293), .B(n289), .Y(n207) );
  NOR2X1 U246 ( .A(n297), .B(n279), .Y(n206) );
  NOR2X1 U247 ( .A(n297), .B(n284), .Y(n205) );
  NOR2X1 U248 ( .A(n297), .B(n288), .Y(n204) );
  NOR2X1 U249 ( .A(n293), .B(n297), .Y(n203) );
  NOR2X1 U250 ( .A(n301), .B(n279), .Y(n202) );
  NOR2X1 U251 ( .A(n301), .B(n283), .Y(n201) );
  NOR2X1 U252 ( .A(n301), .B(n288), .Y(n200) );
  NOR2X1 U253 ( .A(n293), .B(n301), .Y(n199) );
  NOR2X1 U254 ( .A(n297), .B(n301), .Y(n198) );
  NOR2X1 U255 ( .A(n305), .B(n278), .Y(n197) );
  NOR2X1 U256 ( .A(n305), .B(n283), .Y(n196) );
  NOR2X1 U257 ( .A(n305), .B(n288), .Y(n195) );
  NOR2X1 U258 ( .A(n293), .B(n305), .Y(n194) );
  NOR2X1 U259 ( .A(n297), .B(n305), .Y(n193) );
  NOR2X1 U260 ( .A(n305), .B(n301), .Y(n192) );
  NOR2X1 U261 ( .A(n309), .B(n278), .Y(n191) );
  NOR2X1 U262 ( .A(n309), .B(n283), .Y(n190) );
  NOR2X1 U263 ( .A(n309), .B(n288), .Y(n189) );
  NOR2X1 U264 ( .A(n293), .B(n309), .Y(n188) );
  NOR2X1 U265 ( .A(n297), .B(n309), .Y(n187) );
  NOR2X1 U266 ( .A(n309), .B(n301), .Y(n186) );
  NOR2X1 U267 ( .A(n309), .B(n305), .Y(n185) );
  NOR2X1 U268 ( .A(n317), .B(n278), .Y(n184) );
  NOR2X1 U269 ( .A(n317), .B(n283), .Y(n183) );
  NOR2X1 U270 ( .A(n317), .B(n288), .Y(n182) );
  NOR2X1 U271 ( .A(n317), .B(n294), .Y(n181) );
  NOR2X1 U272 ( .A(n317), .B(n297), .Y(n180) );
  NOR2X1 U273 ( .A(n317), .B(n301), .Y(n179) );
  NOR2X1 U274 ( .A(n317), .B(n305), .Y(n178) );
  NOR2X1 U275 ( .A(n317), .B(n309), .Y(n177) );
  NOR2X1 U276 ( .A(n278), .B(n316), .Y(n176) );
  NOR2X1 U277 ( .A(n283), .B(n316), .Y(n175) );
  NOR2X1 U278 ( .A(n288), .B(n316), .Y(n174) );
  NOR2X1 U279 ( .A(n293), .B(n316), .Y(n173) );
  NOR2X1 U280 ( .A(n297), .B(n316), .Y(n172) );
  NOR2X1 U281 ( .A(n301), .B(n316), .Y(n171) );
  NOR2X1 U282 ( .A(n305), .B(n316), .Y(n170) );
  NOR2X1 U283 ( .A(n309), .B(n316), .Y(n169) );
  NOR2X1 U284 ( .A(n317), .B(n316), .Y(n168) );
  NOR2X1 U285 ( .A(n315), .B(n278), .Y(n167) );
  NOR2X1 U286 ( .A(n315), .B(n283), .Y(n166) );
  NOR2X1 U287 ( .A(n315), .B(n288), .Y(n165) );
  NOR2X1 U288 ( .A(n315), .B(n294), .Y(n164) );
  NOR2X1 U289 ( .A(n315), .B(n297), .Y(n163) );
  NOR2X1 U290 ( .A(n315), .B(n301), .Y(n162) );
  NOR2X1 U291 ( .A(n315), .B(n305), .Y(n161) );
  NOR2X1 U292 ( .A(n315), .B(n309), .Y(n160) );
  NOR2X1 U293 ( .A(n314), .B(n278), .Y(n158) );
  NOR2X1 U294 ( .A(n314), .B(n283), .Y(n157) );
  NOR2X1 U295 ( .A(n314), .B(n288), .Y(n156) );
  NOR2X1 U296 ( .A(n293), .B(n314), .Y(n155) );
  NOR2X1 U297 ( .A(n297), .B(n314), .Y(n154) );
  NOR2X1 U298 ( .A(n314), .B(n301), .Y(n153) );
  NOR2X1 U299 ( .A(n314), .B(n305), .Y(n152) );
  NOR2X1 U300 ( .A(n313), .B(n278), .Y(n150) );
  NOR2X1 U301 ( .A(n313), .B(n283), .Y(n149) );
  NOR2X1 U302 ( .A(n313), .B(n288), .Y(n148) );
  NOR2X1 U303 ( .A(n293), .B(n313), .Y(n147) );
  NOR2X1 U304 ( .A(n297), .B(n313), .Y(n146) );
  NOR2X1 U305 ( .A(n313), .B(n301), .Y(n145) );
  NOR2X1 U306 ( .A(n312), .B(n278), .Y(n143) );
  NOR2X1 U307 ( .A(n312), .B(n283), .Y(n142) );
  NOR2X1 U308 ( .A(n312), .B(n288), .Y(n141) );
  NOR2X1 U309 ( .A(n293), .B(n312), .Y(n140) );
  NOR2X1 U310 ( .A(n297), .B(n312), .Y(n139) );
  NOR2X1 U311 ( .A(n311), .B(n278), .Y(n137) );
  NOR2X1 U312 ( .A(n311), .B(n283), .Y(n136) );
  NOR2X1 U313 ( .A(n311), .B(n288), .Y(n135) );
  NOR2X1 U314 ( .A(n293), .B(n311), .Y(n134) );
  NOR2X1 U315 ( .A(n310), .B(n278), .Y(n132) );
  NOR2X1 U316 ( .A(n310), .B(n283), .Y(n131) );
  NOR2X1 U317 ( .A(n310), .B(n288), .Y(n130) );
endmodule


module Control_And_Registers_DW01_add_18 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR3X2 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .Y(SUM[9]) );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X2 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module Control_And_Registers_DW01_add_17 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  XOR3X2 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .Y(SUM[9]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X2 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module Control_And_Registers_DW_mult_uns_0 ( a, b, product );
  input [9:0] a;
  input [9:0] b;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n73, n75,
         n76, n78, n79, n80, n82, n83, n84, n85, n87, n88, n89, n90, n91, n93,
         n94, n95, n96, n97, n98, n100, n101, n102, n103, n104, n105, n106,
         n108, n109, n110, n111, n112, n113, n114, n115, n117, n118, n119,
         n120, n121, n122, n123, n124, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222;

  ADDFX2 U3 ( .A(n26), .B(n36), .CI(n3), .CO(n2), .S(product[8]) );
  ADDFX2 U4 ( .A(n37), .B(n46), .CI(n4), .CO(n3), .S(product[7]) );
  ADDFX2 U5 ( .A(n47), .B(n54), .CI(n5), .CO(n4), .S(product[6]) );
  ADDFX2 U6 ( .A(n55), .B(n61), .CI(n6), .CO(n5), .S(product[5]) );
  ADDFX2 U7 ( .A(n62), .B(n65), .CI(n7), .CO(n6), .S(product[4]) );
  ADDFX2 U8 ( .A(n66), .B(n68), .CI(n8), .CO(n7), .S(product[3]) );
  ADDFX2 U9 ( .A(n9), .B(n106), .CI(n70), .CO(n8), .S(product[2]) );
  ADDHXL U10 ( .A(n115), .B(n124), .CO(n9), .S(product[1]) );
  CMPR42X1 U25 ( .A(n38), .B(n32), .C(n29), .D(n39), .ICI(n35), .S(n26), .ICO(
        n24), .CO(n25) );
  CMPR42X1 U26 ( .A(n93), .B(n100), .C(n41), .D(n43), .ICI(n34), .S(n29), 
        .ICO(n27), .CO(n28) );
  CMPR42X1 U27 ( .A(n78), .B(n117), .C(n87), .D(n82), .ICI(n108), .S(n32), 
        .ICO(n30), .CO(n31) );
  ADDHXL U28 ( .A(n75), .B(n73), .CO(n33), .S(n34) );
  CMPR42X1 U29 ( .A(n44), .B(n42), .C(n40), .D(n49), .ICI(n45), .S(n37), .ICO(
        n35), .CO(n36) );
  CMPR42X1 U30 ( .A(n109), .B(n88), .C(n48), .D(n101), .ICI(n51), .S(n40), 
        .ICO(n38), .CO(n39) );
  ADDFX2 U31 ( .A(n118), .B(n94), .CI(n83), .CO(n41), .S(n42) );
  ADDHXL U32 ( .A(n79), .B(n76), .CO(n43), .S(n44) );
  CMPR42X1 U33 ( .A(n56), .B(n58), .C(n50), .D(n52), .ICI(n53), .S(n47), .ICO(
        n45), .CO(n46) );
  CMPR42X1 U34 ( .A(n89), .B(n119), .C(n102), .D(n95), .ICI(n110), .S(n50), 
        .ICO(n48), .CO(n49) );
  ADDHXL U35 ( .A(n84), .B(n80), .CO(n51), .S(n52) );
  CMPR42X1 U36 ( .A(n63), .B(n111), .C(n59), .D(n57), .ICI(n60), .S(n55), 
        .ICO(n53), .CO(n54) );
  ADDFX2 U37 ( .A(n96), .B(n120), .CI(n103), .CO(n56), .S(n57) );
  ADDHXL U38 ( .A(n90), .B(n85), .CO(n58), .S(n59) );
  CMPR42X1 U39 ( .A(n104), .B(n121), .C(n67), .D(n112), .ICI(n64), .S(n62), 
        .ICO(n60), .CO(n61) );
  ADDHXL U40 ( .A(n97), .B(n91), .CO(n63), .S(n64) );
  ADDFX2 U41 ( .A(n113), .B(n122), .CI(n69), .CO(n65), .S(n66) );
  ADDHXL U42 ( .A(n105), .B(n98), .CO(n67), .S(n68) );
  ADDHXL U43 ( .A(n123), .B(n114), .CO(n69), .S(n70) );
  NAND2XL U121 ( .A(b[9]), .B(a[0]), .Y(n219) );
  CLKINVX2 U122 ( .A(a[0]), .Y(n189) );
  CLKINVX3 U123 ( .A(n179), .Y(n181) );
  INVX1 U124 ( .A(n180), .Y(n179) );
  INVX1 U125 ( .A(b[0]), .Y(n180) );
  CLKINVX3 U126 ( .A(b[1]), .Y(n188) );
  CLKINVX3 U127 ( .A(b[2]), .Y(n187) );
  NOR2BX1 U128 ( .AN(a[8]), .B(n180), .Y(n73) );
  CLKINVX3 U129 ( .A(a[1]), .Y(n190) );
  CLKINVX3 U130 ( .A(a[2]), .Y(n191) );
  CLKINVX3 U131 ( .A(b[3]), .Y(n186) );
  CLKINVX3 U132 ( .A(a[3]), .Y(n192) );
  INVX1 U133 ( .A(b[5]), .Y(n184) );
  INVX1 U134 ( .A(b[4]), .Y(n185) );
  CLKINVX3 U135 ( .A(a[4]), .Y(n193) );
  INVX1 U136 ( .A(a[5]), .Y(n194) );
  INVX1 U137 ( .A(a[6]), .Y(n195) );
  INVX1 U138 ( .A(b[6]), .Y(n183) );
  INVX1 U139 ( .A(b[7]), .Y(n182) );
  INVX1 U140 ( .A(a[7]), .Y(n196) );
  XOR2X1 U141 ( .A(n197), .B(n198), .Y(product[9]) );
  XOR2X1 U142 ( .A(n199), .B(n200), .Y(n198) );
  XOR2X1 U143 ( .A(n201), .B(n202), .Y(n200) );
  NOR2X1 U144 ( .A(n193), .B(n184), .Y(n202) );
  NAND2X1 U145 ( .A(b[6]), .B(a[3]), .Y(n201) );
  XOR2X1 U146 ( .A(n203), .B(n204), .Y(n199) );
  XOR2X1 U147 ( .A(n205), .B(n206), .Y(n204) );
  XOR2X1 U148 ( .A(n207), .B(n208), .Y(n206) );
  NAND2X1 U149 ( .A(n179), .B(a[9]), .Y(n208) );
  NAND2X1 U150 ( .A(b[1]), .B(a[8]), .Y(n207) );
  XOR2X1 U151 ( .A(n28), .B(n24), .Y(n205) );
  XOR2X1 U152 ( .A(n209), .B(n210), .Y(n203) );
  XOR2X1 U153 ( .A(n211), .B(n212), .Y(n210) );
  NAND2X1 U154 ( .A(b[7]), .B(a[2]), .Y(n212) );
  NAND2X1 U155 ( .A(b[4]), .B(a[5]), .Y(n211) );
  XOR2X1 U156 ( .A(n213), .B(n214), .Y(n209) );
  XOR2X1 U157 ( .A(n215), .B(n216), .Y(n214) );
  XNOR2X1 U158 ( .A(n30), .B(n27), .Y(n216) );
  XNOR2X1 U159 ( .A(n33), .B(n31), .Y(n215) );
  XOR2X1 U160 ( .A(n217), .B(n218), .Y(n213) );
  XOR2X1 U161 ( .A(n219), .B(n220), .Y(n218) );
  NAND2X1 U162 ( .A(b[8]), .B(a[1]), .Y(n220) );
  NAND2X1 U163 ( .A(b[2]), .B(a[7]), .Y(n217) );
  XOR2X1 U164 ( .A(n221), .B(n222), .Y(n197) );
  XNOR2X1 U165 ( .A(n25), .B(n2), .Y(n222) );
  NAND2X1 U166 ( .A(b[3]), .B(a[6]), .Y(n221) );
  NOR2X1 U167 ( .A(n181), .B(n189), .Y(product[0]) );
  NOR2X1 U168 ( .A(n192), .B(n181), .Y(n98) );
  NOR2X1 U169 ( .A(n192), .B(n188), .Y(n97) );
  NOR2X1 U170 ( .A(n192), .B(n187), .Y(n96) );
  NOR2X1 U171 ( .A(n186), .B(n192), .Y(n95) );
  NOR2X1 U172 ( .A(n192), .B(n185), .Y(n94) );
  NOR2X1 U173 ( .A(n184), .B(n192), .Y(n93) );
  NOR2X1 U174 ( .A(n193), .B(n181), .Y(n91) );
  NOR2X1 U175 ( .A(n193), .B(n188), .Y(n90) );
  NOR2X1 U176 ( .A(n193), .B(n187), .Y(n89) );
  NOR2X1 U177 ( .A(n186), .B(n193), .Y(n88) );
  NOR2X1 U178 ( .A(n193), .B(n185), .Y(n87) );
  NOR2X1 U179 ( .A(n194), .B(n181), .Y(n85) );
  NOR2X1 U180 ( .A(n194), .B(n188), .Y(n84) );
  NOR2X1 U181 ( .A(n194), .B(n187), .Y(n83) );
  NOR2X1 U182 ( .A(n186), .B(n194), .Y(n82) );
  NOR2X1 U183 ( .A(n195), .B(n181), .Y(n80) );
  NOR2X1 U184 ( .A(n195), .B(n188), .Y(n79) );
  NOR2X1 U185 ( .A(n195), .B(n187), .Y(n78) );
  NOR2X1 U186 ( .A(n181), .B(n196), .Y(n76) );
  NOR2X1 U187 ( .A(n188), .B(n196), .Y(n75) );
  NOR2X1 U188 ( .A(n188), .B(n189), .Y(n124) );
  NOR2X1 U189 ( .A(n187), .B(n189), .Y(n123) );
  NOR2X1 U190 ( .A(n186), .B(n189), .Y(n122) );
  NOR2X1 U191 ( .A(n185), .B(n189), .Y(n121) );
  NOR2X1 U192 ( .A(n184), .B(n189), .Y(n120) );
  NOR2X1 U193 ( .A(n183), .B(n189), .Y(n119) );
  NOR2X1 U194 ( .A(n182), .B(n189), .Y(n118) );
  AND2X1 U195 ( .A(b[8]), .B(a[0]), .Y(n117) );
  NOR2X1 U196 ( .A(n181), .B(n190), .Y(n115) );
  NOR2X1 U197 ( .A(n188), .B(n190), .Y(n114) );
  NOR2X1 U198 ( .A(n187), .B(n190), .Y(n113) );
  NOR2X1 U199 ( .A(n186), .B(n190), .Y(n112) );
  NOR2X1 U200 ( .A(n185), .B(n190), .Y(n111) );
  NOR2X1 U201 ( .A(n184), .B(n190), .Y(n110) );
  NOR2X1 U202 ( .A(n183), .B(n190), .Y(n109) );
  NOR2X1 U203 ( .A(n182), .B(n190), .Y(n108) );
  NOR2X1 U204 ( .A(n191), .B(n181), .Y(n106) );
  NOR2X1 U205 ( .A(n191), .B(n188), .Y(n105) );
  NOR2X1 U206 ( .A(n191), .B(n187), .Y(n104) );
  NOR2X1 U207 ( .A(n186), .B(n191), .Y(n103) );
  NOR2X1 U208 ( .A(n185), .B(n191), .Y(n102) );
  NOR2X1 U209 ( .A(n184), .B(n191), .Y(n101) );
  NOR2X1 U210 ( .A(n183), .B(n191), .Y(n100) );
endmodule


module Control_And_Registers_DW_div_uns_5 ( a, b, quotient, remainder, 
        divide_by_0 );
  input [19:0] a;
  input [19:0] b;
  output [19:0] quotient;
  output [19:0] remainder;
  output divide_by_0;
  wire   \u_div/SumTmp[1][0] , \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] , \u_div/SumTmp[1][5] ,
         \u_div/SumTmp[1][6] , \u_div/SumTmp[1][7] , \u_div/SumTmp[1][8] ,
         \u_div/SumTmp[1][9] , \u_div/SumTmp[1][10] , \u_div/SumTmp[1][11] ,
         \u_div/SumTmp[1][12] , \u_div/SumTmp[1][13] , \u_div/SumTmp[1][14] ,
         \u_div/SumTmp[1][15] , \u_div/SumTmp[1][16] , \u_div/SumTmp[1][17] ,
         \u_div/SumTmp[1][18] , \u_div/SumTmp[2][0] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[2][5] , \u_div/SumTmp[2][6] , \u_div/SumTmp[2][7] ,
         \u_div/SumTmp[2][8] , \u_div/SumTmp[2][9] , \u_div/SumTmp[2][10] ,
         \u_div/SumTmp[2][11] , \u_div/SumTmp[2][12] , \u_div/SumTmp[2][13] ,
         \u_div/SumTmp[2][14] , \u_div/SumTmp[2][15] , \u_div/SumTmp[2][16] ,
         \u_div/SumTmp[2][17] , \u_div/SumTmp[3][0] , \u_div/SumTmp[3][1] ,
         \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] , \u_div/SumTmp[3][4] ,
         \u_div/SumTmp[3][5] , \u_div/SumTmp[3][6] , \u_div/SumTmp[3][7] ,
         \u_div/SumTmp[3][8] , \u_div/SumTmp[3][9] , \u_div/SumTmp[3][10] ,
         \u_div/SumTmp[3][11] , \u_div/SumTmp[3][12] , \u_div/SumTmp[3][13] ,
         \u_div/SumTmp[3][14] , \u_div/SumTmp[3][15] , \u_div/SumTmp[3][16] ,
         \u_div/SumTmp[4][0] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[4][5] ,
         \u_div/SumTmp[4][6] , \u_div/SumTmp[4][7] , \u_div/SumTmp[4][8] ,
         \u_div/SumTmp[4][9] , \u_div/SumTmp[4][10] , \u_div/SumTmp[4][11] ,
         \u_div/SumTmp[4][12] , \u_div/SumTmp[4][13] , \u_div/SumTmp[4][14] ,
         \u_div/SumTmp[4][15] , \u_div/SumTmp[5][0] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] ,
         \u_div/SumTmp[5][5] , \u_div/SumTmp[5][6] , \u_div/SumTmp[5][7] ,
         \u_div/SumTmp[5][8] , \u_div/SumTmp[5][9] , \u_div/SumTmp[5][10] ,
         \u_div/SumTmp[5][11] , \u_div/SumTmp[5][12] , \u_div/SumTmp[5][13] ,
         \u_div/SumTmp[5][14] , \u_div/SumTmp[6][0] , \u_div/SumTmp[6][1] ,
         \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] , \u_div/SumTmp[6][4] ,
         \u_div/SumTmp[6][5] , \u_div/SumTmp[6][6] , \u_div/SumTmp[6][7] ,
         \u_div/SumTmp[6][8] , \u_div/SumTmp[6][9] , \u_div/SumTmp[6][10] ,
         \u_div/SumTmp[6][11] , \u_div/SumTmp[6][12] , \u_div/SumTmp[6][13] ,
         \u_div/SumTmp[7][0] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[7][5] ,
         \u_div/SumTmp[7][6] , \u_div/SumTmp[7][7] , \u_div/SumTmp[7][8] ,
         \u_div/SumTmp[7][9] , \u_div/SumTmp[7][10] , \u_div/SumTmp[7][11] ,
         \u_div/SumTmp[7][12] , \u_div/SumTmp[8][0] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[8][5] , \u_div/SumTmp[8][6] , \u_div/SumTmp[8][7] ,
         \u_div/SumTmp[8][8] , \u_div/SumTmp[8][9] , \u_div/SumTmp[8][10] ,
         \u_div/SumTmp[8][11] , \u_div/SumTmp[9][0] , \u_div/SumTmp[9][1] ,
         \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] , \u_div/SumTmp[9][4] ,
         \u_div/SumTmp[9][5] , \u_div/SumTmp[9][6] , \u_div/SumTmp[9][7] ,
         \u_div/SumTmp[9][8] , \u_div/SumTmp[9][9] , \u_div/SumTmp[9][10] ,
         \u_div/SumTmp[10][0] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[10][5] ,
         \u_div/SumTmp[10][6] , \u_div/SumTmp[10][7] , \u_div/SumTmp[10][8] ,
         \u_div/SumTmp[10][9] , \u_div/SumTmp[11][0] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] ,
         \u_div/SumTmp[11][5] , \u_div/SumTmp[11][6] , \u_div/SumTmp[11][7] ,
         \u_div/SumTmp[11][8] , \u_div/SumTmp[12][0] , \u_div/SumTmp[12][1] ,
         \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] , \u_div/SumTmp[12][4] ,
         \u_div/SumTmp[12][5] , \u_div/SumTmp[12][6] , \u_div/SumTmp[12][7] ,
         \u_div/SumTmp[13][0] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[13][4] , \u_div/SumTmp[13][5] ,
         \u_div/SumTmp[13][6] , \u_div/SumTmp[14][0] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] , \u_div/SumTmp[14][4] ,
         \u_div/SumTmp[14][5] , \u_div/SumTmp[15][0] , \u_div/SumTmp[15][1] ,
         \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] , \u_div/SumTmp[15][4] ,
         \u_div/SumTmp[16][0] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/SumTmp[17][0] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[18][0] , \u_div/SumTmp[18][1] ,
         \u_div/SumTmp[19][0] , \u_div/CryTmp[0][1] , \u_div/CryTmp[0][2] ,
         \u_div/CryTmp[0][3] , \u_div/CryTmp[0][4] , \u_div/CryTmp[0][5] ,
         \u_div/CryTmp[0][6] , \u_div/CryTmp[0][7] , \u_div/CryTmp[0][8] ,
         \u_div/CryTmp[0][9] , \u_div/CryTmp[0][10] , \u_div/CryTmp[0][11] ,
         \u_div/CryTmp[0][12] , \u_div/CryTmp[0][13] , \u_div/CryTmp[0][14] ,
         \u_div/CryTmp[0][15] , \u_div/CryTmp[0][16] , \u_div/CryTmp[0][17] ,
         \u_div/CryTmp[0][18] , \u_div/CryTmp[0][19] , \u_div/CryTmp[1][1] ,
         \u_div/CryTmp[1][2] , \u_div/CryTmp[1][3] , \u_div/CryTmp[1][4] ,
         \u_div/CryTmp[1][5] , \u_div/CryTmp[1][6] , \u_div/CryTmp[1][7] ,
         \u_div/CryTmp[1][8] , \u_div/CryTmp[1][9] , \u_div/CryTmp[1][10] ,
         \u_div/CryTmp[1][11] , \u_div/CryTmp[1][12] , \u_div/CryTmp[1][13] ,
         \u_div/CryTmp[1][14] , \u_div/CryTmp[1][15] , \u_div/CryTmp[1][16] ,
         \u_div/CryTmp[1][17] , \u_div/CryTmp[1][18] , \u_div/CryTmp[1][19] ,
         \u_div/CryTmp[2][1] , \u_div/CryTmp[2][2] , \u_div/CryTmp[2][3] ,
         \u_div/CryTmp[2][4] , \u_div/CryTmp[2][5] , \u_div/CryTmp[2][6] ,
         \u_div/CryTmp[2][7] , \u_div/CryTmp[2][8] , \u_div/CryTmp[2][9] ,
         \u_div/CryTmp[2][10] , \u_div/CryTmp[2][11] , \u_div/CryTmp[2][12] ,
         \u_div/CryTmp[2][13] , \u_div/CryTmp[2][14] , \u_div/CryTmp[2][15] ,
         \u_div/CryTmp[2][16] , \u_div/CryTmp[2][17] , \u_div/CryTmp[2][18] ,
         \u_div/CryTmp[3][1] , \u_div/CryTmp[3][2] , \u_div/CryTmp[3][3] ,
         \u_div/CryTmp[3][4] , \u_div/CryTmp[3][5] , \u_div/CryTmp[3][6] ,
         \u_div/CryTmp[3][7] , \u_div/CryTmp[3][8] , \u_div/CryTmp[3][9] ,
         \u_div/CryTmp[3][10] , \u_div/CryTmp[3][11] , \u_div/CryTmp[3][12] ,
         \u_div/CryTmp[3][13] , \u_div/CryTmp[3][14] , \u_div/CryTmp[3][15] ,
         \u_div/CryTmp[3][16] , \u_div/CryTmp[3][17] , \u_div/CryTmp[4][1] ,
         \u_div/CryTmp[4][2] , \u_div/CryTmp[4][3] , \u_div/CryTmp[4][4] ,
         \u_div/CryTmp[4][5] , \u_div/CryTmp[4][6] , \u_div/CryTmp[4][7] ,
         \u_div/CryTmp[4][8] , \u_div/CryTmp[4][9] , \u_div/CryTmp[4][10] ,
         \u_div/CryTmp[4][11] , \u_div/CryTmp[4][12] , \u_div/CryTmp[4][13] ,
         \u_div/CryTmp[4][14] , \u_div/CryTmp[4][15] , \u_div/CryTmp[4][16] ,
         \u_div/CryTmp[5][1] , \u_div/CryTmp[5][2] , \u_div/CryTmp[5][3] ,
         \u_div/CryTmp[5][4] , \u_div/CryTmp[5][5] , \u_div/CryTmp[5][6] ,
         \u_div/CryTmp[5][7] , \u_div/CryTmp[5][8] , \u_div/CryTmp[5][9] ,
         \u_div/CryTmp[5][10] , \u_div/CryTmp[5][11] , \u_div/CryTmp[5][12] ,
         \u_div/CryTmp[5][13] , \u_div/CryTmp[5][14] , \u_div/CryTmp[5][15] ,
         \u_div/CryTmp[6][1] , \u_div/CryTmp[6][2] , \u_div/CryTmp[6][3] ,
         \u_div/CryTmp[6][4] , \u_div/CryTmp[6][5] , \u_div/CryTmp[6][6] ,
         \u_div/CryTmp[6][7] , \u_div/CryTmp[6][8] , \u_div/CryTmp[6][9] ,
         \u_div/CryTmp[6][10] , \u_div/CryTmp[6][11] , \u_div/CryTmp[6][12] ,
         \u_div/CryTmp[6][13] , \u_div/CryTmp[6][14] , \u_div/CryTmp[7][1] ,
         \u_div/CryTmp[7][2] , \u_div/CryTmp[7][3] , \u_div/CryTmp[7][4] ,
         \u_div/CryTmp[7][5] , \u_div/CryTmp[7][6] , \u_div/CryTmp[7][7] ,
         \u_div/CryTmp[7][8] , \u_div/CryTmp[7][9] , \u_div/CryTmp[7][10] ,
         \u_div/CryTmp[7][11] , \u_div/CryTmp[7][12] , \u_div/CryTmp[7][13] ,
         \u_div/CryTmp[8][1] , \u_div/CryTmp[8][2] , \u_div/CryTmp[8][3] ,
         \u_div/CryTmp[8][4] , \u_div/CryTmp[8][5] , \u_div/CryTmp[8][6] ,
         \u_div/CryTmp[8][7] , \u_div/CryTmp[8][8] , \u_div/CryTmp[8][9] ,
         \u_div/CryTmp[8][10] , \u_div/CryTmp[8][11] , \u_div/CryTmp[8][12] ,
         \u_div/CryTmp[9][1] , \u_div/CryTmp[9][2] , \u_div/CryTmp[9][3] ,
         \u_div/CryTmp[9][4] , \u_div/CryTmp[9][5] , \u_div/CryTmp[9][6] ,
         \u_div/CryTmp[9][7] , \u_div/CryTmp[9][8] , \u_div/CryTmp[9][9] ,
         \u_div/CryTmp[9][10] , \u_div/CryTmp[9][11] , \u_div/CryTmp[10][1] ,
         \u_div/CryTmp[10][2] , \u_div/CryTmp[10][3] , \u_div/CryTmp[10][4] ,
         \u_div/CryTmp[10][5] , \u_div/CryTmp[10][6] , \u_div/CryTmp[10][7] ,
         \u_div/CryTmp[10][8] , \u_div/CryTmp[10][9] , \u_div/CryTmp[10][10] ,
         \u_div/CryTmp[11][1] , \u_div/CryTmp[11][2] , \u_div/CryTmp[11][3] ,
         \u_div/CryTmp[11][4] , \u_div/CryTmp[11][5] , \u_div/CryTmp[11][6] ,
         \u_div/CryTmp[11][7] , \u_div/CryTmp[11][8] , \u_div/CryTmp[11][9] ,
         \u_div/CryTmp[12][1] , \u_div/CryTmp[12][2] , \u_div/CryTmp[12][3] ,
         \u_div/CryTmp[12][4] , \u_div/CryTmp[12][5] , \u_div/CryTmp[12][6] ,
         \u_div/CryTmp[12][7] , \u_div/CryTmp[12][8] , \u_div/CryTmp[13][1] ,
         \u_div/CryTmp[13][2] , \u_div/CryTmp[13][3] , \u_div/CryTmp[13][4] ,
         \u_div/CryTmp[13][5] , \u_div/CryTmp[13][6] , \u_div/CryTmp[13][7] ,
         \u_div/CryTmp[14][1] , \u_div/CryTmp[14][2] , \u_div/CryTmp[14][3] ,
         \u_div/CryTmp[14][4] , \u_div/CryTmp[14][5] , \u_div/CryTmp[14][6] ,
         \u_div/CryTmp[15][1] , \u_div/CryTmp[15][2] , \u_div/CryTmp[15][3] ,
         \u_div/CryTmp[15][4] , \u_div/CryTmp[15][5] , \u_div/CryTmp[16][1] ,
         \u_div/CryTmp[16][2] , \u_div/CryTmp[16][3] , \u_div/CryTmp[16][4] ,
         \u_div/CryTmp[17][1] , \u_div/CryTmp[17][2] , \u_div/CryTmp[17][3] ,
         \u_div/CryTmp[18][1] , \u_div/CryTmp[18][2] , \u_div/CryTmp[19][1] ,
         \u_div/PartRem[1][1] , \u_div/PartRem[1][2] , \u_div/PartRem[1][3] ,
         \u_div/PartRem[1][4] , \u_div/PartRem[1][5] , \u_div/PartRem[1][6] ,
         \u_div/PartRem[1][7] , \u_div/PartRem[1][8] , \u_div/PartRem[1][9] ,
         \u_div/PartRem[1][10] , \u_div/PartRem[1][11] ,
         \u_div/PartRem[1][12] , \u_div/PartRem[1][13] ,
         \u_div/PartRem[1][14] , \u_div/PartRem[1][15] ,
         \u_div/PartRem[1][16] , \u_div/PartRem[1][17] ,
         \u_div/PartRem[1][18] , \u_div/PartRem[1][19] , \u_div/PartRem[2][1] ,
         \u_div/PartRem[2][2] , \u_div/PartRem[2][3] , \u_div/PartRem[2][4] ,
         \u_div/PartRem[2][5] , \u_div/PartRem[2][6] , \u_div/PartRem[2][7] ,
         \u_div/PartRem[2][8] , \u_div/PartRem[2][9] , \u_div/PartRem[2][10] ,
         \u_div/PartRem[2][11] , \u_div/PartRem[2][12] ,
         \u_div/PartRem[2][13] , \u_div/PartRem[2][14] ,
         \u_div/PartRem[2][15] , \u_div/PartRem[2][16] ,
         \u_div/PartRem[2][17] , \u_div/PartRem[2][18] , n1, n2, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224;
  wire   [19:0] \u_div/BInv ;

  ADDFX2 \u_div/u_fa_PartRem_0_2_1  ( .A(n7), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[2][1] ), .CO(\u_div/CryTmp[2][2] ), .S(
        \u_div/SumTmp[2][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_1  ( .A(n10), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[3][1] ), .CO(\u_div/CryTmp[3][2] ), .S(
        \u_div/SumTmp[3][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_1  ( .A(n9), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[4][1] ), .CO(\u_div/CryTmp[4][2] ), .S(
        \u_div/SumTmp[4][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_1  ( .A(n15), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[5][1] ), .CO(\u_div/CryTmp[5][2] ), .S(
        \u_div/SumTmp[5][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_1  ( .A(n16), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[6][1] ), .CO(\u_div/CryTmp[6][2] ), .S(
        \u_div/SumTmp[6][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_1  ( .A(n8), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[7][1] ), .CO(\u_div/CryTmp[7][2] ), .S(
        \u_div/SumTmp[7][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_1  ( .A(n13), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[8][1] ), .CO(\u_div/CryTmp[8][2] ), .S(
        \u_div/SumTmp[8][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_1  ( .A(n11), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[9][1] ), .CO(\u_div/CryTmp[9][2] ), .S(
        \u_div/SumTmp[9][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_1  ( .A(n18), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[10][1] ), .CO(\u_div/CryTmp[10][2] ), .S(
        \u_div/SumTmp[10][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_1  ( .A(n17), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[11][2] ), .S(
        \u_div/SumTmp[11][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_1  ( .A(n12), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[12][1] ), .CO(\u_div/CryTmp[12][2] ), .S(
        \u_div/SumTmp[12][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_1  ( .A(n21), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[13][1] ), .CO(\u_div/CryTmp[13][2] ), .S(
        \u_div/SumTmp[13][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_1  ( .A(n23), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[14][1] ), .CO(\u_div/CryTmp[14][2] ), .S(
        \u_div/SumTmp[14][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_1  ( .A(n19), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[15][1] ), .CO(\u_div/CryTmp[15][2] ), .S(
        \u_div/SumTmp[15][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_1  ( .A(n22), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[16][1] ), .CO(\u_div/CryTmp[16][2] ), .S(
        \u_div/SumTmp[16][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_1  ( .A(n20), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[17][1] ), .CO(\u_div/CryTmp[17][2] ), .S(
        \u_div/SumTmp[17][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_18_1  ( .A(n14), .B(\u_div/BInv [1]), .CI(
        \u_div/CryTmp[18][1] ), .CO(\u_div/CryTmp[18][2] ), .S(
        \u_div/SumTmp[18][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        \u_div/BInv [1]), .CI(\u_div/CryTmp[1][1] ), .CO(\u_div/CryTmp[1][2] ), 
        .S(\u_div/SumTmp[1][1] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_19  ( .A(\u_div/PartRem[1][19] ), .B(
        \u_div/BInv [19]), .CI(\u_div/CryTmp[0][19] ), .CO(quotient[0]) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_17  ( .A(\u_div/PartRem[1][17] ), .B(
        \u_div/BInv [17]), .CI(\u_div/CryTmp[0][17] ), .CO(
        \u_div/CryTmp[0][18] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_18  ( .A(\u_div/PartRem[1][18] ), .B(
        \u_div/BInv [18]), .CI(\u_div/CryTmp[0][18] ), .CO(
        \u_div/CryTmp[0][19] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_17  ( .A(\u_div/PartRem[2][17] ), .B(
        \u_div/BInv [17]), .CI(\u_div/CryTmp[1][17] ), .CO(
        \u_div/CryTmp[1][18] ), .S(\u_div/SumTmp[1][17] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_16  ( .A(\u_div/PartRem[2][16] ), .B(
        \u_div/BInv [16]), .CI(\u_div/CryTmp[1][16] ), .CO(
        \u_div/CryTmp[1][17] ), .S(\u_div/SumTmp[1][16] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_16  ( .A(n142), .B(\u_div/BInv [16]), .CI(
        \u_div/CryTmp[2][16] ), .CO(\u_div/CryTmp[2][17] ), .S(
        \u_div/SumTmp[2][16] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_15  ( .A(\u_div/PartRem[1][15] ), .B(
        \u_div/BInv [15]), .CI(\u_div/CryTmp[0][15] ), .CO(
        \u_div/CryTmp[0][16] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_16  ( .A(\u_div/PartRem[1][16] ), .B(
        \u_div/BInv [16]), .CI(\u_div/CryTmp[0][16] ), .CO(
        \u_div/CryTmp[0][17] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_15  ( .A(\u_div/PartRem[2][15] ), .B(
        \u_div/BInv [15]), .CI(\u_div/CryTmp[1][15] ), .CO(
        \u_div/CryTmp[1][16] ), .S(\u_div/SumTmp[1][15] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_15  ( .A(n141), .B(\u_div/BInv [15]), .CI(
        \u_div/CryTmp[2][15] ), .CO(\u_div/CryTmp[2][16] ), .S(
        \u_div/SumTmp[2][15] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_15  ( .A(n138), .B(\u_div/BInv [15]), .CI(
        \u_div/CryTmp[3][15] ), .CO(\u_div/CryTmp[3][16] ), .S(
        \u_div/SumTmp[3][15] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_14  ( .A(\u_div/PartRem[2][14] ), .B(
        \u_div/BInv [14]), .CI(\u_div/CryTmp[1][14] ), .CO(
        \u_div/CryTmp[1][15] ), .S(\u_div/SumTmp[1][14] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_14  ( .A(n137), .B(\u_div/BInv [14]), .CI(
        \u_div/CryTmp[2][14] ), .CO(\u_div/CryTmp[2][15] ), .S(
        \u_div/SumTmp[2][14] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_14  ( .A(n126), .B(\u_div/BInv [14]), .CI(
        \u_div/CryTmp[3][14] ), .CO(\u_div/CryTmp[3][15] ), .S(
        \u_div/SumTmp[3][14] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_14  ( .A(n129), .B(\u_div/BInv [14]), .CI(
        \u_div/CryTmp[4][14] ), .CO(\u_div/CryTmp[4][15] ), .S(
        \u_div/SumTmp[4][14] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_13  ( .A(\u_div/PartRem[1][13] ), .B(
        \u_div/BInv [13]), .CI(\u_div/CryTmp[0][13] ), .CO(
        \u_div/CryTmp[0][14] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_14  ( .A(\u_div/PartRem[1][14] ), .B(
        \u_div/BInv [14]), .CI(\u_div/CryTmp[0][14] ), .CO(
        \u_div/CryTmp[0][15] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_13  ( .A(\u_div/PartRem[2][13] ), .B(
        \u_div/BInv [13]), .CI(\u_div/CryTmp[1][13] ), .CO(
        \u_div/CryTmp[1][14] ), .S(\u_div/SumTmp[1][13] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_13  ( .A(n136), .B(\u_div/BInv [13]), .CI(
        \u_div/CryTmp[2][13] ), .CO(\u_div/CryTmp[2][14] ), .S(
        \u_div/SumTmp[2][13] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_13  ( .A(n125), .B(\u_div/BInv [13]), .CI(
        \u_div/CryTmp[3][13] ), .CO(\u_div/CryTmp[3][14] ), .S(
        \u_div/SumTmp[3][13] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_13  ( .A(n128), .B(\u_div/BInv [13]), .CI(
        \u_div/CryTmp[4][13] ), .CO(\u_div/CryTmp[4][14] ), .S(
        \u_div/SumTmp[4][13] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_13  ( .A(n131), .B(\u_div/BInv [13]), .CI(
        \u_div/CryTmp[5][13] ), .CO(\u_div/CryTmp[5][14] ), .S(
        \u_div/SumTmp[5][13] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_11  ( .A(\u_div/PartRem[1][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[0][11] ), .CO(
        \u_div/CryTmp[0][12] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_12  ( .A(\u_div/PartRem[1][12] ), .B(
        \u_div/BInv [12]), .CI(\u_div/CryTmp[0][12] ), .CO(
        \u_div/CryTmp[0][13] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_12  ( .A(\u_div/PartRem[2][12] ), .B(
        \u_div/BInv [12]), .CI(\u_div/CryTmp[1][12] ), .CO(
        \u_div/CryTmp[1][13] ), .S(\u_div/SumTmp[1][12] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_12  ( .A(n135), .B(\u_div/BInv [12]), .CI(
        \u_div/CryTmp[2][12] ), .CO(\u_div/CryTmp[2][13] ), .S(
        \u_div/SumTmp[2][12] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_12  ( .A(n124), .B(\u_div/BInv [12]), .CI(
        \u_div/CryTmp[3][12] ), .CO(\u_div/CryTmp[3][13] ), .S(
        \u_div/SumTmp[3][12] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_12  ( .A(n127), .B(\u_div/BInv [12]), .CI(
        \u_div/CryTmp[4][12] ), .CO(\u_div/CryTmp[4][13] ), .S(
        \u_div/SumTmp[4][12] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_12  ( .A(n130), .B(\u_div/BInv [12]), .CI(
        \u_div/CryTmp[5][12] ), .CO(\u_div/CryTmp[5][13] ), .S(
        \u_div/SumTmp[5][12] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_12  ( .A(n133), .B(\u_div/BInv [12]), .CI(
        \u_div/CryTmp[6][12] ), .CO(\u_div/CryTmp[6][13] ), .S(
        \u_div/SumTmp[6][12] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_11  ( .A(\u_div/PartRem[2][11] ), .B(
        \u_div/BInv [11]), .CI(\u_div/CryTmp[1][11] ), .CO(
        \u_div/CryTmp[1][12] ), .S(\u_div/SumTmp[1][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_11  ( .A(n122), .B(\u_div/BInv [11]), .CI(
        \u_div/CryTmp[2][11] ), .CO(\u_div/CryTmp[2][12] ), .S(
        \u_div/SumTmp[2][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_11  ( .A(n106), .B(\u_div/BInv [11]), .CI(
        \u_div/CryTmp[3][11] ), .CO(\u_div/CryTmp[3][12] ), .S(
        \u_div/SumTmp[3][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_11  ( .A(n109), .B(\u_div/BInv [11]), .CI(
        \u_div/CryTmp[4][11] ), .CO(\u_div/CryTmp[4][12] ), .S(
        \u_div/SumTmp[4][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_11  ( .A(n112), .B(\u_div/BInv [11]), .CI(
        \u_div/CryTmp[5][11] ), .CO(\u_div/CryTmp[5][12] ), .S(
        \u_div/SumTmp[5][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_11  ( .A(n115), .B(\u_div/BInv [11]), .CI(
        \u_div/CryTmp[6][11] ), .CO(\u_div/CryTmp[6][12] ), .S(
        \u_div/SumTmp[6][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_11  ( .A(n101), .B(\u_div/BInv [11]), .CI(
        \u_div/CryTmp[7][11] ), .CO(\u_div/CryTmp[7][12] ), .S(
        \u_div/SumTmp[7][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_9  ( .A(\u_div/PartRem[1][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[0][9] ), .CO(\u_div/CryTmp[0][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_10  ( .A(\u_div/PartRem[1][10] ), .B(
        \u_div/BInv [10]), .CI(\u_div/CryTmp[0][10] ), .CO(
        \u_div/CryTmp[0][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_10  ( .A(\u_div/PartRem[2][10] ), .B(
        \u_div/BInv [10]), .CI(\u_div/CryTmp[1][10] ), .CO(
        \u_div/CryTmp[1][11] ), .S(\u_div/SumTmp[1][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_10  ( .A(n121), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[2][10] ), .CO(\u_div/CryTmp[2][11] ), .S(
        \u_div/SumTmp[2][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_10  ( .A(n105), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[3][10] ), .CO(\u_div/CryTmp[3][11] ), .S(
        \u_div/SumTmp[3][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_10  ( .A(n108), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[4][10] ), .CO(\u_div/CryTmp[4][11] ), .S(
        \u_div/SumTmp[4][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_10  ( .A(n111), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[5][10] ), .CO(\u_div/CryTmp[5][11] ), .S(
        \u_div/SumTmp[5][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_10  ( .A(n114), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[6][10] ), .CO(\u_div/CryTmp[6][11] ), .S(
        \u_div/SumTmp[6][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_10  ( .A(n100), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[7][10] ), .CO(\u_div/CryTmp[7][11] ), .S(
        \u_div/SumTmp[7][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_10  ( .A(n117), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[8][10] ), .CO(\u_div/CryTmp[8][11] ), .S(
        \u_div/SumTmp[8][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_9  ( .A(\u_div/PartRem[2][9] ), .B(
        \u_div/BInv [9]), .CI(\u_div/CryTmp[1][9] ), .CO(\u_div/CryTmp[1][10] ), .S(\u_div/SumTmp[1][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_9  ( .A(n120), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[2][9] ), .CO(\u_div/CryTmp[2][10] ), .S(
        \u_div/SumTmp[2][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_9  ( .A(n104), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[3][9] ), .CO(\u_div/CryTmp[3][10] ), .S(
        \u_div/SumTmp[3][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_9  ( .A(n107), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[4][9] ), .CO(\u_div/CryTmp[4][10] ), .S(
        \u_div/SumTmp[4][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_9  ( .A(n110), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[5][9] ), .CO(\u_div/CryTmp[5][10] ), .S(
        \u_div/SumTmp[5][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_9  ( .A(n113), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[6][9] ), .CO(\u_div/CryTmp[6][10] ), .S(
        \u_div/SumTmp[6][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_9  ( .A(n99), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[7][9] ), .CO(\u_div/CryTmp[7][10] ), .S(
        \u_div/SumTmp[7][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_9  ( .A(n116), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[8][9] ), .CO(\u_div/CryTmp[8][10] ), .S(
        \u_div/SumTmp[8][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_9  ( .A(n102), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[9][9] ), .CO(\u_div/CryTmp[9][10] ), .S(
        \u_div/SumTmp[9][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_7  ( .A(\u_div/PartRem[1][7] ), .B(
        \u_div/BInv [7]), .CI(\u_div/CryTmp[0][7] ), .CO(\u_div/CryTmp[0][8] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_8  ( .A(\u_div/PartRem[1][8] ), .B(
        \u_div/BInv [8]), .CI(\u_div/CryTmp[0][8] ), .CO(\u_div/CryTmp[0][9] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_8  ( .A(\u_div/PartRem[2][8] ), .B(
        \u_div/BInv [8]), .CI(\u_div/CryTmp[1][8] ), .CO(\u_div/CryTmp[1][9] ), 
        .S(\u_div/SumTmp[1][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_8  ( .A(n98), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[2][8] ), .CO(\u_div/CryTmp[2][9] ), .S(
        \u_div/SumTmp[2][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_8  ( .A(n83), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[3][8] ), .CO(\u_div/CryTmp[3][9] ), .S(
        \u_div/SumTmp[3][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_8  ( .A(n85), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[4][8] ), .CO(\u_div/CryTmp[4][9] ), .S(
        \u_div/SumTmp[4][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_8  ( .A(n87), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[5][8] ), .CO(\u_div/CryTmp[5][9] ), .S(
        \u_div/SumTmp[5][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_8  ( .A(n89), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[6][8] ), .CO(\u_div/CryTmp[6][9] ), .S(
        \u_div/SumTmp[6][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_8  ( .A(n79), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[7][8] ), .CO(\u_div/CryTmp[7][9] ), .S(
        \u_div/SumTmp[7][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_8  ( .A(n91), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[8][8] ), .CO(\u_div/CryTmp[8][9] ), .S(
        \u_div/SumTmp[8][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_8  ( .A(n81), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[9][8] ), .CO(\u_div/CryTmp[9][9] ), .S(
        \u_div/SumTmp[9][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_8  ( .A(n93), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[10][8] ), .CO(\u_div/CryTmp[10][9] ), .S(
        \u_div/SumTmp[10][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_7  ( .A(\u_div/PartRem[2][7] ), .B(
        \u_div/BInv [7]), .CI(\u_div/CryTmp[1][7] ), .CO(\u_div/CryTmp[1][8] ), 
        .S(\u_div/SumTmp[1][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_7  ( .A(n97), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[2][7] ), .CO(\u_div/CryTmp[2][8] ), .S(
        \u_div/SumTmp[2][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_7  ( .A(n82), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[3][7] ), .CO(\u_div/CryTmp[3][8] ), .S(
        \u_div/SumTmp[3][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_7  ( .A(n84), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[4][7] ), .CO(\u_div/CryTmp[4][8] ), .S(
        \u_div/SumTmp[4][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_7  ( .A(n86), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[5][7] ), .CO(\u_div/CryTmp[5][8] ), .S(
        \u_div/SumTmp[5][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_7  ( .A(n88), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[6][7] ), .CO(\u_div/CryTmp[6][8] ), .S(
        \u_div/SumTmp[6][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_7  ( .A(n78), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[7][7] ), .CO(\u_div/CryTmp[7][8] ), .S(
        \u_div/SumTmp[7][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_7  ( .A(n90), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[8][7] ), .CO(\u_div/CryTmp[8][8] ), .S(
        \u_div/SumTmp[8][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_7  ( .A(n80), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[9][7] ), .CO(\u_div/CryTmp[9][8] ), .S(
        \u_div/SumTmp[9][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_7  ( .A(n92), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[10][7] ), .CO(\u_div/CryTmp[10][8] ), .S(
        \u_div/SumTmp[10][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_7  ( .A(n94), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[11][7] ), .CO(\u_div/CryTmp[11][8] ), .S(
        \u_div/SumTmp[11][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_5  ( .A(\u_div/PartRem[1][5] ), .B(
        \u_div/BInv [5]), .CI(\u_div/CryTmp[0][5] ), .CO(\u_div/CryTmp[0][6] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_6  ( .A(\u_div/PartRem[1][6] ), .B(
        \u_div/BInv [6]), .CI(\u_div/CryTmp[0][6] ), .CO(\u_div/CryTmp[0][7] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_6  ( .A(\u_div/PartRem[2][6] ), .B(
        \u_div/BInv [6]), .CI(\u_div/CryTmp[1][6] ), .CO(\u_div/CryTmp[1][7] ), 
        .S(\u_div/SumTmp[1][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_6  ( .A(n77), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[2][6] ), .CO(\u_div/CryTmp[2][7] ), .S(
        \u_div/SumTmp[2][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_6  ( .A(n47), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[3][6] ), .CO(\u_div/CryTmp[3][7] ), .S(
        \u_div/SumTmp[3][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_6  ( .A(n50), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[4][6] ), .CO(\u_div/CryTmp[4][7] ), .S(
        \u_div/SumTmp[4][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_6  ( .A(n53), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[5][6] ), .CO(\u_div/CryTmp[5][7] ), .S(
        \u_div/SumTmp[5][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_6  ( .A(n56), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[6][6] ), .CO(\u_div/CryTmp[6][7] ), .S(
        \u_div/SumTmp[6][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_6  ( .A(n41), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[7][6] ), .CO(\u_div/CryTmp[7][7] ), .S(
        \u_div/SumTmp[7][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_6  ( .A(n59), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[8][6] ), .CO(\u_div/CryTmp[8][7] ), .S(
        \u_div/SumTmp[8][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_6  ( .A(n44), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[9][6] ), .CO(\u_div/CryTmp[9][7] ), .S(
        \u_div/SumTmp[9][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_6  ( .A(n62), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[10][6] ), .CO(\u_div/CryTmp[10][7] ), .S(
        \u_div/SumTmp[10][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_6  ( .A(n65), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[11][6] ), .CO(\u_div/CryTmp[11][7] ), .S(
        \u_div/SumTmp[11][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_6  ( .A(n71), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[12][6] ), .CO(\u_div/CryTmp[12][7] ), .S(
        \u_div/SumTmp[12][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_5  ( .A(\u_div/PartRem[2][5] ), .B(
        \u_div/BInv [5]), .CI(\u_div/CryTmp[1][5] ), .CO(\u_div/CryTmp[1][6] ), 
        .S(\u_div/SumTmp[1][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_5  ( .A(n76), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[2][5] ), .CO(\u_div/CryTmp[2][6] ), .S(
        \u_div/SumTmp[2][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_5  ( .A(n46), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[3][5] ), .CO(\u_div/CryTmp[3][6] ), .S(
        \u_div/SumTmp[3][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_5  ( .A(n49), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[4][5] ), .CO(\u_div/CryTmp[4][6] ), .S(
        \u_div/SumTmp[4][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_5  ( .A(n52), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[5][5] ), .CO(\u_div/CryTmp[5][6] ), .S(
        \u_div/SumTmp[5][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_5  ( .A(n55), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[6][5] ), .CO(\u_div/CryTmp[6][6] ), .S(
        \u_div/SumTmp[6][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_5  ( .A(n40), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[7][5] ), .CO(\u_div/CryTmp[7][6] ), .S(
        \u_div/SumTmp[7][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_5  ( .A(n58), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[8][5] ), .CO(\u_div/CryTmp[8][6] ), .S(
        \u_div/SumTmp[8][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_5  ( .A(n43), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[9][5] ), .CO(\u_div/CryTmp[9][6] ), .S(
        \u_div/SumTmp[9][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_5  ( .A(n61), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[10][5] ), .CO(\u_div/CryTmp[10][6] ), .S(
        \u_div/SumTmp[10][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_5  ( .A(n64), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[11][5] ), .CO(\u_div/CryTmp[11][6] ), .S(
        \u_div/SumTmp[11][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_5  ( .A(n70), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[12][5] ), .CO(\u_div/CryTmp[12][6] ), .S(
        \u_div/SumTmp[12][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_5  ( .A(n67), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[13][5] ), .CO(\u_div/CryTmp[13][6] ), .S(
        \u_div/SumTmp[13][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/BInv [4]), .CI(\u_div/CryTmp[1][4] ), .CO(\u_div/CryTmp[1][5] ), 
        .S(\u_div/SumTmp[1][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_4  ( .A(n75), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[2][4] ), .CO(\u_div/CryTmp[2][5] ), .S(
        \u_div/SumTmp[2][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_4  ( .A(n45), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[3][4] ), .CO(\u_div/CryTmp[3][5] ), .S(
        \u_div/SumTmp[3][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_4  ( .A(n48), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[4][4] ), .CO(\u_div/CryTmp[4][5] ), .S(
        \u_div/SumTmp[4][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_4  ( .A(n51), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[5][4] ), .CO(\u_div/CryTmp[5][5] ), .S(
        \u_div/SumTmp[5][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_4  ( .A(n54), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[6][4] ), .CO(\u_div/CryTmp[6][5] ), .S(
        \u_div/SumTmp[6][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_4  ( .A(n39), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[7][4] ), .CO(\u_div/CryTmp[7][5] ), .S(
        \u_div/SumTmp[7][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_4  ( .A(n57), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[8][4] ), .CO(\u_div/CryTmp[8][5] ), .S(
        \u_div/SumTmp[8][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_4  ( .A(n42), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[9][4] ), .CO(\u_div/CryTmp[9][5] ), .S(
        \u_div/SumTmp[9][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_4  ( .A(n60), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[10][4] ), .CO(\u_div/CryTmp[10][5] ), .S(
        \u_div/SumTmp[10][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_4  ( .A(n63), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[11][4] ), .CO(\u_div/CryTmp[11][5] ), .S(
        \u_div/SumTmp[11][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_4  ( .A(n69), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[12][4] ), .CO(\u_div/CryTmp[12][5] ), .S(
        \u_div/SumTmp[12][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_4  ( .A(n66), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[13][4] ), .CO(\u_div/CryTmp[13][5] ), .S(
        \u_div/SumTmp[13][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_4  ( .A(n72), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[14][4] ), .CO(\u_div/CryTmp[14][5] ), .S(
        \u_div/SumTmp[14][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_3  ( .A(\u_div/PartRem[1][3] ), .B(
        \u_div/BInv [3]), .CI(\u_div/CryTmp[0][3] ), .CO(\u_div/CryTmp[0][4] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_4  ( .A(\u_div/PartRem[1][4] ), .B(
        \u_div/BInv [4]), .CI(\u_div/CryTmp[0][4] ), .CO(\u_div/CryTmp[0][5] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        \u_div/BInv [3]), .CI(\u_div/CryTmp[1][3] ), .CO(\u_div/CryTmp[1][4] ), 
        .S(\u_div/SumTmp[1][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_3  ( .A(n38), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[2][3] ), .CO(\u_div/CryTmp[2][4] ), .S(
        \u_div/SumTmp[2][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_3  ( .A(n27), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[3][3] ), .CO(\u_div/CryTmp[3][4] ), .S(
        \u_div/SumTmp[3][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_3  ( .A(n28), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[4][3] ), .CO(\u_div/CryTmp[4][4] ), .S(
        \u_div/SumTmp[4][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_3  ( .A(n29), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[5][3] ), .CO(\u_div/CryTmp[5][4] ), .S(
        \u_div/SumTmp[5][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_3  ( .A(n30), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[6][3] ), .CO(\u_div/CryTmp[6][4] ), .S(
        \u_div/SumTmp[6][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_3  ( .A(n24), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[7][3] ), .CO(\u_div/CryTmp[7][4] ), .S(
        \u_div/SumTmp[7][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_3  ( .A(n31), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[8][3] ), .CO(\u_div/CryTmp[8][4] ), .S(
        \u_div/SumTmp[8][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_3  ( .A(n25), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[9][3] ), .CO(\u_div/CryTmp[9][4] ), .S(
        \u_div/SumTmp[9][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_3  ( .A(n32), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[10][3] ), .CO(\u_div/CryTmp[10][4] ), .S(
        \u_div/SumTmp[10][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_3  ( .A(n33), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[11][3] ), .CO(\u_div/CryTmp[11][4] ), .S(
        \u_div/SumTmp[11][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_3  ( .A(n35), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[12][3] ), .CO(\u_div/CryTmp[12][4] ), .S(
        \u_div/SumTmp[12][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_3  ( .A(n34), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[13][3] ), .CO(\u_div/CryTmp[13][4] ), .S(
        \u_div/SumTmp[13][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_3  ( .A(n36), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[14][3] ), .CO(\u_div/CryTmp[14][4] ), .S(
        \u_div/SumTmp[14][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_3  ( .A(n37), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[15][3] ), .CO(\u_div/CryTmp[15][4] ), .S(
        \u_div/SumTmp[15][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/BInv [2]), .CI(\u_div/CryTmp[1][2] ), .CO(\u_div/CryTmp[1][3] ), 
        .S(\u_div/SumTmp[1][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_2  ( .A(n160), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[2][2] ), .CO(\u_div/CryTmp[2][3] ), .S(
        \u_div/SumTmp[2][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_2  ( .A(n148), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[3][2] ), .CO(\u_div/CryTmp[3][3] ), .S(
        \u_div/SumTmp[3][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_2  ( .A(n149), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[4][2] ), .CO(\u_div/CryTmp[4][3] ), .S(
        \u_div/SumTmp[4][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_2  ( .A(n150), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[5][2] ), .CO(\u_div/CryTmp[5][3] ), .S(
        \u_div/SumTmp[5][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_6_2  ( .A(n151), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[6][2] ), .CO(\u_div/CryTmp[6][3] ), .S(
        \u_div/SumTmp[6][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_2  ( .A(n145), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[7][2] ), .CO(\u_div/CryTmp[7][3] ), .S(
        \u_div/SumTmp[7][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_2  ( .A(n152), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[8][2] ), .CO(\u_div/CryTmp[8][3] ), .S(
        \u_div/SumTmp[8][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_2  ( .A(n146), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[9][2] ), .CO(\u_div/CryTmp[9][3] ), .S(
        \u_div/SumTmp[9][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_2  ( .A(n153), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[10][2] ), .CO(\u_div/CryTmp[10][3] ), .S(
        \u_div/SumTmp[10][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_2  ( .A(n154), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[11][2] ), .CO(\u_div/CryTmp[11][3] ), .S(
        \u_div/SumTmp[11][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_2  ( .A(n156), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[12][2] ), .CO(\u_div/CryTmp[12][3] ), .S(
        \u_div/SumTmp[12][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_2  ( .A(n155), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[13][2] ), .CO(\u_div/CryTmp[13][3] ), .S(
        \u_div/SumTmp[13][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_2  ( .A(n157), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[14][2] ), .CO(\u_div/CryTmp[14][3] ), .S(
        \u_div/SumTmp[14][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_2  ( .A(n158), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[15][2] ), .CO(\u_div/CryTmp[15][3] ), .S(
        \u_div/SumTmp[15][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_2  ( .A(n147), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[16][2] ), .CO(\u_div/CryTmp[16][3] ), .S(
        \u_div/SumTmp[16][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_0_1  ( .A(\u_div/PartRem[1][1] ), .B(
        \u_div/BInv [1]), .CI(\u_div/CryTmp[0][1] ), .CO(\u_div/CryTmp[0][2] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/BInv [2]), .CI(\u_div/CryTmp[0][2] ), .CO(\u_div/CryTmp[0][3] )
         );
  ADDFX2 \u_div/u_fa_PartRem_0_6_13  ( .A(n134), .B(\u_div/BInv [13]), .CI(
        \u_div/CryTmp[6][13] ), .CO(\u_div/CryTmp[6][14] ), .S(
        \u_div/SumTmp[6][13] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_9_10  ( .A(n103), .B(\u_div/BInv [10]), .CI(
        \u_div/CryTmp[9][10] ), .CO(\u_div/CryTmp[9][11] ), .S(
        \u_div/SumTmp[9][10] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_12_7  ( .A(n96), .B(\u_div/BInv [7]), .CI(
        \u_div/CryTmp[12][7] ), .CO(\u_div/CryTmp[12][8] ), .S(
        \u_div/SumTmp[12][7] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_15_4  ( .A(n74), .B(\u_div/BInv [4]), .CI(
        \u_div/CryTmp[15][4] ), .CO(\u_div/CryTmp[15][5] ), .S(
        \u_div/SumTmp[15][4] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_1_18  ( .A(\u_div/PartRem[2][18] ), .B(
        \u_div/BInv [18]), .CI(\u_div/CryTmp[1][18] ), .CO(
        \u_div/CryTmp[1][19] ), .S(\u_div/SumTmp[1][18] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_5_14  ( .A(n132), .B(\u_div/BInv [14]), .CI(
        \u_div/CryTmp[5][14] ), .CO(\u_div/CryTmp[5][15] ), .S(
        \u_div/SumTmp[5][14] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_8_11  ( .A(n118), .B(\u_div/BInv [11]), .CI(
        \u_div/CryTmp[8][11] ), .CO(\u_div/CryTmp[8][12] ), .S(
        \u_div/SumTmp[8][11] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_11_8  ( .A(n95), .B(\u_div/BInv [8]), .CI(
        \u_div/CryTmp[11][8] ), .CO(\u_div/CryTmp[11][9] ), .S(
        \u_div/SumTmp[11][8] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_4_15  ( .A(n140), .B(\u_div/BInv [15]), .CI(
        \u_div/CryTmp[4][15] ), .CO(\u_div/CryTmp[4][16] ), .S(
        \u_div/SumTmp[4][15] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_7_12  ( .A(n123), .B(\u_div/BInv [12]), .CI(
        \u_div/CryTmp[7][12] ), .CO(\u_div/CryTmp[7][13] ), .S(
        \u_div/SumTmp[7][12] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_10_9  ( .A(n119), .B(\u_div/BInv [9]), .CI(
        \u_div/CryTmp[10][9] ), .CO(\u_div/CryTmp[10][10] ), .S(
        \u_div/SumTmp[10][9] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_14_5  ( .A(n73), .B(\u_div/BInv [5]), .CI(
        \u_div/CryTmp[14][5] ), .CO(\u_div/CryTmp[14][6] ), .S(
        \u_div/SumTmp[14][5] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_13_6  ( .A(n68), .B(\u_div/BInv [6]), .CI(
        \u_div/CryTmp[13][6] ), .CO(\u_div/CryTmp[13][7] ), .S(
        \u_div/SumTmp[13][6] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_17_2  ( .A(n159), .B(\u_div/BInv [2]), .CI(
        \u_div/CryTmp[17][2] ), .CO(\u_div/CryTmp[17][3] ), .S(
        \u_div/SumTmp[17][2] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_16_3  ( .A(n26), .B(\u_div/BInv [3]), .CI(
        \u_div/CryTmp[16][3] ), .CO(\u_div/CryTmp[16][4] ), .S(
        \u_div/SumTmp[16][3] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_2_17  ( .A(n143), .B(\u_div/BInv [17]), .CI(
        \u_div/CryTmp[2][17] ), .CO(\u_div/CryTmp[2][18] ), .S(
        \u_div/SumTmp[2][17] ) );
  ADDFX2 \u_div/u_fa_PartRem_0_3_16  ( .A(n139), .B(\u_div/BInv [16]), .CI(
        \u_div/CryTmp[3][16] ), .CO(\u_div/CryTmp[3][17] ), .S(
        \u_div/SumTmp[3][16] ) );
  CLKINVX3 U1 ( .A(n203), .Y(quotient[6]) );
  INVX4 U2 ( .A(b[1]), .Y(\u_div/BInv [1]) );
  INVX4 U3 ( .A(b[3]), .Y(\u_div/BInv [3]) );
  INVX4 U4 ( .A(b[2]), .Y(\u_div/BInv [2]) );
  NOR2X2 U5 ( .A(n207), .B(n209), .Y(n1) );
  NOR3X2 U6 ( .A(b[17]), .B(n207), .C(n208), .Y(n2) );
  AND2X4 U7 ( .A(\u_div/CryTmp[4][16] ), .B(n206), .Y(quotient[4]) );
  AND2X4 U8 ( .A(\u_div/CryTmp[10][10] ), .B(n224), .Y(quotient[10]) );
  AND2X4 U9 ( .A(\u_div/CryTmp[7][13] ), .B(n202), .Y(quotient[7]) );
  AND2X2 U10 ( .A(n211), .B(n212), .Y(quotient[19]) );
  MX2X1 U11 ( .A(a[3]), .B(\u_div/SumTmp[3][0] ), .S0(quotient[3]), .Y(n7) );
  MX2X1 U12 ( .A(a[8]), .B(\u_div/SumTmp[8][0] ), .S0(quotient[8]), .Y(n8) );
  MX2X1 U13 ( .A(a[5]), .B(\u_div/SumTmp[5][0] ), .S0(quotient[5]), .Y(n9) );
  MX2X1 U14 ( .A(a[4]), .B(\u_div/SumTmp[4][0] ), .S0(quotient[4]), .Y(n10) );
  MX2X1 U15 ( .A(a[10]), .B(\u_div/SumTmp[10][0] ), .S0(quotient[10]), .Y(n11)
         );
  MX2X1 U16 ( .A(a[13]), .B(\u_div/SumTmp[13][0] ), .S0(quotient[13]), .Y(n12)
         );
  MX2X1 U17 ( .A(a[9]), .B(\u_div/SumTmp[9][0] ), .S0(quotient[9]), .Y(n13) );
  MX2X1 U18 ( .A(a[19]), .B(\u_div/SumTmp[19][0] ), .S0(quotient[19]), .Y(n14)
         );
  MX2X1 U19 ( .A(a[6]), .B(\u_div/SumTmp[6][0] ), .S0(quotient[6]), .Y(n15) );
  MX2X1 U20 ( .A(a[7]), .B(\u_div/SumTmp[7][0] ), .S0(quotient[7]), .Y(n16) );
  MX2X1 U21 ( .A(a[12]), .B(\u_div/SumTmp[12][0] ), .S0(quotient[12]), .Y(n17)
         );
  MX2X1 U22 ( .A(a[11]), .B(\u_div/SumTmp[11][0] ), .S0(quotient[11]), .Y(n18)
         );
  MX2X1 U23 ( .A(a[16]), .B(\u_div/SumTmp[16][0] ), .S0(quotient[16]), .Y(n19)
         );
  MX2X1 U24 ( .A(a[18]), .B(\u_div/SumTmp[18][0] ), .S0(quotient[18]), .Y(n20)
         );
  MX2X1 U25 ( .A(a[14]), .B(\u_div/SumTmp[14][0] ), .S0(quotient[14]), .Y(n21)
         );
  MX2X1 U26 ( .A(a[17]), .B(\u_div/SumTmp[17][0] ), .S0(quotient[17]), .Y(n22)
         );
  MX2X1 U27 ( .A(a[15]), .B(\u_div/SumTmp[15][0] ), .S0(quotient[15]), .Y(n23)
         );
  CLKINVX3 U28 ( .A(b[6]), .Y(\u_div/BInv [6]) );
  CLKINVX3 U29 ( .A(b[4]), .Y(\u_div/BInv [4]) );
  CLKINVX3 U30 ( .A(b[5]), .Y(\u_div/BInv [5]) );
  CLKINVX3 U31 ( .A(b[7]), .Y(\u_div/BInv [7]) );
  CLKINVX3 U32 ( .A(b[8]), .Y(\u_div/BInv [8]) );
  CLKINVX3 U33 ( .A(n201), .Y(quotient[8]) );
  NAND2BX1 U34 ( .AN(n200), .B(\u_div/CryTmp[8][12] ), .Y(n201) );
  CLKINVX3 U35 ( .A(n223), .Y(quotient[11]) );
  NAND2BX1 U36 ( .AN(n221), .B(\u_div/CryTmp[11][9] ), .Y(n223) );
  CLKINVX3 U37 ( .A(n219), .Y(quotient[14]) );
  NAND2BX1 U38 ( .AN(n217), .B(\u_div/CryTmp[14][6] ), .Y(n219) );
  CLKINVX3 U39 ( .A(n215), .Y(quotient[17]) );
  NAND2BX1 U40 ( .AN(n213), .B(\u_div/CryTmp[17][3] ), .Y(n215) );
  MXI2X1 U41 ( .A(n160), .B(\u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(n169)
         );
  MX2X1 U42 ( .A(n152), .B(\u_div/SumTmp[8][2] ), .S0(quotient[8]), .Y(n24) );
  MX2X1 U43 ( .A(n153), .B(\u_div/SumTmp[10][2] ), .S0(quotient[10]), .Y(n25)
         );
  MX2X1 U44 ( .A(n159), .B(\u_div/SumTmp[17][2] ), .S0(quotient[17]), .Y(n26)
         );
  MXI2X1 U45 ( .A(n170), .B(n187), .S0(quotient[1]), .Y(\u_div/PartRem[1][3] )
         );
  INVX1 U46 ( .A(\u_div/SumTmp[1][2] ), .Y(n187) );
  MX2X1 U47 ( .A(n149), .B(\u_div/SumTmp[4][2] ), .S0(quotient[4]), .Y(n27) );
  MX2X1 U48 ( .A(n150), .B(\u_div/SumTmp[5][2] ), .S0(quotient[5]), .Y(n28) );
  MX2X1 U49 ( .A(n151), .B(\u_div/SumTmp[6][2] ), .S0(quotient[6]), .Y(n29) );
  MX2X1 U50 ( .A(n145), .B(\u_div/SumTmp[7][2] ), .S0(quotient[7]), .Y(n30) );
  MX2X1 U51 ( .A(n146), .B(\u_div/SumTmp[9][2] ), .S0(quotient[9]), .Y(n31) );
  MX2X1 U52 ( .A(n154), .B(\u_div/SumTmp[11][2] ), .S0(quotient[11]), .Y(n32)
         );
  MX2X1 U53 ( .A(n156), .B(\u_div/SumTmp[12][2] ), .S0(quotient[12]), .Y(n33)
         );
  MX2X1 U54 ( .A(n157), .B(\u_div/SumTmp[14][2] ), .S0(quotient[14]), .Y(n34)
         );
  MX2X1 U55 ( .A(n155), .B(\u_div/SumTmp[13][2] ), .S0(quotient[13]), .Y(n35)
         );
  MX2X1 U56 ( .A(n158), .B(\u_div/SumTmp[15][2] ), .S0(quotient[15]), .Y(n36)
         );
  MX2X1 U57 ( .A(n147), .B(\u_div/SumTmp[16][2] ), .S0(quotient[16]), .Y(n37)
         );
  MX2X1 U58 ( .A(n148), .B(\u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(n38) );
  BUFX3 U59 ( .A(n1), .Y(quotient[2]) );
  NAND2BX1 U60 ( .AN(n204), .B(\u_div/CryTmp[5][15] ), .Y(n205) );
  MXI2X1 U61 ( .A(n38), .B(\u_div/SumTmp[2][3] ), .S0(quotient[2]), .Y(n168)
         );
  MXI2X1 U62 ( .A(n75), .B(\u_div/SumTmp[2][4] ), .S0(quotient[2]), .Y(n167)
         );
  MX2X1 U63 ( .A(n31), .B(\u_div/SumTmp[8][3] ), .S0(quotient[8]), .Y(n39) );
  MX2X1 U64 ( .A(n57), .B(\u_div/SumTmp[8][4] ), .S0(quotient[8]), .Y(n40) );
  MX2X1 U65 ( .A(n58), .B(\u_div/SumTmp[8][5] ), .S0(quotient[8]), .Y(n41) );
  MX2X1 U66 ( .A(n32), .B(\u_div/SumTmp[10][3] ), .S0(quotient[10]), .Y(n42)
         );
  MX2X1 U67 ( .A(n60), .B(\u_div/SumTmp[10][4] ), .S0(quotient[10]), .Y(n43)
         );
  MX2X1 U68 ( .A(n61), .B(\u_div/SumTmp[10][5] ), .S0(quotient[10]), .Y(n44)
         );
  MXI2X1 U69 ( .A(n168), .B(n185), .S0(quotient[1]), .Y(\u_div/PartRem[1][5] )
         );
  INVX1 U70 ( .A(\u_div/SumTmp[1][4] ), .Y(n185) );
  MX2X1 U71 ( .A(n28), .B(\u_div/SumTmp[4][3] ), .S0(quotient[4]), .Y(n45) );
  MX2X1 U72 ( .A(n48), .B(\u_div/SumTmp[4][4] ), .S0(quotient[4]), .Y(n46) );
  MX2X1 U73 ( .A(n49), .B(\u_div/SumTmp[4][5] ), .S0(quotient[4]), .Y(n47) );
  MX2X1 U74 ( .A(n29), .B(\u_div/SumTmp[5][3] ), .S0(quotient[5]), .Y(n48) );
  MX2X1 U75 ( .A(n51), .B(\u_div/SumTmp[5][4] ), .S0(quotient[5]), .Y(n49) );
  MX2X1 U76 ( .A(n52), .B(\u_div/SumTmp[5][5] ), .S0(quotient[5]), .Y(n50) );
  MX2X1 U77 ( .A(n30), .B(\u_div/SumTmp[6][3] ), .S0(quotient[6]), .Y(n51) );
  MX2X1 U78 ( .A(n54), .B(\u_div/SumTmp[6][4] ), .S0(quotient[6]), .Y(n52) );
  MX2X1 U79 ( .A(n55), .B(\u_div/SumTmp[6][5] ), .S0(quotient[6]), .Y(n53) );
  MX2X1 U80 ( .A(n24), .B(\u_div/SumTmp[7][3] ), .S0(quotient[7]), .Y(n54) );
  MX2X1 U81 ( .A(n39), .B(\u_div/SumTmp[7][4] ), .S0(quotient[7]), .Y(n55) );
  MX2X1 U82 ( .A(n40), .B(\u_div/SumTmp[7][5] ), .S0(quotient[7]), .Y(n56) );
  MX2X1 U83 ( .A(n25), .B(\u_div/SumTmp[9][3] ), .S0(quotient[9]), .Y(n57) );
  MX2X1 U84 ( .A(n42), .B(\u_div/SumTmp[9][4] ), .S0(quotient[9]), .Y(n58) );
  MX2X1 U85 ( .A(n43), .B(\u_div/SumTmp[9][5] ), .S0(quotient[9]), .Y(n59) );
  MX2X1 U86 ( .A(n33), .B(\u_div/SumTmp[11][3] ), .S0(quotient[11]), .Y(n60)
         );
  MX2X1 U87 ( .A(n63), .B(\u_div/SumTmp[11][4] ), .S0(quotient[11]), .Y(n61)
         );
  MX2X1 U88 ( .A(n64), .B(\u_div/SumTmp[11][5] ), .S0(quotient[11]), .Y(n62)
         );
  MX2X1 U89 ( .A(n35), .B(\u_div/SumTmp[12][3] ), .S0(quotient[12]), .Y(n63)
         );
  MX2X1 U90 ( .A(n69), .B(\u_div/SumTmp[12][4] ), .S0(quotient[12]), .Y(n64)
         );
  MX2X1 U91 ( .A(n70), .B(\u_div/SumTmp[12][5] ), .S0(quotient[12]), .Y(n65)
         );
  MX2X1 U92 ( .A(n36), .B(\u_div/SumTmp[14][3] ), .S0(quotient[14]), .Y(n66)
         );
  MX2X1 U93 ( .A(n72), .B(\u_div/SumTmp[14][4] ), .S0(quotient[14]), .Y(n67)
         );
  MX2X1 U94 ( .A(n73), .B(\u_div/SumTmp[14][5] ), .S0(quotient[14]), .Y(n68)
         );
  MX2X1 U95 ( .A(n34), .B(\u_div/SumTmp[13][3] ), .S0(quotient[13]), .Y(n69)
         );
  MX2X1 U96 ( .A(n66), .B(\u_div/SumTmp[13][4] ), .S0(quotient[13]), .Y(n70)
         );
  MX2X1 U97 ( .A(n67), .B(\u_div/SumTmp[13][5] ), .S0(quotient[13]), .Y(n71)
         );
  MX2X1 U98 ( .A(n37), .B(\u_div/SumTmp[15][3] ), .S0(quotient[15]), .Y(n72)
         );
  MX2X1 U99 ( .A(n74), .B(\u_div/SumTmp[15][4] ), .S0(quotient[15]), .Y(n73)
         );
  MX2X1 U100 ( .A(n26), .B(\u_div/SumTmp[16][3] ), .S0(quotient[16]), .Y(n74)
         );
  MX2X1 U101 ( .A(n27), .B(\u_div/SumTmp[3][3] ), .S0(quotient[3]), .Y(n75) );
  MX2X1 U102 ( .A(n45), .B(\u_div/SumTmp[3][4] ), .S0(quotient[3]), .Y(n76) );
  MX2X1 U103 ( .A(n46), .B(\u_div/SumTmp[3][5] ), .S0(quotient[3]), .Y(n77) );
  MXI2X1 U104 ( .A(n76), .B(\u_div/SumTmp[2][5] ), .S0(quotient[2]), .Y(n166)
         );
  MXI2X1 U105 ( .A(n97), .B(\u_div/SumTmp[2][7] ), .S0(quotient[2]), .Y(n164)
         );
  MXI2X1 U106 ( .A(n77), .B(\u_div/SumTmp[2][6] ), .S0(quotient[2]), .Y(n165)
         );
  MX2X1 U107 ( .A(n59), .B(\u_div/SumTmp[8][6] ), .S0(quotient[8]), .Y(n78) );
  MX2X1 U108 ( .A(n90), .B(\u_div/SumTmp[8][7] ), .S0(quotient[8]), .Y(n79) );
  MX2X1 U109 ( .A(n62), .B(\u_div/SumTmp[10][6] ), .S0(quotient[10]), .Y(n80)
         );
  MX2X1 U110 ( .A(n92), .B(\u_div/SumTmp[10][7] ), .S0(quotient[10]), .Y(n81)
         );
  MXI2X1 U111 ( .A(n166), .B(n183), .S0(quotient[1]), .Y(\u_div/PartRem[1][7] ) );
  INVX1 U112 ( .A(\u_div/SumTmp[1][6] ), .Y(n183) );
  MX2X1 U113 ( .A(n50), .B(\u_div/SumTmp[4][6] ), .S0(quotient[4]), .Y(n82) );
  MX2X1 U114 ( .A(n84), .B(\u_div/SumTmp[4][7] ), .S0(quotient[4]), .Y(n83) );
  MX2X1 U115 ( .A(n53), .B(\u_div/SumTmp[5][6] ), .S0(quotient[5]), .Y(n84) );
  MX2X1 U116 ( .A(n86), .B(\u_div/SumTmp[5][7] ), .S0(quotient[5]), .Y(n85) );
  MX2X1 U117 ( .A(n56), .B(\u_div/SumTmp[6][6] ), .S0(quotient[6]), .Y(n86) );
  MX2X1 U118 ( .A(n88), .B(\u_div/SumTmp[6][7] ), .S0(quotient[6]), .Y(n87) );
  MX2X1 U119 ( .A(n41), .B(\u_div/SumTmp[7][6] ), .S0(quotient[7]), .Y(n88) );
  MX2X1 U120 ( .A(n78), .B(\u_div/SumTmp[7][7] ), .S0(quotient[7]), .Y(n89) );
  MX2X1 U121 ( .A(n44), .B(\u_div/SumTmp[9][6] ), .S0(quotient[9]), .Y(n90) );
  MX2X1 U122 ( .A(n80), .B(\u_div/SumTmp[9][7] ), .S0(quotient[9]), .Y(n91) );
  MX2X1 U123 ( .A(n65), .B(\u_div/SumTmp[11][6] ), .S0(quotient[11]), .Y(n92)
         );
  MX2X1 U124 ( .A(n94), .B(\u_div/SumTmp[11][7] ), .S0(quotient[11]), .Y(n93)
         );
  MX2X1 U125 ( .A(n71), .B(\u_div/SumTmp[12][6] ), .S0(quotient[12]), .Y(n94)
         );
  MX2X1 U126 ( .A(n96), .B(\u_div/SumTmp[12][7] ), .S0(quotient[12]), .Y(n95)
         );
  MX2X1 U127 ( .A(n68), .B(\u_div/SumTmp[13][6] ), .S0(quotient[13]), .Y(n96)
         );
  MX2X1 U128 ( .A(n47), .B(\u_div/SumTmp[3][6] ), .S0(quotient[3]), .Y(n97) );
  MX2X1 U129 ( .A(n82), .B(\u_div/SumTmp[3][7] ), .S0(quotient[3]), .Y(n98) );
  MXI2X1 U130 ( .A(n120), .B(\u_div/SumTmp[2][9] ), .S0(quotient[2]), .Y(n180)
         );
  MXI2X1 U131 ( .A(n98), .B(\u_div/SumTmp[2][8] ), .S0(quotient[2]), .Y(n163)
         );
  MXI2X1 U132 ( .A(n121), .B(\u_div/SumTmp[2][10] ), .S0(n1), .Y(n179) );
  MX2X1 U133 ( .A(n91), .B(\u_div/SumTmp[8][8] ), .S0(quotient[8]), .Y(n99) );
  MX2X1 U134 ( .A(n116), .B(\u_div/SumTmp[8][9] ), .S0(quotient[8]), .Y(n100)
         );
  MX2X1 U135 ( .A(n117), .B(\u_div/SumTmp[8][10] ), .S0(quotient[8]), .Y(n101)
         );
  MX2X1 U136 ( .A(n93), .B(\u_div/SumTmp[10][8] ), .S0(quotient[10]), .Y(n102)
         );
  MX2X1 U137 ( .A(n119), .B(\u_div/SumTmp[10][9] ), .S0(quotient[10]), .Y(n103) );
  MXI2X1 U138 ( .A(n180), .B(n197), .S0(n162), .Y(\u_div/PartRem[1][11] ) );
  INVX1 U139 ( .A(\u_div/SumTmp[1][10] ), .Y(n197) );
  MXI2X1 U140 ( .A(n164), .B(n181), .S0(quotient[1]), .Y(\u_div/PartRem[1][9] ) );
  INVX1 U141 ( .A(\u_div/SumTmp[1][8] ), .Y(n181) );
  MX2X1 U142 ( .A(n85), .B(\u_div/SumTmp[4][8] ), .S0(quotient[4]), .Y(n104)
         );
  MX2X1 U143 ( .A(n107), .B(\u_div/SumTmp[4][9] ), .S0(quotient[4]), .Y(n105)
         );
  MX2X1 U144 ( .A(n108), .B(\u_div/SumTmp[4][10] ), .S0(quotient[4]), .Y(n106)
         );
  MX2X1 U145 ( .A(n87), .B(\u_div/SumTmp[5][8] ), .S0(quotient[5]), .Y(n107)
         );
  MX2X1 U146 ( .A(n110), .B(\u_div/SumTmp[5][9] ), .S0(quotient[5]), .Y(n108)
         );
  MX2X1 U147 ( .A(n111), .B(\u_div/SumTmp[5][10] ), .S0(quotient[5]), .Y(n109)
         );
  MX2X1 U148 ( .A(n89), .B(\u_div/SumTmp[6][8] ), .S0(quotient[6]), .Y(n110)
         );
  MX2X1 U149 ( .A(n113), .B(\u_div/SumTmp[6][9] ), .S0(quotient[6]), .Y(n111)
         );
  MX2X1 U150 ( .A(n114), .B(\u_div/SumTmp[6][10] ), .S0(quotient[6]), .Y(n112)
         );
  MX2X1 U151 ( .A(n79), .B(\u_div/SumTmp[7][8] ), .S0(quotient[7]), .Y(n113)
         );
  MX2X1 U152 ( .A(n99), .B(\u_div/SumTmp[7][9] ), .S0(quotient[7]), .Y(n114)
         );
  MX2X1 U153 ( .A(n100), .B(\u_div/SumTmp[7][10] ), .S0(quotient[7]), .Y(n115)
         );
  MX2X1 U154 ( .A(n81), .B(\u_div/SumTmp[9][8] ), .S0(quotient[9]), .Y(n116)
         );
  MX2X1 U155 ( .A(n102), .B(\u_div/SumTmp[9][9] ), .S0(quotient[9]), .Y(n117)
         );
  MX2X1 U156 ( .A(n103), .B(\u_div/SumTmp[9][10] ), .S0(quotient[9]), .Y(n118)
         );
  MX2X1 U157 ( .A(n95), .B(\u_div/SumTmp[11][8] ), .S0(quotient[11]), .Y(n119)
         );
  MX2X1 U158 ( .A(n83), .B(\u_div/SumTmp[3][8] ), .S0(quotient[3]), .Y(n120)
         );
  MX2X1 U159 ( .A(n104), .B(\u_div/SumTmp[3][9] ), .S0(n2), .Y(n121) );
  MX2X1 U160 ( .A(n105), .B(\u_div/SumTmp[3][10] ), .S0(n2), .Y(n122) );
  MXI2X1 U161 ( .A(n122), .B(\u_div/SumTmp[2][11] ), .S0(n1), .Y(n178) );
  MXI2X1 U162 ( .A(n136), .B(\u_div/SumTmp[2][13] ), .S0(n1), .Y(n176) );
  MXI2X1 U163 ( .A(n135), .B(\u_div/SumTmp[2][12] ), .S0(n1), .Y(n177) );
  MX2X1 U164 ( .A(n118), .B(\u_div/SumTmp[8][11] ), .S0(quotient[8]), .Y(n123)
         );
  MXI2X1 U165 ( .A(n178), .B(n195), .S0(n162), .Y(\u_div/PartRem[1][13] ) );
  INVX1 U166 ( .A(\u_div/SumTmp[1][12] ), .Y(n195) );
  MX2X1 U167 ( .A(n109), .B(\u_div/SumTmp[4][11] ), .S0(quotient[4]), .Y(n124)
         );
  MX2X1 U168 ( .A(n127), .B(\u_div/SumTmp[4][12] ), .S0(quotient[4]), .Y(n125)
         );
  MX2X1 U169 ( .A(n128), .B(\u_div/SumTmp[4][13] ), .S0(quotient[4]), .Y(n126)
         );
  MX2X1 U170 ( .A(n112), .B(\u_div/SumTmp[5][11] ), .S0(quotient[5]), .Y(n127)
         );
  MX2X1 U171 ( .A(n130), .B(\u_div/SumTmp[5][12] ), .S0(quotient[5]), .Y(n128)
         );
  MX2X1 U172 ( .A(n131), .B(\u_div/SumTmp[5][13] ), .S0(quotient[5]), .Y(n129)
         );
  MX2X1 U173 ( .A(n115), .B(\u_div/SumTmp[6][11] ), .S0(quotient[6]), .Y(n130)
         );
  MX2X1 U174 ( .A(n133), .B(\u_div/SumTmp[6][12] ), .S0(quotient[6]), .Y(n131)
         );
  MX2X1 U175 ( .A(n134), .B(\u_div/SumTmp[6][13] ), .S0(quotient[6]), .Y(n132)
         );
  MX2X1 U176 ( .A(n101), .B(\u_div/SumTmp[7][11] ), .S0(quotient[7]), .Y(n133)
         );
  MX2X1 U177 ( .A(n123), .B(\u_div/SumTmp[7][12] ), .S0(quotient[7]), .Y(n134)
         );
  MX2X1 U178 ( .A(n106), .B(\u_div/SumTmp[3][11] ), .S0(n2), .Y(n135) );
  MX2X1 U179 ( .A(n124), .B(\u_div/SumTmp[3][12] ), .S0(n2), .Y(n136) );
  MX2X1 U180 ( .A(n125), .B(\u_div/SumTmp[3][13] ), .S0(quotient[3]), .Y(n137)
         );
  MXI2X1 U181 ( .A(n141), .B(\u_div/SumTmp[2][15] ), .S0(quotient[2]), .Y(n174) );
  MXI2X1 U182 ( .A(n137), .B(\u_div/SumTmp[2][14] ), .S0(quotient[2]), .Y(n175) );
  MXI2X1 U183 ( .A(n142), .B(\u_div/SumTmp[2][16] ), .S0(quotient[2]), .Y(n173) );
  MXI2X1 U184 ( .A(n176), .B(n193), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][15] ) );
  INVX1 U185 ( .A(\u_div/SumTmp[1][14] ), .Y(n193) );
  MXI2X1 U186 ( .A(n174), .B(n191), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][17] ) );
  INVX1 U187 ( .A(\u_div/SumTmp[1][16] ), .Y(n191) );
  MX2X1 U188 ( .A(n129), .B(\u_div/SumTmp[4][14] ), .S0(quotient[4]), .Y(n138)
         );
  MX2X1 U189 ( .A(n140), .B(\u_div/SumTmp[4][15] ), .S0(quotient[4]), .Y(n139)
         );
  MX2X1 U190 ( .A(n132), .B(\u_div/SumTmp[5][14] ), .S0(quotient[5]), .Y(n140)
         );
  MX2X1 U191 ( .A(n126), .B(\u_div/SumTmp[3][14] ), .S0(quotient[3]), .Y(n141)
         );
  MX2X1 U192 ( .A(n138), .B(\u_div/SumTmp[3][15] ), .S0(quotient[3]), .Y(n142)
         );
  MX2X1 U193 ( .A(n139), .B(\u_div/SumTmp[3][16] ), .S0(quotient[3]), .Y(n143)
         );
  MXI2X1 U194 ( .A(n143), .B(\u_div/SumTmp[2][17] ), .S0(quotient[2]), .Y(n172) );
  MXI2X1 U195 ( .A(n172), .B(n189), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][19] ) );
  INVX1 U196 ( .A(\u_div/SumTmp[1][18] ), .Y(n189) );
  NAND3BX1 U197 ( .AN(n204), .B(\u_div/BInv [14]), .C(\u_div/CryTmp[6][14] ), 
        .Y(n203) );
  CLKINVX3 U198 ( .A(n199), .Y(quotient[9]) );
  NAND3BX1 U199 ( .AN(n200), .B(\u_div/BInv [11]), .C(\u_div/CryTmp[9][11] ), 
        .Y(n199) );
  CLKINVX3 U200 ( .A(n222), .Y(quotient[12]) );
  NAND3BX1 U201 ( .AN(n221), .B(\u_div/BInv [8]), .C(\u_div/CryTmp[12][8] ), 
        .Y(n222) );
  CLKINVX3 U202 ( .A(n218), .Y(quotient[15]) );
  NAND3BX1 U203 ( .AN(n217), .B(\u_div/BInv [5]), .C(\u_div/CryTmp[15][5] ), 
        .Y(n218) );
  AND2X2 U204 ( .A(\u_div/CryTmp[16][4] ), .B(n216), .Y(quotient[16]) );
  NAND2X1 U205 ( .A(n216), .B(\u_div/BInv [3]), .Y(n213) );
  MXI2X1 U206 ( .A(n7), .B(\u_div/SumTmp[2][1] ), .S0(quotient[2]), .Y(n170)
         );
  NAND2X1 U207 ( .A(n220), .B(\u_div/BInv [6]), .Y(n217) );
  MX2X1 U208 ( .A(n13), .B(\u_div/SumTmp[8][1] ), .S0(quotient[8]), .Y(n145)
         );
  NAND2X1 U209 ( .A(n224), .B(\u_div/BInv [9]), .Y(n221) );
  MX2X1 U210 ( .A(n18), .B(\u_div/SumTmp[10][1] ), .S0(quotient[10]), .Y(n146)
         );
  NAND2X1 U211 ( .A(n202), .B(\u_div/BInv [12]), .Y(n200) );
  NAND2X1 U212 ( .A(n206), .B(\u_div/BInv [15]), .Y(n204) );
  INVX1 U213 ( .A(n214), .Y(quotient[18]) );
  NAND3BX1 U214 ( .AN(n213), .B(\u_div/BInv [2]), .C(\u_div/CryTmp[18][2] ), 
        .Y(n214) );
  MX2X1 U215 ( .A(n20), .B(\u_div/SumTmp[17][1] ), .S0(quotient[17]), .Y(n147)
         );
  MX2X1 U216 ( .A(n9), .B(\u_div/SumTmp[4][1] ), .S0(quotient[4]), .Y(n148) );
  MX2X1 U217 ( .A(n15), .B(\u_div/SumTmp[5][1] ), .S0(quotient[5]), .Y(n149)
         );
  BUFX3 U218 ( .A(n162), .Y(quotient[1]) );
  MX2X1 U219 ( .A(n16), .B(\u_div/SumTmp[6][1] ), .S0(quotient[6]), .Y(n150)
         );
  MX2X1 U220 ( .A(n8), .B(\u_div/SumTmp[7][1] ), .S0(quotient[7]), .Y(n151) );
  MX2X1 U221 ( .A(n11), .B(\u_div/SumTmp[9][1] ), .S0(quotient[9]), .Y(n152)
         );
  MX2X1 U222 ( .A(n17), .B(\u_div/SumTmp[11][1] ), .S0(quotient[11]), .Y(n153)
         );
  MX2X1 U223 ( .A(n12), .B(\u_div/SumTmp[12][1] ), .S0(quotient[12]), .Y(n154)
         );
  MX2X1 U224 ( .A(n23), .B(\u_div/SumTmp[14][1] ), .S0(quotient[14]), .Y(n155)
         );
  MX2X1 U225 ( .A(n21), .B(\u_div/SumTmp[13][1] ), .S0(quotient[13]), .Y(n156)
         );
  MX2X1 U226 ( .A(n19), .B(\u_div/SumTmp[15][1] ), .S0(quotient[15]), .Y(n157)
         );
  MX2X1 U227 ( .A(n22), .B(\u_div/SumTmp[16][1] ), .S0(quotient[16]), .Y(n158)
         );
  MX2X1 U228 ( .A(n14), .B(\u_div/SumTmp[18][1] ), .S0(quotient[18]), .Y(n159)
         );
  MX2X1 U229 ( .A(n10), .B(\u_div/SumTmp[3][1] ), .S0(quotient[3]), .Y(n160)
         );
  AND2X2 U230 ( .A(\u_div/CryTmp[13][7] ), .B(n220), .Y(quotient[13]) );
  INVX1 U231 ( .A(\u_div/CryTmp[2][18] ), .Y(n209) );
  BUFX3 U232 ( .A(n2), .Y(quotient[3]) );
  INVX1 U233 ( .A(n172), .Y(\u_div/PartRem[2][18] ) );
  MXI2X1 U234 ( .A(n171), .B(n188), .S0(quotient[1]), .Y(\u_div/PartRem[1][2] ) );
  INVX1 U235 ( .A(\u_div/SumTmp[1][1] ), .Y(n188) );
  INVX1 U236 ( .A(n170), .Y(\u_div/PartRem[2][2] ) );
  INVX1 U237 ( .A(n169), .Y(\u_div/PartRem[2][3] ) );
  MXI2X1 U238 ( .A(n169), .B(n186), .S0(quotient[1]), .Y(\u_div/PartRem[1][4] ) );
  INVX1 U239 ( .A(\u_div/SumTmp[1][3] ), .Y(n186) );
  INVX1 U240 ( .A(n168), .Y(\u_div/PartRem[2][4] ) );
  INVX1 U241 ( .A(n167), .Y(\u_div/PartRem[2][5] ) );
  INVX1 U242 ( .A(n166), .Y(\u_div/PartRem[2][6] ) );
  MXI2X1 U243 ( .A(n167), .B(n184), .S0(quotient[1]), .Y(\u_div/PartRem[1][6] ) );
  INVX1 U244 ( .A(\u_div/SumTmp[1][5] ), .Y(n184) );
  INVX1 U245 ( .A(n165), .Y(\u_div/PartRem[2][7] ) );
  INVX1 U246 ( .A(n164), .Y(\u_div/PartRem[2][8] ) );
  MXI2X1 U247 ( .A(n165), .B(n182), .S0(quotient[1]), .Y(\u_div/PartRem[1][8] ) );
  INVX1 U248 ( .A(\u_div/SumTmp[1][7] ), .Y(n182) );
  INVX1 U249 ( .A(n163), .Y(\u_div/PartRem[2][9] ) );
  INVX1 U250 ( .A(n180), .Y(\u_div/PartRem[2][10] ) );
  MXI2X1 U251 ( .A(n163), .B(n198), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][10] ) );
  INVX1 U252 ( .A(\u_div/SumTmp[1][9] ), .Y(n198) );
  INVX1 U253 ( .A(n179), .Y(\u_div/PartRem[2][11] ) );
  INVX1 U254 ( .A(n178), .Y(\u_div/PartRem[2][12] ) );
  MXI2X1 U255 ( .A(n179), .B(n196), .S0(n162), .Y(\u_div/PartRem[1][12] ) );
  INVX1 U256 ( .A(\u_div/SumTmp[1][11] ), .Y(n196) );
  INVX1 U257 ( .A(n177), .Y(\u_div/PartRem[2][13] ) );
  MXI2X1 U258 ( .A(n177), .B(n194), .S0(n162), .Y(\u_div/PartRem[1][14] ) );
  INVX1 U259 ( .A(\u_div/SumTmp[1][13] ), .Y(n194) );
  INVX1 U260 ( .A(n176), .Y(\u_div/PartRem[2][14] ) );
  INVX1 U261 ( .A(n175), .Y(\u_div/PartRem[2][15] ) );
  MXI2X1 U262 ( .A(n175), .B(n192), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][16] ) );
  INVX1 U263 ( .A(\u_div/SumTmp[1][15] ), .Y(n192) );
  INVX1 U264 ( .A(n174), .Y(\u_div/PartRem[2][16] ) );
  INVX1 U265 ( .A(n173), .Y(\u_div/PartRem[2][17] ) );
  MXI2X1 U266 ( .A(n173), .B(n190), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][18] ) );
  INVX1 U267 ( .A(\u_div/SumTmp[1][17] ), .Y(n190) );
  NOR3X1 U268 ( .A(n221), .B(b[8]), .C(b[7]), .Y(n220) );
  NOR3X1 U269 ( .A(n217), .B(b[5]), .C(b[4]), .Y(n216) );
  NOR3X1 U270 ( .A(n207), .B(b[17]), .C(b[16]), .Y(n206) );
  NOR3X1 U271 ( .A(n200), .B(b[11]), .C(b[10]), .Y(n224) );
  NOR3X1 U272 ( .A(n204), .B(b[14]), .C(b[13]), .Y(n202) );
  MXI2X1 U273 ( .A(a[2]), .B(\u_div/SumTmp[2][0] ), .S0(quotient[2]), .Y(n171)
         );
  XNOR2X1 U274 ( .A(\u_div/BInv [0]), .B(a[2]), .Y(\u_div/SumTmp[2][0] ) );
  XNOR2X1 U275 ( .A(\u_div/BInv [0]), .B(a[8]), .Y(\u_div/SumTmp[8][0] ) );
  NOR3BX1 U276 ( .AN(\u_div/CryTmp[19][1] ), .B(b[2]), .C(b[1]), .Y(n211) );
  INVX1 U277 ( .A(n213), .Y(n212) );
  XNOR2X1 U278 ( .A(\u_div/BInv [0]), .B(a[10]), .Y(\u_div/SumTmp[10][0] ) );
  OR2X2 U279 ( .A(b[19]), .B(b[18]), .Y(n207) );
  XNOR2X1 U280 ( .A(\u_div/BInv [0]), .B(a[17]), .Y(\u_div/SumTmp[17][0] ) );
  XNOR2X1 U281 ( .A(\u_div/BInv [0]), .B(a[19]), .Y(\u_div/SumTmp[19][0] ) );
  MX2X1 U282 ( .A(a[1]), .B(\u_div/SumTmp[1][0] ), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][1] ) );
  XNOR2X1 U283 ( .A(\u_div/BInv [0]), .B(a[1]), .Y(\u_div/SumTmp[1][0] ) );
  XNOR2X1 U284 ( .A(\u_div/BInv [0]), .B(a[4]), .Y(\u_div/SumTmp[4][0] ) );
  XNOR2X1 U285 ( .A(\u_div/BInv [0]), .B(a[5]), .Y(\u_div/SumTmp[5][0] ) );
  XNOR2X1 U286 ( .A(\u_div/BInv [0]), .B(a[6]), .Y(\u_div/SumTmp[6][0] ) );
  XNOR2X1 U287 ( .A(\u_div/BInv [0]), .B(a[7]), .Y(\u_div/SumTmp[7][0] ) );
  XNOR2X1 U288 ( .A(\u_div/BInv [0]), .B(a[9]), .Y(\u_div/SumTmp[9][0] ) );
  XNOR2X1 U289 ( .A(\u_div/BInv [0]), .B(a[11]), .Y(\u_div/SumTmp[11][0] ) );
  XNOR2X1 U290 ( .A(\u_div/BInv [0]), .B(a[12]), .Y(\u_div/SumTmp[12][0] ) );
  XNOR2X1 U291 ( .A(\u_div/BInv [0]), .B(a[14]), .Y(\u_div/SumTmp[14][0] ) );
  XNOR2X1 U292 ( .A(\u_div/BInv [0]), .B(a[13]), .Y(\u_div/SumTmp[13][0] ) );
  XNOR2X1 U293 ( .A(\u_div/BInv [0]), .B(a[15]), .Y(\u_div/SumTmp[15][0] ) );
  XNOR2X1 U294 ( .A(\u_div/BInv [0]), .B(a[16]), .Y(\u_div/SumTmp[16][0] ) );
  XNOR2X1 U295 ( .A(\u_div/BInv [0]), .B(a[3]), .Y(\u_div/SumTmp[3][0] ) );
  XNOR2X1 U296 ( .A(\u_div/BInv [0]), .B(a[18]), .Y(\u_div/SumTmp[18][0] ) );
  OR2X2 U297 ( .A(a[1]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[1][1] ) );
  INVX1 U298 ( .A(n171), .Y(\u_div/PartRem[2][1] ) );
  INVX1 U299 ( .A(\u_div/CryTmp[3][17] ), .Y(n208) );
  INVX1 U300 ( .A(n210), .Y(n162) );
  NAND2BX1 U301 ( .AN(b[19]), .B(\u_div/CryTmp[1][19] ), .Y(n210) );
  OR2X2 U302 ( .A(a[18]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[18][1] ) );
  OR2X2 U303 ( .A(a[17]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[17][1] ) );
  OR2X2 U304 ( .A(a[16]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[16][1] ) );
  OR2X2 U305 ( .A(a[15]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[15][1] ) );
  OR2X2 U306 ( .A(a[14]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[14][1] ) );
  OR2X2 U307 ( .A(a[13]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[13][1] ) );
  OR2X2 U308 ( .A(a[12]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[12][1] ) );
  OR2X2 U309 ( .A(a[11]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[11][1] ) );
  OR2X2 U310 ( .A(a[10]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[10][1] ) );
  OR2X2 U311 ( .A(a[9]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[9][1] ) );
  OR2X2 U312 ( .A(a[8]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[8][1] ) );
  OR2X2 U313 ( .A(a[7]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[7][1] ) );
  OR2X2 U314 ( .A(a[6]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[6][1] ) );
  OR2X2 U315 ( .A(a[5]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[5][1] ) );
  OR2X2 U316 ( .A(a[4]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[4][1] ) );
  OR2X2 U317 ( .A(a[3]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[3][1] ) );
  OR2X2 U318 ( .A(a[2]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[2][1] ) );
  CLKINVX3 U319 ( .A(b[12]), .Y(\u_div/BInv [12]) );
  CLKINVX3 U320 ( .A(b[15]), .Y(\u_div/BInv [15]) );
  CLKINVX3 U321 ( .A(b[9]), .Y(\u_div/BInv [9]) );
  OR2X2 U322 ( .A(a[19]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[19][1] ) );
  CLKINVX3 U323 ( .A(b[10]), .Y(\u_div/BInv [10]) );
  CLKINVX3 U324 ( .A(b[11]), .Y(\u_div/BInv [11]) );
  CLKINVX3 U325 ( .A(b[13]), .Y(\u_div/BInv [13]) );
  CLKINVX3 U326 ( .A(b[14]), .Y(\u_div/BInv [14]) );
  INVX1 U327 ( .A(b[16]), .Y(\u_div/BInv [16]) );
  INVX1 U328 ( .A(b[17]), .Y(\u_div/BInv [17]) );
  OR2X2 U329 ( .A(a[0]), .B(\u_div/BInv [0]), .Y(\u_div/CryTmp[0][1] ) );
  INVX1 U330 ( .A(b[18]), .Y(\u_div/BInv [18]) );
  INVX1 U331 ( .A(b[19]), .Y(\u_div/BInv [19]) );
  CLKINVX8 U332 ( .A(b[0]), .Y(\u_div/BInv [0]) );
  CLKINVX4 U333 ( .A(n205), .Y(quotient[5]) );
endmodule


module Control_And_Registers ( clk, rst, ena_in, Address, data_in, ena_out, 
        Image_Done, Block_Done, params, Im_block, W_block );
  input [9:0] Address;
  input [15:0] data_in;
  output [46:0] params;
  output [31:0] Im_block;
  output [31:0] W_block;
  input clk, rst, ena_in, Block_Done;
  output ena_out, Image_Done;
  wire   N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N84, N85, N86, N87, \registers[31][7] , \registers[31][6] ,
         \registers[31][5] , \registers[31][4] , \registers[31][3] ,
         \registers[31][2] , \registers[31][1] , \registers[31][0] ,
         \registers[30][7] , \registers[30][6] , \registers[30][5] ,
         \registers[30][4] , \registers[30][3] , \registers[30][2] ,
         \registers[30][1] , \registers[30][0] , \registers[29][7] ,
         \registers[29][6] , \registers[29][5] , \registers[29][4] ,
         \registers[29][3] , \registers[29][2] , \registers[29][1] ,
         \registers[29][0] , \registers[28][7] , \registers[28][6] ,
         \registers[28][5] , \registers[28][4] , \registers[28][3] ,
         \registers[28][2] , \registers[28][1] , \registers[28][0] ,
         \registers[27][7] , \registers[27][6] , \registers[27][5] ,
         \registers[27][4] , \registers[27][3] , \registers[27][2] ,
         \registers[27][1] , \registers[27][0] , \registers[26][7] ,
         \registers[26][6] , \registers[26][5] , \registers[26][4] ,
         \registers[26][3] , \registers[26][2] , \registers[26][1] ,
         \registers[26][0] , \registers[25][7] , \registers[25][6] ,
         \registers[25][5] , \registers[25][4] , \registers[25][3] ,
         \registers[25][2] , \registers[25][1] , \registers[25][0] ,
         \registers[24][7] , \registers[24][6] , \registers[24][5] ,
         \registers[24][4] , \registers[24][3] , \registers[24][2] ,
         \registers[24][1] , \registers[24][0] , \registers[23][7] ,
         \registers[23][6] , \registers[23][5] , \registers[23][4] ,
         \registers[23][3] , \registers[23][2] , \registers[23][1] ,
         \registers[23][0] , \registers[22][7] , \registers[22][6] ,
         \registers[22][5] , \registers[22][4] , \registers[22][3] ,
         \registers[22][2] , \registers[22][1] , \registers[22][0] ,
         \registers[21][7] , \registers[21][6] , \registers[21][5] ,
         \registers[21][4] , \registers[21][3] , \registers[21][2] ,
         \registers[21][1] , \registers[21][0] , \registers[20][7] ,
         \registers[20][6] , \registers[20][5] , \registers[20][4] ,
         \registers[20][3] , \registers[20][2] , \registers[20][1] ,
         \registers[20][0] , \registers[19][7] , \registers[19][6] ,
         \registers[19][5] , \registers[19][4] , \registers[19][3] ,
         \registers[19][2] , \registers[19][1] , \registers[19][0] ,
         \registers[18][7] , \registers[18][6] , \registers[18][5] ,
         \registers[18][4] , \registers[18][3] , \registers[18][2] ,
         \registers[18][1] , \registers[18][0] , \registers[17][7] ,
         \registers[17][6] , \registers[17][5] , \registers[17][4] ,
         \registers[17][3] , \registers[17][2] , \registers[17][1] ,
         \registers[17][0] , \registers[16][7] , \registers[16][6] ,
         \registers[16][5] , \registers[16][4] , \registers[16][3] ,
         \registers[16][2] , \registers[16][1] , \registers[16][0] ,
         \registers[15][7] , \registers[15][6] , \registers[15][5] ,
         \registers[15][4] , \registers[15][3] , \registers[15][2] ,
         \registers[15][1] , \registers[15][0] , \registers[14][7] ,
         \registers[14][6] , \registers[14][5] , \registers[14][4] ,
         \registers[14][3] , \registers[14][2] , \registers[14][1] ,
         \registers[14][0] , \registers[13][7] , \registers[13][6] ,
         \registers[13][5] , \registers[13][4] , \registers[13][3] ,
         \registers[13][2] , \registers[13][1] , \registers[13][0] ,
         \registers[12][7] , \registers[12][6] , \registers[12][5] ,
         \registers[12][4] , \registers[12][3] , \registers[12][2] ,
         \registers[12][1] , \registers[12][0] , \registers[11][7] ,
         \registers[11][6] , \registers[11][5] , \registers[11][4] ,
         \registers[11][3] , \registers[11][2] , \registers[11][1] ,
         \registers[11][0] , \registers[10][7] , \registers[10][6] ,
         \registers[10][5] , \registers[10][4] , \registers[10][3] ,
         \registers[10][2] , \registers[10][1] , \registers[10][0] ,
         \registers[9][7] , \registers[9][6] , \registers[9][5] ,
         \registers[9][4] , \registers[9][3] , \registers[9][2] ,
         \registers[9][1] , \registers[9][0] , \registers[8][7] ,
         \registers[8][6] , \registers[8][5] , \registers[8][4] ,
         \registers[8][3] , \registers[8][2] , \registers[8][1] ,
         \registers[8][0] , \registers[7][7] , \registers[7][6] ,
         \registers[7][5] , \registers[7][4] , \registers[7][3] ,
         \registers[7][2] , \registers[7][1] , \registers[7][0] ,
         \registers[6][7] , \registers[6][6] , \registers[6][5] ,
         \registers[6][4] , \registers[6][3] , \registers[6][2] ,
         \registers[6][1] , \registers[6][0] , \registers[5][7] ,
         \registers[5][6] , \registers[5][5] , \registers[5][4] ,
         \registers[5][3] , \registers[5][2] , \registers[5][1] ,
         \registers[5][0] , \registers[4][7] , \registers[4][6] ,
         \registers[4][5] , \registers[4][4] , \registers[4][3] ,
         \registers[4][2] , \registers[4][1] , \registers[4][0] ,
         \registers[3][7] , \registers[3][6] , \registers[3][5] ,
         \registers[3][4] , \registers[3][3] , \registers[3][2] ,
         \registers[3][1] , \registers[3][0] , \registers[2][7] ,
         \registers[2][6] , \registers[2][5] , \registers[2][4] ,
         \registers[2][3] , \registers[2][2] , \registers[2][1] ,
         \registers[2][0] , \registers[1][7] , \registers[1][6] ,
         \registers[1][5] , \registers[1][4] , \registers[1][3] ,
         \registers[1][2] , \registers[1][1] , \registers[1][0] ,
         \registers[0][7] , \registers[0][6] , \registers[0][5] ,
         \registers[0][4] , \registers[0][3] , \registers[0][2] ,
         \registers[0][1] , \registers[0][0] , \registers[63][7] ,
         \registers[63][6] , \registers[63][5] , \registers[63][4] ,
         \registers[63][3] , \registers[63][2] , \registers[63][1] ,
         \registers[63][0] , \registers[62][7] , \registers[62][6] ,
         \registers[62][5] , \registers[62][4] , \registers[62][3] ,
         \registers[62][2] , \registers[62][1] , \registers[62][0] ,
         \registers[61][7] , \registers[61][6] , \registers[61][5] ,
         \registers[61][4] , \registers[61][3] , \registers[61][2] ,
         \registers[61][1] , \registers[61][0] , \registers[60][7] ,
         \registers[60][6] , \registers[60][5] , \registers[60][4] ,
         \registers[60][3] , \registers[60][2] , \registers[60][1] ,
         \registers[60][0] , \registers[59][7] , \registers[59][6] ,
         \registers[59][5] , \registers[59][4] , \registers[59][3] ,
         \registers[59][2] , \registers[59][1] , \registers[59][0] ,
         \registers[58][7] , \registers[58][6] , \registers[58][5] ,
         \registers[58][4] , \registers[58][3] , \registers[58][2] ,
         \registers[58][1] , \registers[58][0] , \registers[57][7] ,
         \registers[57][6] , \registers[57][5] , \registers[57][4] ,
         \registers[57][3] , \registers[57][2] , \registers[57][1] ,
         \registers[57][0] , \registers[56][7] , \registers[56][6] ,
         \registers[56][5] , \registers[56][4] , \registers[56][3] ,
         \registers[56][2] , \registers[56][1] , \registers[56][0] ,
         \registers[55][7] , \registers[55][6] , \registers[55][5] ,
         \registers[55][4] , \registers[55][3] , \registers[55][2] ,
         \registers[55][1] , \registers[55][0] , \registers[54][7] ,
         \registers[54][6] , \registers[54][5] , \registers[54][4] ,
         \registers[54][3] , \registers[54][2] , \registers[54][1] ,
         \registers[54][0] , \registers[53][7] , \registers[53][6] ,
         \registers[53][5] , \registers[53][4] , \registers[53][3] ,
         \registers[53][2] , \registers[53][1] , \registers[53][0] ,
         \registers[52][7] , \registers[52][6] , \registers[52][5] ,
         \registers[52][4] , \registers[52][3] , \registers[52][2] ,
         \registers[52][1] , \registers[52][0] , \registers[51][7] ,
         \registers[51][6] , \registers[51][5] , \registers[51][4] ,
         \registers[51][3] , \registers[51][2] , \registers[51][1] ,
         \registers[51][0] , \registers[50][7] , \registers[50][6] ,
         \registers[50][5] , \registers[50][4] , \registers[50][3] ,
         \registers[50][2] , \registers[50][1] , \registers[50][0] ,
         \registers[49][7] , \registers[49][6] , \registers[49][5] ,
         \registers[49][4] , \registers[49][3] , \registers[49][2] ,
         \registers[49][1] , \registers[49][0] , \registers[48][7] ,
         \registers[48][6] , \registers[48][5] , \registers[48][4] ,
         \registers[48][3] , \registers[48][2] , \registers[48][1] ,
         \registers[48][0] , \registers[47][7] , \registers[47][6] ,
         \registers[47][5] , \registers[47][4] , \registers[47][3] ,
         \registers[47][2] , \registers[47][1] , \registers[47][0] ,
         \registers[46][7] , \registers[46][6] , \registers[46][5] ,
         \registers[46][4] , \registers[46][3] , \registers[46][2] ,
         \registers[46][1] , \registers[46][0] , \registers[45][7] ,
         \registers[45][6] , \registers[45][5] , \registers[45][4] ,
         \registers[45][3] , \registers[45][2] , \registers[45][1] ,
         \registers[45][0] , \registers[44][7] , \registers[44][6] ,
         \registers[44][5] , \registers[44][4] , \registers[44][3] ,
         \registers[44][2] , \registers[44][1] , \registers[44][0] ,
         \registers[43][7] , \registers[43][6] , \registers[43][5] ,
         \registers[43][4] , \registers[43][3] , \registers[43][2] ,
         \registers[43][1] , \registers[43][0] , \registers[42][7] ,
         \registers[42][6] , \registers[42][5] , \registers[42][4] ,
         \registers[42][3] , \registers[42][2] , \registers[42][1] ,
         \registers[42][0] , \registers[41][7] , \registers[41][6] ,
         \registers[41][5] , \registers[41][4] , \registers[41][3] ,
         \registers[41][2] , \registers[41][1] , \registers[41][0] ,
         \registers[40][7] , \registers[40][6] , \registers[40][5] ,
         \registers[40][4] , \registers[40][3] , \registers[40][2] ,
         \registers[40][1] , \registers[40][0] , \registers[39][7] ,
         \registers[39][6] , \registers[39][5] , \registers[39][4] ,
         \registers[39][3] , \registers[39][2] , \registers[39][1] ,
         \registers[39][0] , \registers[38][7] , \registers[38][6] ,
         \registers[38][5] , \registers[38][4] , \registers[38][3] ,
         \registers[38][2] , \registers[38][1] , \registers[38][0] ,
         \registers[37][7] , \registers[37][6] , \registers[37][5] ,
         \registers[37][4] , \registers[37][3] , \registers[37][2] ,
         \registers[37][1] , \registers[37][0] , \registers[36][7] ,
         \registers[36][6] , \registers[36][5] , \registers[36][4] ,
         \registers[36][3] , \registers[36][2] , \registers[36][1] ,
         \registers[36][0] , \registers[35][7] , \registers[35][6] ,
         \registers[35][5] , \registers[35][4] , \registers[35][3] ,
         \registers[35][2] , \registers[35][1] , \registers[35][0] ,
         \registers[34][7] , \registers[34][6] , \registers[34][5] ,
         \registers[34][4] , \registers[34][3] , \registers[34][2] ,
         \registers[34][1] , \registers[34][0] , \registers[33][7] ,
         \registers[33][6] , \registers[33][5] , \registers[33][4] ,
         \registers[33][3] , \registers[33][2] , \registers[33][1] ,
         \registers[33][0] , \registers[32][7] , \registers[32][6] ,
         \registers[32][5] , \registers[32][4] , \registers[32][3] ,
         \registers[32][2] , \registers[32][1] , \registers[32][0] ,
         \registers[95][7] , \registers[95][6] , \registers[95][5] ,
         \registers[95][4] , \registers[95][3] , \registers[95][2] ,
         \registers[95][1] , \registers[95][0] , \registers[94][7] ,
         \registers[94][6] , \registers[94][5] , \registers[94][4] ,
         \registers[94][3] , \registers[94][2] , \registers[94][1] ,
         \registers[94][0] , \registers[93][7] , \registers[93][6] ,
         \registers[93][5] , \registers[93][4] , \registers[93][3] ,
         \registers[93][2] , \registers[93][1] , \registers[93][0] ,
         \registers[92][7] , \registers[92][6] , \registers[92][5] ,
         \registers[92][4] , \registers[92][3] , \registers[92][2] ,
         \registers[92][1] , \registers[92][0] , \registers[91][7] ,
         \registers[91][6] , \registers[91][5] , \registers[91][4] ,
         \registers[91][3] , \registers[91][2] , \registers[91][1] ,
         \registers[91][0] , \registers[90][7] , \registers[90][6] ,
         \registers[90][5] , \registers[90][4] , \registers[90][3] ,
         \registers[90][2] , \registers[90][1] , \registers[90][0] ,
         \registers[89][7] , \registers[89][6] , \registers[89][5] ,
         \registers[89][4] , \registers[89][3] , \registers[89][2] ,
         \registers[89][1] , \registers[89][0] , \registers[88][7] ,
         \registers[88][6] , \registers[88][5] , \registers[88][4] ,
         \registers[88][3] , \registers[88][2] , \registers[88][1] ,
         \registers[88][0] , \registers[87][7] , \registers[87][6] ,
         \registers[87][5] , \registers[87][4] , \registers[87][3] ,
         \registers[87][2] , \registers[87][1] , \registers[87][0] ,
         \registers[86][7] , \registers[86][6] , \registers[86][5] ,
         \registers[86][4] , \registers[86][3] , \registers[86][2] ,
         \registers[86][1] , \registers[86][0] , \registers[85][7] ,
         \registers[85][6] , \registers[85][5] , \registers[85][4] ,
         \registers[85][3] , \registers[85][2] , \registers[85][1] ,
         \registers[85][0] , \registers[84][7] , \registers[84][6] ,
         \registers[84][5] , \registers[84][4] , \registers[84][3] ,
         \registers[84][2] , \registers[84][1] , \registers[84][0] ,
         \registers[83][7] , \registers[83][6] , \registers[83][5] ,
         \registers[83][4] , \registers[83][3] , \registers[83][2] ,
         \registers[83][1] , \registers[83][0] , \registers[82][7] ,
         \registers[82][6] , \registers[82][5] , \registers[82][4] ,
         \registers[82][3] , \registers[82][2] , \registers[82][1] ,
         \registers[82][0] , \registers[81][7] , \registers[81][6] ,
         \registers[81][5] , \registers[81][4] , \registers[81][3] ,
         \registers[81][2] , \registers[81][1] , \registers[81][0] ,
         \registers[80][7] , \registers[80][6] , \registers[80][5] ,
         \registers[80][4] , \registers[80][3] , \registers[80][2] ,
         \registers[80][1] , \registers[80][0] , \registers[79][7] ,
         \registers[79][6] , \registers[79][5] , \registers[79][4] ,
         \registers[79][3] , \registers[79][2] , \registers[79][1] ,
         \registers[79][0] , \registers[78][7] , \registers[78][6] ,
         \registers[78][5] , \registers[78][4] , \registers[78][3] ,
         \registers[78][2] , \registers[78][1] , \registers[78][0] ,
         \registers[77][7] , \registers[77][6] , \registers[77][5] ,
         \registers[77][4] , \registers[77][3] , \registers[77][2] ,
         \registers[77][1] , \registers[77][0] , \registers[76][7] ,
         \registers[76][6] , \registers[76][5] , \registers[76][4] ,
         \registers[76][3] , \registers[76][2] , \registers[76][1] ,
         \registers[76][0] , \registers[75][7] , \registers[75][6] ,
         \registers[75][5] , \registers[75][4] , \registers[75][3] ,
         \registers[75][2] , \registers[75][1] , \registers[75][0] ,
         \registers[74][7] , \registers[74][6] , \registers[74][5] ,
         \registers[74][4] , \registers[74][3] , \registers[74][2] ,
         \registers[74][1] , \registers[74][0] , \registers[73][7] ,
         \registers[73][6] , \registers[73][5] , \registers[73][4] ,
         \registers[73][3] , \registers[73][2] , \registers[73][1] ,
         \registers[73][0] , \registers[72][7] , \registers[72][6] ,
         \registers[72][5] , \registers[72][4] , \registers[72][3] ,
         \registers[72][2] , \registers[72][1] , \registers[72][0] ,
         \registers[71][7] , \registers[71][6] , \registers[71][5] ,
         \registers[71][4] , \registers[71][3] , \registers[71][2] ,
         \registers[71][1] , \registers[71][0] , \registers[70][7] ,
         \registers[70][6] , \registers[70][5] , \registers[70][4] ,
         \registers[70][3] , \registers[70][2] , \registers[70][1] ,
         \registers[70][0] , \registers[69][7] , \registers[69][6] ,
         \registers[69][5] , \registers[69][4] , \registers[69][3] ,
         \registers[69][2] , \registers[69][1] , \registers[69][0] ,
         \registers[68][7] , \registers[68][6] , \registers[68][5] ,
         \registers[68][4] , \registers[68][3] , \registers[68][2] ,
         \registers[68][1] , \registers[68][0] , \registers[67][7] ,
         \registers[67][6] , \registers[67][5] , \registers[67][4] ,
         \registers[67][3] , \registers[67][2] , \registers[67][1] ,
         \registers[67][0] , \registers[66][7] , \registers[66][6] ,
         \registers[66][5] , \registers[66][4] , \registers[66][3] ,
         \registers[66][2] , \registers[66][1] , \registers[66][0] ,
         \registers[65][7] , \registers[65][6] , \registers[65][5] ,
         \registers[65][4] , \registers[65][3] , \registers[65][2] ,
         \registers[65][1] , \registers[65][0] , \registers[64][7] ,
         \registers[64][6] , \registers[64][5] , \registers[64][4] ,
         \registers[64][3] , \registers[64][2] , \registers[64][1] ,
         \registers[64][0] , \registers[127][7] , \registers[127][6] ,
         \registers[127][5] , \registers[127][4] , \registers[127][3] ,
         \registers[127][2] , \registers[127][1] , \registers[127][0] ,
         \registers[126][7] , \registers[126][6] , \registers[126][5] ,
         \registers[126][4] , \registers[126][3] , \registers[126][2] ,
         \registers[126][1] , \registers[126][0] , \registers[125][7] ,
         \registers[125][6] , \registers[125][5] , \registers[125][4] ,
         \registers[125][3] , \registers[125][2] , \registers[125][1] ,
         \registers[125][0] , \registers[124][7] , \registers[124][6] ,
         \registers[124][5] , \registers[124][4] , \registers[124][3] ,
         \registers[124][2] , \registers[124][1] , \registers[124][0] ,
         \registers[123][7] , \registers[123][6] , \registers[123][5] ,
         \registers[123][4] , \registers[123][3] , \registers[123][2] ,
         \registers[123][1] , \registers[123][0] , \registers[122][7] ,
         \registers[122][6] , \registers[122][5] , \registers[122][4] ,
         \registers[122][3] , \registers[122][2] , \registers[122][1] ,
         \registers[122][0] , \registers[121][7] , \registers[121][6] ,
         \registers[121][5] , \registers[121][4] , \registers[121][3] ,
         \registers[121][2] , \registers[121][1] , \registers[121][0] ,
         \registers[120][7] , \registers[120][6] , \registers[120][5] ,
         \registers[120][4] , \registers[120][3] , \registers[120][2] ,
         \registers[120][1] , \registers[120][0] , \registers[119][7] ,
         \registers[119][6] , \registers[119][5] , \registers[119][4] ,
         \registers[119][3] , \registers[119][2] , \registers[119][1] ,
         \registers[119][0] , \registers[118][7] , \registers[118][6] ,
         \registers[118][5] , \registers[118][4] , \registers[118][3] ,
         \registers[118][2] , \registers[118][1] , \registers[118][0] ,
         \registers[117][7] , \registers[117][6] , \registers[117][5] ,
         \registers[117][4] , \registers[117][3] , \registers[117][2] ,
         \registers[117][1] , \registers[117][0] , \registers[116][7] ,
         \registers[116][6] , \registers[116][5] , \registers[116][4] ,
         \registers[116][3] , \registers[116][2] , \registers[116][1] ,
         \registers[116][0] , \registers[115][7] , \registers[115][6] ,
         \registers[115][5] , \registers[115][4] , \registers[115][3] ,
         \registers[115][2] , \registers[115][1] , \registers[115][0] ,
         \registers[114][7] , \registers[114][6] , \registers[114][5] ,
         \registers[114][4] , \registers[114][3] , \registers[114][2] ,
         \registers[114][1] , \registers[114][0] , \registers[113][7] ,
         \registers[113][6] , \registers[113][5] , \registers[113][4] ,
         \registers[113][3] , \registers[113][2] , \registers[113][1] ,
         \registers[113][0] , \registers[112][7] , \registers[112][6] ,
         \registers[112][5] , \registers[112][4] , \registers[112][3] ,
         \registers[112][2] , \registers[112][1] , \registers[112][0] ,
         \registers[111][7] , \registers[111][6] , \registers[111][5] ,
         \registers[111][4] , \registers[111][3] , \registers[111][2] ,
         \registers[111][1] , \registers[111][0] , \registers[110][7] ,
         \registers[110][6] , \registers[110][5] , \registers[110][4] ,
         \registers[110][3] , \registers[110][2] , \registers[110][1] ,
         \registers[110][0] , \registers[109][7] , \registers[109][6] ,
         \registers[109][5] , \registers[109][4] , \registers[109][3] ,
         \registers[109][2] , \registers[109][1] , \registers[109][0] ,
         \registers[108][7] , \registers[108][6] , \registers[108][5] ,
         \registers[108][4] , \registers[108][3] , \registers[108][2] ,
         \registers[108][1] , \registers[108][0] , \registers[107][7] ,
         \registers[107][6] , \registers[107][5] , \registers[107][4] ,
         \registers[107][3] , \registers[107][2] , \registers[107][1] ,
         \registers[107][0] , \registers[106][7] , \registers[106][6] ,
         \registers[106][5] , \registers[106][4] , \registers[106][3] ,
         \registers[106][2] , \registers[106][1] , \registers[106][0] ,
         \registers[105][7] , \registers[105][6] , \registers[105][5] ,
         \registers[105][4] , \registers[105][3] , \registers[105][2] ,
         \registers[105][1] , \registers[105][0] , \registers[104][7] ,
         \registers[104][6] , \registers[104][5] , \registers[104][4] ,
         \registers[104][3] , \registers[104][2] , \registers[104][1] ,
         \registers[104][0] , \registers[103][7] , \registers[103][6] ,
         \registers[103][5] , \registers[103][4] , \registers[103][3] ,
         \registers[103][2] , \registers[103][1] , \registers[103][0] ,
         \registers[102][7] , \registers[102][6] , \registers[102][5] ,
         \registers[102][4] , \registers[102][3] , \registers[102][2] ,
         \registers[102][1] , \registers[102][0] , \registers[101][7] ,
         \registers[101][6] , \registers[101][5] , \registers[101][4] ,
         \registers[101][3] , \registers[101][2] , \registers[101][1] ,
         \registers[101][0] , \registers[100][7] , \registers[100][6] ,
         \registers[100][5] , \registers[100][4] , \registers[100][3] ,
         \registers[100][2] , \registers[100][1] , \registers[100][0] ,
         \registers[99][7] , \registers[99][6] , \registers[99][5] ,
         \registers[99][4] , \registers[99][3] , \registers[99][2] ,
         \registers[99][1] , \registers[99][0] , \registers[98][7] ,
         \registers[98][6] , \registers[98][5] , \registers[98][4] ,
         \registers[98][3] , \registers[98][2] , \registers[98][1] ,
         \registers[98][0] , \registers[97][7] , \registers[97][6] ,
         \registers[97][5] , \registers[97][4] , \registers[97][3] ,
         \registers[97][2] , \registers[97][1] , \registers[97][0] ,
         \registers[96][7] , \registers[96][6] , \registers[96][5] ,
         \registers[96][4] , \registers[96][3] , \registers[96][2] ,
         \registers[96][1] , \registers[96][0] , \registers[159][7] ,
         \registers[159][6] , \registers[159][5] , \registers[159][4] ,
         \registers[159][3] , \registers[159][2] , \registers[159][1] ,
         \registers[159][0] , \registers[158][7] , \registers[158][6] ,
         \registers[158][5] , \registers[158][4] , \registers[158][3] ,
         \registers[158][2] , \registers[158][1] , \registers[158][0] ,
         \registers[157][7] , \registers[157][6] , \registers[157][5] ,
         \registers[157][4] , \registers[157][3] , \registers[157][2] ,
         \registers[157][1] , \registers[157][0] , \registers[156][7] ,
         \registers[156][6] , \registers[156][5] , \registers[156][4] ,
         \registers[156][3] , \registers[156][2] , \registers[156][1] ,
         \registers[156][0] , \registers[155][7] , \registers[155][6] ,
         \registers[155][5] , \registers[155][4] , \registers[155][3] ,
         \registers[155][2] , \registers[155][1] , \registers[155][0] ,
         \registers[154][7] , \registers[154][6] , \registers[154][5] ,
         \registers[154][4] , \registers[154][3] , \registers[154][2] ,
         \registers[154][1] , \registers[154][0] , \registers[153][7] ,
         \registers[153][6] , \registers[153][5] , \registers[153][4] ,
         \registers[153][3] , \registers[153][2] , \registers[153][1] ,
         \registers[153][0] , \registers[152][7] , \registers[152][6] ,
         \registers[152][5] , \registers[152][4] , \registers[152][3] ,
         \registers[152][2] , \registers[152][1] , \registers[152][0] ,
         \registers[151][7] , \registers[151][6] , \registers[151][5] ,
         \registers[151][4] , \registers[151][3] , \registers[151][2] ,
         \registers[151][1] , \registers[151][0] , \registers[150][7] ,
         \registers[150][6] , \registers[150][5] , \registers[150][4] ,
         \registers[150][3] , \registers[150][2] , \registers[150][1] ,
         \registers[150][0] , \registers[149][7] , \registers[149][6] ,
         \registers[149][5] , \registers[149][4] , \registers[149][3] ,
         \registers[149][2] , \registers[149][1] , \registers[149][0] ,
         \registers[148][7] , \registers[148][6] , \registers[148][5] ,
         \registers[148][4] , \registers[148][3] , \registers[148][2] ,
         \registers[148][1] , \registers[148][0] , \registers[147][7] ,
         \registers[147][6] , \registers[147][5] , \registers[147][4] ,
         \registers[147][3] , \registers[147][2] , \registers[147][1] ,
         \registers[147][0] , \registers[146][7] , \registers[146][6] ,
         \registers[146][5] , \registers[146][4] , \registers[146][3] ,
         \registers[146][2] , \registers[146][1] , \registers[146][0] ,
         \registers[145][7] , \registers[145][6] , \registers[145][5] ,
         \registers[145][4] , \registers[145][3] , \registers[145][2] ,
         \registers[145][1] , \registers[145][0] , \registers[144][7] ,
         \registers[144][6] , \registers[144][5] , \registers[144][4] ,
         \registers[144][3] , \registers[144][2] , \registers[144][1] ,
         \registers[144][0] , \registers[143][7] , \registers[143][6] ,
         \registers[143][5] , \registers[143][4] , \registers[143][3] ,
         \registers[143][2] , \registers[143][1] , \registers[143][0] ,
         \registers[142][7] , \registers[142][6] , \registers[142][5] ,
         \registers[142][4] , \registers[142][3] , \registers[142][2] ,
         \registers[142][1] , \registers[142][0] , \registers[141][7] ,
         \registers[141][6] , \registers[141][5] , \registers[141][4] ,
         \registers[141][3] , \registers[141][2] , \registers[141][1] ,
         \registers[141][0] , \registers[140][7] , \registers[140][6] ,
         \registers[140][5] , \registers[140][4] , \registers[140][3] ,
         \registers[140][2] , \registers[140][1] , \registers[140][0] ,
         \registers[139][7] , \registers[139][6] , \registers[139][5] ,
         \registers[139][4] , \registers[139][3] , \registers[139][2] ,
         \registers[139][1] , \registers[139][0] , \registers[138][7] ,
         \registers[138][6] , \registers[138][5] , \registers[138][4] ,
         \registers[138][3] , \registers[138][2] , \registers[138][1] ,
         \registers[138][0] , \registers[137][7] , \registers[137][6] ,
         \registers[137][5] , \registers[137][4] , \registers[137][3] ,
         \registers[137][2] , \registers[137][1] , \registers[137][0] ,
         \registers[136][7] , \registers[136][6] , \registers[136][5] ,
         \registers[136][4] , \registers[136][3] , \registers[136][2] ,
         \registers[136][1] , \registers[136][0] , \registers[135][7] ,
         \registers[135][6] , \registers[135][5] , \registers[135][4] ,
         \registers[135][3] , \registers[135][2] , \registers[135][1] ,
         \registers[135][0] , \registers[134][7] , \registers[134][6] ,
         \registers[134][5] , \registers[134][4] , \registers[134][3] ,
         \registers[134][2] , \registers[134][1] , \registers[134][0] ,
         \registers[133][7] , \registers[133][6] , \registers[133][5] ,
         \registers[133][4] , \registers[133][3] , \registers[133][2] ,
         \registers[133][1] , \registers[133][0] , \registers[132][7] ,
         \registers[132][6] , \registers[132][5] , \registers[132][4] ,
         \registers[132][3] , \registers[132][2] , \registers[132][1] ,
         \registers[132][0] , \registers[131][7] , \registers[131][6] ,
         \registers[131][5] , \registers[131][4] , \registers[131][3] ,
         \registers[131][2] , \registers[131][1] , \registers[131][0] ,
         \registers[130][7] , \registers[130][6] , \registers[130][5] ,
         \registers[130][4] , \registers[130][3] , \registers[130][2] ,
         \registers[130][1] , \registers[130][0] , \registers[129][7] ,
         \registers[129][6] , \registers[129][5] , \registers[129][4] ,
         \registers[129][3] , \registers[129][2] , \registers[129][1] ,
         \registers[129][0] , \registers[128][7] , \registers[128][6] ,
         \registers[128][5] , \registers[128][4] , \registers[128][3] ,
         \registers[128][2] , \registers[128][1] , \registers[128][0] ,
         \registers[191][7] , \registers[191][6] , \registers[191][5] ,
         \registers[191][4] , \registers[191][3] , \registers[191][2] ,
         \registers[191][1] , \registers[191][0] , \registers[190][7] ,
         \registers[190][6] , \registers[190][5] , \registers[190][4] ,
         \registers[190][3] , \registers[190][2] , \registers[190][1] ,
         \registers[190][0] , \registers[189][7] , \registers[189][6] ,
         \registers[189][5] , \registers[189][4] , \registers[189][3] ,
         \registers[189][2] , \registers[189][1] , \registers[189][0] ,
         \registers[188][7] , \registers[188][6] , \registers[188][5] ,
         \registers[188][4] , \registers[188][3] , \registers[188][2] ,
         \registers[188][1] , \registers[188][0] , \registers[187][7] ,
         \registers[187][6] , \registers[187][5] , \registers[187][4] ,
         \registers[187][3] , \registers[187][2] , \registers[187][1] ,
         \registers[187][0] , \registers[186][7] , \registers[186][6] ,
         \registers[186][5] , \registers[186][4] , \registers[186][3] ,
         \registers[186][2] , \registers[186][1] , \registers[186][0] ,
         \registers[185][7] , \registers[185][6] , \registers[185][5] ,
         \registers[185][4] , \registers[185][3] , \registers[185][2] ,
         \registers[185][1] , \registers[185][0] , \registers[184][7] ,
         \registers[184][6] , \registers[184][5] , \registers[184][4] ,
         \registers[184][3] , \registers[184][2] , \registers[184][1] ,
         \registers[184][0] , \registers[183][7] , \registers[183][6] ,
         \registers[183][5] , \registers[183][4] , \registers[183][3] ,
         \registers[183][2] , \registers[183][1] , \registers[183][0] ,
         \registers[182][7] , \registers[182][6] , \registers[182][5] ,
         \registers[182][4] , \registers[182][3] , \registers[182][2] ,
         \registers[182][1] , \registers[182][0] , \registers[181][7] ,
         \registers[181][6] , \registers[181][5] , \registers[181][4] ,
         \registers[181][3] , \registers[181][2] , \registers[181][1] ,
         \registers[181][0] , \registers[180][7] , \registers[180][6] ,
         \registers[180][5] , \registers[180][4] , \registers[180][3] ,
         \registers[180][2] , \registers[180][1] , \registers[180][0] ,
         \registers[179][7] , \registers[179][6] , \registers[179][5] ,
         \registers[179][4] , \registers[179][3] , \registers[179][2] ,
         \registers[179][1] , \registers[179][0] , \registers[178][7] ,
         \registers[178][6] , \registers[178][5] , \registers[178][4] ,
         \registers[178][3] , \registers[178][2] , \registers[178][1] ,
         \registers[178][0] , \registers[177][7] , \registers[177][6] ,
         \registers[177][5] , \registers[177][4] , \registers[177][3] ,
         \registers[177][2] , \registers[177][1] , \registers[177][0] ,
         \registers[176][7] , \registers[176][6] , \registers[176][5] ,
         \registers[176][4] , \registers[176][3] , \registers[176][2] ,
         \registers[176][1] , \registers[176][0] , \registers[175][7] ,
         \registers[175][6] , \registers[175][5] , \registers[175][4] ,
         \registers[175][3] , \registers[175][2] , \registers[175][1] ,
         \registers[175][0] , \registers[174][7] , \registers[174][6] ,
         \registers[174][5] , \registers[174][4] , \registers[174][3] ,
         \registers[174][2] , \registers[174][1] , \registers[174][0] ,
         \registers[173][7] , \registers[173][6] , \registers[173][5] ,
         \registers[173][4] , \registers[173][3] , \registers[173][2] ,
         \registers[173][1] , \registers[173][0] , \registers[172][7] ,
         \registers[172][6] , \registers[172][5] , \registers[172][4] ,
         \registers[172][3] , \registers[172][2] , \registers[172][1] ,
         \registers[172][0] , \registers[171][7] , \registers[171][6] ,
         \registers[171][5] , \registers[171][4] , \registers[171][3] ,
         \registers[171][2] , \registers[171][1] , \registers[171][0] ,
         \registers[170][7] , \registers[170][6] , \registers[170][5] ,
         \registers[170][4] , \registers[170][3] , \registers[170][2] ,
         \registers[170][1] , \registers[170][0] , \registers[169][7] ,
         \registers[169][6] , \registers[169][5] , \registers[169][4] ,
         \registers[169][3] , \registers[169][2] , \registers[169][1] ,
         \registers[169][0] , \registers[168][7] , \registers[168][6] ,
         \registers[168][5] , \registers[168][4] , \registers[168][3] ,
         \registers[168][2] , \registers[168][1] , \registers[168][0] ,
         \registers[167][7] , \registers[167][6] , \registers[167][5] ,
         \registers[167][4] , \registers[167][3] , \registers[167][2] ,
         \registers[167][1] , \registers[167][0] , \registers[166][7] ,
         \registers[166][6] , \registers[166][5] , \registers[166][4] ,
         \registers[166][3] , \registers[166][2] , \registers[166][1] ,
         \registers[166][0] , \registers[165][7] , \registers[165][6] ,
         \registers[165][5] , \registers[165][4] , \registers[165][3] ,
         \registers[165][2] , \registers[165][1] , \registers[165][0] ,
         \registers[164][7] , \registers[164][6] , \registers[164][5] ,
         \registers[164][4] , \registers[164][3] , \registers[164][2] ,
         \registers[164][1] , \registers[164][0] , \registers[163][7] ,
         \registers[163][6] , \registers[163][5] , \registers[163][4] ,
         \registers[163][3] , \registers[163][2] , \registers[163][1] ,
         \registers[163][0] , \registers[162][7] , \registers[162][6] ,
         \registers[162][5] , \registers[162][4] , \registers[162][3] ,
         \registers[162][2] , \registers[162][1] , \registers[162][0] ,
         \registers[161][7] , \registers[161][6] , \registers[161][5] ,
         \registers[161][4] , \registers[161][3] , \registers[161][2] ,
         \registers[161][1] , \registers[161][0] , \registers[160][7] ,
         \registers[160][6] , \registers[160][5] , \registers[160][4] ,
         \registers[160][3] , \registers[160][2] , \registers[160][1] ,
         \registers[160][0] , \registers[223][7] , \registers[223][6] ,
         \registers[223][5] , \registers[223][4] , \registers[223][3] ,
         \registers[223][2] , \registers[223][1] , \registers[223][0] ,
         \registers[222][7] , \registers[222][6] , \registers[222][5] ,
         \registers[222][4] , \registers[222][3] , \registers[222][2] ,
         \registers[222][1] , \registers[222][0] , \registers[221][7] ,
         \registers[221][6] , \registers[221][5] , \registers[221][4] ,
         \registers[221][3] , \registers[221][2] , \registers[221][1] ,
         \registers[221][0] , \registers[220][7] , \registers[220][6] ,
         \registers[220][5] , \registers[220][4] , \registers[220][3] ,
         \registers[220][2] , \registers[220][1] , \registers[220][0] ,
         \registers[219][7] , \registers[219][6] , \registers[219][5] ,
         \registers[219][4] , \registers[219][3] , \registers[219][2] ,
         \registers[219][1] , \registers[219][0] , \registers[218][7] ,
         \registers[218][6] , \registers[218][5] , \registers[218][4] ,
         \registers[218][3] , \registers[218][2] , \registers[218][1] ,
         \registers[218][0] , \registers[217][7] , \registers[217][6] ,
         \registers[217][5] , \registers[217][4] , \registers[217][3] ,
         \registers[217][2] , \registers[217][1] , \registers[217][0] ,
         \registers[216][7] , \registers[216][6] , \registers[216][5] ,
         \registers[216][4] , \registers[216][3] , \registers[216][2] ,
         \registers[216][1] , \registers[216][0] , \registers[215][7] ,
         \registers[215][6] , \registers[215][5] , \registers[215][4] ,
         \registers[215][3] , \registers[215][2] , \registers[215][1] ,
         \registers[215][0] , \registers[214][7] , \registers[214][6] ,
         \registers[214][5] , \registers[214][4] , \registers[214][3] ,
         \registers[214][2] , \registers[214][1] , \registers[214][0] ,
         \registers[213][7] , \registers[213][6] , \registers[213][5] ,
         \registers[213][4] , \registers[213][3] , \registers[213][2] ,
         \registers[213][1] , \registers[213][0] , \registers[212][7] ,
         \registers[212][6] , \registers[212][5] , \registers[212][4] ,
         \registers[212][3] , \registers[212][2] , \registers[212][1] ,
         \registers[212][0] , \registers[211][7] , \registers[211][6] ,
         \registers[211][5] , \registers[211][4] , \registers[211][3] ,
         \registers[211][2] , \registers[211][1] , \registers[211][0] ,
         \registers[210][7] , \registers[210][6] , \registers[210][5] ,
         \registers[210][4] , \registers[210][3] , \registers[210][2] ,
         \registers[210][1] , \registers[210][0] , \registers[209][7] ,
         \registers[209][6] , \registers[209][5] , \registers[209][4] ,
         \registers[209][3] , \registers[209][2] , \registers[209][1] ,
         \registers[209][0] , \registers[208][7] , \registers[208][6] ,
         \registers[208][5] , \registers[208][4] , \registers[208][3] ,
         \registers[208][2] , \registers[208][1] , \registers[208][0] ,
         \registers[207][7] , \registers[207][6] , \registers[207][5] ,
         \registers[207][4] , \registers[207][3] , \registers[207][2] ,
         \registers[207][1] , \registers[207][0] , \registers[206][7] ,
         \registers[206][6] , \registers[206][5] , \registers[206][4] ,
         \registers[206][3] , \registers[206][2] , \registers[206][1] ,
         \registers[206][0] , \registers[205][7] , \registers[205][6] ,
         \registers[205][5] , \registers[205][4] , \registers[205][3] ,
         \registers[205][2] , \registers[205][1] , \registers[205][0] ,
         \registers[204][7] , \registers[204][6] , \registers[204][5] ,
         \registers[204][4] , \registers[204][3] , \registers[204][2] ,
         \registers[204][1] , \registers[204][0] , \registers[203][7] ,
         \registers[203][6] , \registers[203][5] , \registers[203][4] ,
         \registers[203][3] , \registers[203][2] , \registers[203][1] ,
         \registers[203][0] , \registers[202][7] , \registers[202][6] ,
         \registers[202][5] , \registers[202][4] , \registers[202][3] ,
         \registers[202][2] , \registers[202][1] , \registers[202][0] ,
         \registers[201][7] , \registers[201][6] , \registers[201][5] ,
         \registers[201][4] , \registers[201][3] , \registers[201][2] ,
         \registers[201][1] , \registers[201][0] , \registers[200][7] ,
         \registers[200][6] , \registers[200][5] , \registers[200][4] ,
         \registers[200][3] , \registers[200][2] , \registers[200][1] ,
         \registers[200][0] , \registers[199][7] , \registers[199][6] ,
         \registers[199][5] , \registers[199][4] , \registers[199][3] ,
         \registers[199][2] , \registers[199][1] , \registers[199][0] ,
         \registers[198][7] , \registers[198][6] , \registers[198][5] ,
         \registers[198][4] , \registers[198][3] , \registers[198][2] ,
         \registers[198][1] , \registers[198][0] , \registers[197][7] ,
         \registers[197][6] , \registers[197][5] , \registers[197][4] ,
         \registers[197][3] , \registers[197][2] , \registers[197][1] ,
         \registers[197][0] , \registers[196][7] , \registers[196][6] ,
         \registers[196][5] , \registers[196][4] , \registers[196][3] ,
         \registers[196][2] , \registers[196][1] , \registers[196][0] ,
         \registers[195][7] , \registers[195][6] , \registers[195][5] ,
         \registers[195][4] , \registers[195][3] , \registers[195][2] ,
         \registers[195][1] , \registers[195][0] , \registers[194][7] ,
         \registers[194][6] , \registers[194][5] , \registers[194][4] ,
         \registers[194][3] , \registers[194][2] , \registers[194][1] ,
         \registers[194][0] , \registers[193][7] , \registers[193][6] ,
         \registers[193][5] , \registers[193][4] , \registers[193][3] ,
         \registers[193][2] , \registers[193][1] , \registers[193][0] ,
         \registers[192][7] , \registers[192][6] , \registers[192][5] ,
         \registers[192][4] , \registers[192][3] , \registers[192][2] ,
         \registers[192][1] , \registers[192][0] , \registers[255][7] ,
         \registers[255][6] , \registers[255][5] , \registers[255][4] ,
         \registers[255][3] , \registers[255][2] , \registers[255][1] ,
         \registers[255][0] , \registers[254][7] , \registers[254][6] ,
         \registers[254][5] , \registers[254][4] , \registers[254][3] ,
         \registers[254][2] , \registers[254][1] , \registers[254][0] ,
         \registers[253][7] , \registers[253][6] , \registers[253][5] ,
         \registers[253][4] , \registers[253][3] , \registers[253][2] ,
         \registers[253][1] , \registers[253][0] , \registers[252][7] ,
         \registers[252][6] , \registers[252][5] , \registers[252][4] ,
         \registers[252][3] , \registers[252][2] , \registers[252][1] ,
         \registers[252][0] , \registers[251][7] , \registers[251][6] ,
         \registers[251][5] , \registers[251][4] , \registers[251][3] ,
         \registers[251][2] , \registers[251][1] , \registers[251][0] ,
         \registers[250][7] , \registers[250][6] , \registers[250][5] ,
         \registers[250][4] , \registers[250][3] , \registers[250][2] ,
         \registers[250][1] , \registers[250][0] , \registers[249][7] ,
         \registers[249][6] , \registers[249][5] , \registers[249][4] ,
         \registers[249][3] , \registers[249][2] , \registers[249][1] ,
         \registers[249][0] , \registers[248][7] , \registers[248][6] ,
         \registers[248][5] , \registers[248][4] , \registers[248][3] ,
         \registers[248][2] , \registers[248][1] , \registers[248][0] ,
         \registers[247][7] , \registers[247][6] , \registers[247][5] ,
         \registers[247][4] , \registers[247][3] , \registers[247][2] ,
         \registers[247][1] , \registers[247][0] , \registers[246][7] ,
         \registers[246][6] , \registers[246][5] , \registers[246][4] ,
         \registers[246][3] , \registers[246][2] , \registers[246][1] ,
         \registers[246][0] , \registers[245][7] , \registers[245][6] ,
         \registers[245][5] , \registers[245][4] , \registers[245][3] ,
         \registers[245][2] , \registers[245][1] , \registers[245][0] ,
         \registers[244][7] , \registers[244][6] , \registers[244][5] ,
         \registers[244][4] , \registers[244][3] , \registers[244][2] ,
         \registers[244][1] , \registers[244][0] , \registers[243][7] ,
         \registers[243][6] , \registers[243][5] , \registers[243][4] ,
         \registers[243][3] , \registers[243][2] , \registers[243][1] ,
         \registers[243][0] , \registers[242][7] , \registers[242][6] ,
         \registers[242][5] , \registers[242][4] , \registers[242][3] ,
         \registers[242][2] , \registers[242][1] , \registers[242][0] ,
         \registers[241][7] , \registers[241][6] , \registers[241][5] ,
         \registers[241][4] , \registers[241][3] , \registers[241][2] ,
         \registers[241][1] , \registers[241][0] , \registers[240][7] ,
         \registers[240][6] , \registers[240][5] , \registers[240][4] ,
         \registers[240][3] , \registers[240][2] , \registers[240][1] ,
         \registers[240][0] , \registers[239][7] , \registers[239][6] ,
         \registers[239][5] , \registers[239][4] , \registers[239][3] ,
         \registers[239][2] , \registers[239][1] , \registers[239][0] ,
         \registers[238][7] , \registers[238][6] , \registers[238][5] ,
         \registers[238][4] , \registers[238][3] , \registers[238][2] ,
         \registers[238][1] , \registers[238][0] , \registers[237][7] ,
         \registers[237][6] , \registers[237][5] , \registers[237][4] ,
         \registers[237][3] , \registers[237][2] , \registers[237][1] ,
         \registers[237][0] , \registers[236][7] , \registers[236][6] ,
         \registers[236][5] , \registers[236][4] , \registers[236][3] ,
         \registers[236][2] , \registers[236][1] , \registers[236][0] ,
         \registers[235][7] , \registers[235][6] , \registers[235][5] ,
         \registers[235][4] , \registers[235][3] , \registers[235][2] ,
         \registers[235][1] , \registers[235][0] , \registers[234][7] ,
         \registers[234][6] , \registers[234][5] , \registers[234][4] ,
         \registers[234][3] , \registers[234][2] , \registers[234][1] ,
         \registers[234][0] , \registers[233][7] , \registers[233][6] ,
         \registers[233][5] , \registers[233][4] , \registers[233][3] ,
         \registers[233][2] , \registers[233][1] , \registers[233][0] ,
         \registers[232][7] , \registers[232][6] , \registers[232][5] ,
         \registers[232][4] , \registers[232][3] , \registers[232][2] ,
         \registers[232][1] , \registers[232][0] , \registers[231][7] ,
         \registers[231][6] , \registers[231][5] , \registers[231][4] ,
         \registers[231][3] , \registers[231][2] , \registers[231][1] ,
         \registers[231][0] , \registers[230][7] , \registers[230][6] ,
         \registers[230][5] , \registers[230][4] , \registers[230][3] ,
         \registers[230][2] , \registers[230][1] , \registers[230][0] ,
         \registers[229][7] , \registers[229][6] , \registers[229][5] ,
         \registers[229][4] , \registers[229][3] , \registers[229][2] ,
         \registers[229][1] , \registers[229][0] , \registers[228][7] ,
         \registers[228][6] , \registers[228][5] , \registers[228][4] ,
         \registers[228][3] , \registers[228][2] , \registers[228][1] ,
         \registers[228][0] , \registers[227][7] , \registers[227][6] ,
         \registers[227][5] , \registers[227][4] , \registers[227][3] ,
         \registers[227][2] , \registers[227][1] , \registers[227][0] ,
         \registers[226][7] , \registers[226][6] , \registers[226][5] ,
         \registers[226][4] , \registers[226][3] , \registers[226][2] ,
         \registers[226][1] , \registers[226][0] , \registers[225][7] ,
         \registers[225][6] , \registers[225][5] , \registers[225][4] ,
         \registers[225][3] , \registers[225][2] , \registers[225][1] ,
         \registers[225][0] , \registers[224][7] , \registers[224][6] ,
         \registers[224][5] , \registers[224][4] , \registers[224][3] ,
         \registers[224][2] , \registers[224][1] , \registers[224][0] ,
         \registers[287][7] , \registers[287][6] , \registers[287][5] ,
         \registers[287][4] , \registers[287][3] , \registers[287][2] ,
         \registers[287][1] , \registers[287][0] , \registers[286][7] ,
         \registers[286][6] , \registers[286][5] , \registers[286][4] ,
         \registers[286][3] , \registers[286][2] , \registers[286][1] ,
         \registers[286][0] , \registers[285][7] , \registers[285][6] ,
         \registers[285][5] , \registers[285][4] , \registers[285][3] ,
         \registers[285][2] , \registers[285][1] , \registers[285][0] ,
         \registers[284][7] , \registers[284][6] , \registers[284][5] ,
         \registers[284][4] , \registers[284][3] , \registers[284][2] ,
         \registers[284][1] , \registers[284][0] , \registers[283][7] ,
         \registers[283][6] , \registers[283][5] , \registers[283][4] ,
         \registers[283][3] , \registers[283][2] , \registers[283][1] ,
         \registers[283][0] , \registers[282][7] , \registers[282][6] ,
         \registers[282][5] , \registers[282][4] , \registers[282][3] ,
         \registers[282][2] , \registers[282][1] , \registers[282][0] ,
         \registers[281][7] , \registers[281][6] , \registers[281][5] ,
         \registers[281][4] , \registers[281][3] , \registers[281][2] ,
         \registers[281][1] , \registers[281][0] , \registers[280][7] ,
         \registers[280][6] , \registers[280][5] , \registers[280][4] ,
         \registers[280][3] , \registers[280][2] , \registers[280][1] ,
         \registers[280][0] , \registers[279][7] , \registers[279][6] ,
         \registers[279][5] , \registers[279][4] , \registers[279][3] ,
         \registers[279][2] , \registers[279][1] , \registers[279][0] ,
         \registers[278][7] , \registers[278][6] , \registers[278][5] ,
         \registers[278][4] , \registers[278][3] , \registers[278][2] ,
         \registers[278][1] , \registers[278][0] , \registers[277][7] ,
         \registers[277][6] , \registers[277][5] , \registers[277][4] ,
         \registers[277][3] , \registers[277][2] , \registers[277][1] ,
         \registers[277][0] , \registers[276][7] , \registers[276][6] ,
         \registers[276][5] , \registers[276][4] , \registers[276][3] ,
         \registers[276][2] , \registers[276][1] , \registers[276][0] ,
         \registers[275][7] , \registers[275][6] , \registers[275][5] ,
         \registers[275][4] , \registers[275][3] , \registers[275][2] ,
         \registers[275][1] , \registers[275][0] , \registers[274][7] ,
         \registers[274][6] , \registers[274][5] , \registers[274][4] ,
         \registers[274][3] , \registers[274][2] , \registers[274][1] ,
         \registers[274][0] , \registers[273][7] , \registers[273][6] ,
         \registers[273][5] , \registers[273][4] , \registers[273][3] ,
         \registers[273][2] , \registers[273][1] , \registers[273][0] ,
         \registers[272][7] , \registers[272][6] , \registers[272][5] ,
         \registers[272][4] , \registers[272][3] , \registers[272][2] ,
         \registers[272][1] , \registers[272][0] , \registers[271][7] ,
         \registers[271][6] , \registers[271][5] , \registers[271][4] ,
         \registers[271][3] , \registers[271][2] , \registers[271][1] ,
         \registers[271][0] , \registers[270][7] , \registers[270][6] ,
         \registers[270][5] , \registers[270][4] , \registers[270][3] ,
         \registers[270][2] , \registers[270][1] , \registers[270][0] ,
         \registers[269][7] , \registers[269][6] , \registers[269][5] ,
         \registers[269][4] , \registers[269][3] , \registers[269][2] ,
         \registers[269][1] , \registers[269][0] , \registers[268][7] ,
         \registers[268][6] , \registers[268][5] , \registers[268][4] ,
         \registers[268][3] , \registers[268][2] , \registers[268][1] ,
         \registers[268][0] , \registers[267][7] , \registers[267][6] ,
         \registers[267][5] , \registers[267][4] , \registers[267][3] ,
         \registers[267][2] , \registers[267][1] , \registers[267][0] ,
         \registers[266][7] , \registers[266][6] , \registers[266][5] ,
         \registers[266][4] , \registers[266][3] , \registers[266][2] ,
         \registers[266][1] , \registers[266][0] , \registers[265][7] ,
         \registers[265][6] , \registers[265][5] , \registers[265][4] ,
         \registers[265][3] , \registers[265][2] , \registers[265][1] ,
         \registers[265][0] , \registers[264][7] , \registers[264][6] ,
         \registers[264][5] , \registers[264][4] , \registers[264][3] ,
         \registers[264][2] , \registers[264][1] , \registers[264][0] ,
         \registers[263][7] , \registers[263][6] , \registers[263][5] ,
         \registers[263][4] , \registers[263][3] , \registers[263][2] ,
         \registers[263][1] , \registers[263][0] , \registers[262][7] ,
         \registers[262][6] , \registers[262][5] , \registers[262][4] ,
         \registers[262][3] , \registers[262][2] , \registers[262][1] ,
         \registers[262][0] , \registers[261][7] , \registers[261][6] ,
         \registers[261][5] , \registers[261][4] , \registers[261][3] ,
         \registers[261][2] , \registers[261][1] , \registers[261][0] ,
         \registers[260][7] , \registers[260][6] , \registers[260][5] ,
         \registers[260][4] , \registers[260][3] , \registers[260][2] ,
         \registers[260][1] , \registers[260][0] , \registers[259][7] ,
         \registers[259][6] , \registers[259][5] , \registers[259][4] ,
         \registers[259][3] , \registers[259][2] , \registers[259][1] ,
         \registers[259][0] , \registers[258][7] , \registers[258][6] ,
         \registers[258][5] , \registers[258][4] , \registers[258][3] ,
         \registers[258][2] , \registers[258][1] , \registers[258][0] ,
         \registers[257][7] , \registers[257][6] , \registers[257][5] ,
         \registers[257][4] , \registers[257][3] , \registers[257][2] ,
         \registers[257][1] , \registers[257][0] , \registers[256][7] ,
         \registers[256][6] , \registers[256][5] , \registers[256][4] ,
         \registers[256][3] , \registers[256][2] , \registers[256][1] ,
         \registers[256][0] , \registers[319][7] , \registers[319][6] ,
         \registers[319][5] , \registers[319][4] , \registers[319][3] ,
         \registers[319][2] , \registers[319][1] , \registers[319][0] ,
         \registers[318][7] , \registers[318][6] , \registers[318][5] ,
         \registers[318][4] , \registers[318][3] , \registers[318][2] ,
         \registers[318][1] , \registers[318][0] , \registers[317][7] ,
         \registers[317][6] , \registers[317][5] , \registers[317][4] ,
         \registers[317][3] , \registers[317][2] , \registers[317][1] ,
         \registers[317][0] , \registers[316][7] , \registers[316][6] ,
         \registers[316][5] , \registers[316][4] , \registers[316][3] ,
         \registers[316][2] , \registers[316][1] , \registers[316][0] ,
         \registers[315][7] , \registers[315][6] , \registers[315][5] ,
         \registers[315][4] , \registers[315][3] , \registers[315][2] ,
         \registers[315][1] , \registers[315][0] , \registers[314][7] ,
         \registers[314][6] , \registers[314][5] , \registers[314][4] ,
         \registers[314][3] , \registers[314][2] , \registers[314][1] ,
         \registers[314][0] , \registers[313][7] , \registers[313][6] ,
         \registers[313][5] , \registers[313][4] , \registers[313][3] ,
         \registers[313][2] , \registers[313][1] , \registers[313][0] ,
         \registers[312][7] , \registers[312][6] , \registers[312][5] ,
         \registers[312][4] , \registers[312][3] , \registers[312][2] ,
         \registers[312][1] , \registers[312][0] , \registers[311][7] ,
         \registers[311][6] , \registers[311][5] , \registers[311][4] ,
         \registers[311][3] , \registers[311][2] , \registers[311][1] ,
         \registers[311][0] , \registers[310][7] , \registers[310][6] ,
         \registers[310][5] , \registers[310][4] , \registers[310][3] ,
         \registers[310][2] , \registers[310][1] , \registers[310][0] ,
         \registers[309][7] , \registers[309][6] , \registers[309][5] ,
         \registers[309][4] , \registers[309][3] , \registers[309][2] ,
         \registers[309][1] , \registers[309][0] , \registers[308][7] ,
         \registers[308][6] , \registers[308][5] , \registers[308][4] ,
         \registers[308][3] , \registers[308][2] , \registers[308][1] ,
         \registers[308][0] , \registers[307][7] , \registers[307][6] ,
         \registers[307][5] , \registers[307][4] , \registers[307][3] ,
         \registers[307][2] , \registers[307][1] , \registers[307][0] ,
         \registers[306][7] , \registers[306][6] , \registers[306][5] ,
         \registers[306][4] , \registers[306][3] , \registers[306][2] ,
         \registers[306][1] , \registers[306][0] , \registers[305][7] ,
         \registers[305][6] , \registers[305][5] , \registers[305][4] ,
         \registers[305][3] , \registers[305][2] , \registers[305][1] ,
         \registers[305][0] , \registers[304][7] , \registers[304][6] ,
         \registers[304][5] , \registers[304][4] , \registers[304][3] ,
         \registers[304][2] , \registers[304][1] , \registers[304][0] ,
         \registers[303][7] , \registers[303][6] , \registers[303][5] ,
         \registers[303][4] , \registers[303][3] , \registers[303][2] ,
         \registers[303][1] , \registers[303][0] , \registers[302][7] ,
         \registers[302][6] , \registers[302][5] , \registers[302][4] ,
         \registers[302][3] , \registers[302][2] , \registers[302][1] ,
         \registers[302][0] , \registers[301][7] , \registers[301][6] ,
         \registers[301][5] , \registers[301][4] , \registers[301][3] ,
         \registers[301][2] , \registers[301][1] , \registers[301][0] ,
         \registers[300][7] , \registers[300][6] , \registers[300][5] ,
         \registers[300][4] , \registers[300][3] , \registers[300][2] ,
         \registers[300][1] , \registers[300][0] , \registers[299][7] ,
         \registers[299][6] , \registers[299][5] , \registers[299][4] ,
         \registers[299][3] , \registers[299][2] , \registers[299][1] ,
         \registers[299][0] , \registers[298][7] , \registers[298][6] ,
         \registers[298][5] , \registers[298][4] , \registers[298][3] ,
         \registers[298][2] , \registers[298][1] , \registers[298][0] ,
         \registers[297][7] , \registers[297][6] , \registers[297][5] ,
         \registers[297][4] , \registers[297][3] , \registers[297][2] ,
         \registers[297][1] , \registers[297][0] , \registers[296][7] ,
         \registers[296][6] , \registers[296][5] , \registers[296][4] ,
         \registers[296][3] , \registers[296][2] , \registers[296][1] ,
         \registers[296][0] , \registers[295][7] , \registers[295][6] ,
         \registers[295][5] , \registers[295][4] , \registers[295][3] ,
         \registers[295][2] , \registers[295][1] , \registers[295][0] ,
         \registers[294][7] , \registers[294][6] , \registers[294][5] ,
         \registers[294][4] , \registers[294][3] , \registers[294][2] ,
         \registers[294][1] , \registers[294][0] , \registers[293][7] ,
         \registers[293][6] , \registers[293][5] , \registers[293][4] ,
         \registers[293][3] , \registers[293][2] , \registers[293][1] ,
         \registers[293][0] , \registers[292][7] , \registers[292][6] ,
         \registers[292][5] , \registers[292][4] , \registers[292][3] ,
         \registers[292][2] , \registers[292][1] , \registers[292][0] ,
         \registers[291][7] , \registers[291][6] , \registers[291][5] ,
         \registers[291][4] , \registers[291][3] , \registers[291][2] ,
         \registers[291][1] , \registers[291][0] , \registers[290][7] ,
         \registers[290][6] , \registers[290][5] , \registers[290][4] ,
         \registers[290][3] , \registers[290][2] , \registers[290][1] ,
         \registers[290][0] , \registers[289][7] , \registers[289][6] ,
         \registers[289][5] , \registers[289][4] , \registers[289][3] ,
         \registers[289][2] , \registers[289][1] , \registers[289][0] ,
         \registers[288][7] , \registers[288][6] , \registers[288][5] ,
         \registers[288][4] , \registers[288][3] , \registers[288][2] ,
         \registers[288][1] , \registers[288][0] , \registers[351][7] ,
         \registers[351][6] , \registers[351][5] , \registers[351][4] ,
         \registers[351][3] , \registers[351][2] , \registers[351][1] ,
         \registers[351][0] , \registers[350][7] , \registers[350][6] ,
         \registers[350][5] , \registers[350][4] , \registers[350][3] ,
         \registers[350][2] , \registers[350][1] , \registers[350][0] ,
         \registers[349][7] , \registers[349][6] , \registers[349][5] ,
         \registers[349][4] , \registers[349][3] , \registers[349][2] ,
         \registers[349][1] , \registers[349][0] , \registers[348][7] ,
         \registers[348][6] , \registers[348][5] , \registers[348][4] ,
         \registers[348][3] , \registers[348][2] , \registers[348][1] ,
         \registers[348][0] , \registers[347][7] , \registers[347][6] ,
         \registers[347][5] , \registers[347][4] , \registers[347][3] ,
         \registers[347][2] , \registers[347][1] , \registers[347][0] ,
         \registers[346][7] , \registers[346][6] , \registers[346][5] ,
         \registers[346][4] , \registers[346][3] , \registers[346][2] ,
         \registers[346][1] , \registers[346][0] , \registers[345][7] ,
         \registers[345][6] , \registers[345][5] , \registers[345][4] ,
         \registers[345][3] , \registers[345][2] , \registers[345][1] ,
         \registers[345][0] , \registers[344][7] , \registers[344][6] ,
         \registers[344][5] , \registers[344][4] , \registers[344][3] ,
         \registers[344][2] , \registers[344][1] , \registers[344][0] ,
         \registers[343][7] , \registers[343][6] , \registers[343][5] ,
         \registers[343][4] , \registers[343][3] , \registers[343][2] ,
         \registers[343][1] , \registers[343][0] , \registers[342][7] ,
         \registers[342][6] , \registers[342][5] , \registers[342][4] ,
         \registers[342][3] , \registers[342][2] , \registers[342][1] ,
         \registers[342][0] , \registers[341][7] , \registers[341][6] ,
         \registers[341][5] , \registers[341][4] , \registers[341][3] ,
         \registers[341][2] , \registers[341][1] , \registers[341][0] ,
         \registers[340][7] , \registers[340][6] , \registers[340][5] ,
         \registers[340][4] , \registers[340][3] , \registers[340][2] ,
         \registers[340][1] , \registers[340][0] , \registers[339][7] ,
         \registers[339][6] , \registers[339][5] , \registers[339][4] ,
         \registers[339][3] , \registers[339][2] , \registers[339][1] ,
         \registers[339][0] , \registers[338][7] , \registers[338][6] ,
         \registers[338][5] , \registers[338][4] , \registers[338][3] ,
         \registers[338][2] , \registers[338][1] , \registers[338][0] ,
         \registers[337][7] , \registers[337][6] , \registers[337][5] ,
         \registers[337][4] , \registers[337][3] , \registers[337][2] ,
         \registers[337][1] , \registers[337][0] , \registers[336][7] ,
         \registers[336][6] , \registers[336][5] , \registers[336][4] ,
         \registers[336][3] , \registers[336][2] , \registers[336][1] ,
         \registers[336][0] , \registers[335][7] , \registers[335][6] ,
         \registers[335][5] , \registers[335][4] , \registers[335][3] ,
         \registers[335][2] , \registers[335][1] , \registers[335][0] ,
         \registers[334][7] , \registers[334][6] , \registers[334][5] ,
         \registers[334][4] , \registers[334][3] , \registers[334][2] ,
         \registers[334][1] , \registers[334][0] , \registers[333][7] ,
         \registers[333][6] , \registers[333][5] , \registers[333][4] ,
         \registers[333][3] , \registers[333][2] , \registers[333][1] ,
         \registers[333][0] , \registers[332][7] , \registers[332][6] ,
         \registers[332][5] , \registers[332][4] , \registers[332][3] ,
         \registers[332][2] , \registers[332][1] , \registers[332][0] ,
         \registers[331][7] , \registers[331][6] , \registers[331][5] ,
         \registers[331][4] , \registers[331][3] , \registers[331][2] ,
         \registers[331][1] , \registers[331][0] , \registers[330][7] ,
         \registers[330][6] , \registers[330][5] , \registers[330][4] ,
         \registers[330][3] , \registers[330][2] , \registers[330][1] ,
         \registers[330][0] , \registers[329][7] , \registers[329][6] ,
         \registers[329][5] , \registers[329][4] , \registers[329][3] ,
         \registers[329][2] , \registers[329][1] , \registers[329][0] ,
         \registers[328][7] , \registers[328][6] , \registers[328][5] ,
         \registers[328][4] , \registers[328][3] , \registers[328][2] ,
         \registers[328][1] , \registers[328][0] , \registers[327][7] ,
         \registers[327][6] , \registers[327][5] , \registers[327][4] ,
         \registers[327][3] , \registers[327][2] , \registers[327][1] ,
         \registers[327][0] , \registers[326][7] , \registers[326][6] ,
         \registers[326][5] , \registers[326][4] , \registers[326][3] ,
         \registers[326][2] , \registers[326][1] , \registers[326][0] ,
         \registers[325][7] , \registers[325][6] , \registers[325][5] ,
         \registers[325][4] , \registers[325][3] , \registers[325][2] ,
         \registers[325][1] , \registers[325][0] , \registers[324][7] ,
         \registers[324][6] , \registers[324][5] , \registers[324][4] ,
         \registers[324][3] , \registers[324][2] , \registers[324][1] ,
         \registers[324][0] , \registers[323][7] , \registers[323][6] ,
         \registers[323][5] , \registers[323][4] , \registers[323][3] ,
         \registers[323][2] , \registers[323][1] , \registers[323][0] ,
         \registers[322][7] , \registers[322][6] , \registers[322][5] ,
         \registers[322][4] , \registers[322][3] , \registers[322][2] ,
         \registers[322][1] , \registers[322][0] , \registers[321][7] ,
         \registers[321][6] , \registers[321][5] , \registers[321][4] ,
         \registers[321][3] , \registers[321][2] , \registers[321][1] ,
         \registers[321][0] , \registers[320][7] , \registers[320][6] ,
         \registers[320][5] , \registers[320][4] , \registers[320][3] ,
         \registers[320][2] , \registers[320][1] , \registers[320][0] ,
         \registers[383][7] , \registers[383][6] , \registers[383][5] ,
         \registers[383][4] , \registers[383][3] , \registers[383][2] ,
         \registers[383][1] , \registers[383][0] , \registers[382][7] ,
         \registers[382][6] , \registers[382][5] , \registers[382][4] ,
         \registers[382][3] , \registers[382][2] , \registers[382][1] ,
         \registers[382][0] , \registers[381][7] , \registers[381][6] ,
         \registers[381][5] , \registers[381][4] , \registers[381][3] ,
         \registers[381][2] , \registers[381][1] , \registers[381][0] ,
         \registers[380][7] , \registers[380][6] , \registers[380][5] ,
         \registers[380][4] , \registers[380][3] , \registers[380][2] ,
         \registers[380][1] , \registers[380][0] , \registers[379][7] ,
         \registers[379][6] , \registers[379][5] , \registers[379][4] ,
         \registers[379][3] , \registers[379][2] , \registers[379][1] ,
         \registers[379][0] , \registers[378][7] , \registers[378][6] ,
         \registers[378][5] , \registers[378][4] , \registers[378][3] ,
         \registers[378][2] , \registers[378][1] , \registers[378][0] ,
         \registers[377][7] , \registers[377][6] , \registers[377][5] ,
         \registers[377][4] , \registers[377][3] , \registers[377][2] ,
         \registers[377][1] , \registers[377][0] , \registers[376][7] ,
         \registers[376][6] , \registers[376][5] , \registers[376][4] ,
         \registers[376][3] , \registers[376][2] , \registers[376][1] ,
         \registers[376][0] , \registers[375][7] , \registers[375][6] ,
         \registers[375][5] , \registers[375][4] , \registers[375][3] ,
         \registers[375][2] , \registers[375][1] , \registers[375][0] ,
         \registers[374][7] , \registers[374][6] , \registers[374][5] ,
         \registers[374][4] , \registers[374][3] , \registers[374][2] ,
         \registers[374][1] , \registers[374][0] , \registers[373][7] ,
         \registers[373][6] , \registers[373][5] , \registers[373][4] ,
         \registers[373][3] , \registers[373][2] , \registers[373][1] ,
         \registers[373][0] , \registers[372][7] , \registers[372][6] ,
         \registers[372][5] , \registers[372][4] , \registers[372][3] ,
         \registers[372][2] , \registers[372][1] , \registers[372][0] ,
         \registers[371][7] , \registers[371][6] , \registers[371][5] ,
         \registers[371][4] , \registers[371][3] , \registers[371][2] ,
         \registers[371][1] , \registers[371][0] , \registers[370][7] ,
         \registers[370][6] , \registers[370][5] , \registers[370][4] ,
         \registers[370][3] , \registers[370][2] , \registers[370][1] ,
         \registers[370][0] , \registers[369][7] , \registers[369][6] ,
         \registers[369][5] , \registers[369][4] , \registers[369][3] ,
         \registers[369][2] , \registers[369][1] , \registers[369][0] ,
         \registers[368][7] , \registers[368][6] , \registers[368][5] ,
         \registers[368][4] , \registers[368][3] , \registers[368][2] ,
         \registers[368][1] , \registers[368][0] , \registers[367][7] ,
         \registers[367][6] , \registers[367][5] , \registers[367][4] ,
         \registers[367][3] , \registers[367][2] , \registers[367][1] ,
         \registers[367][0] , \registers[366][7] , \registers[366][6] ,
         \registers[366][5] , \registers[366][4] , \registers[366][3] ,
         \registers[366][2] , \registers[366][1] , \registers[366][0] ,
         \registers[365][7] , \registers[365][6] , \registers[365][5] ,
         \registers[365][4] , \registers[365][3] , \registers[365][2] ,
         \registers[365][1] , \registers[365][0] , \registers[364][7] ,
         \registers[364][6] , \registers[364][5] , \registers[364][4] ,
         \registers[364][3] , \registers[364][2] , \registers[364][1] ,
         \registers[364][0] , \registers[363][7] , \registers[363][6] ,
         \registers[363][5] , \registers[363][4] , \registers[363][3] ,
         \registers[363][2] , \registers[363][1] , \registers[363][0] ,
         \registers[362][7] , \registers[362][6] , \registers[362][5] ,
         \registers[362][4] , \registers[362][3] , \registers[362][2] ,
         \registers[362][1] , \registers[362][0] , \registers[361][7] ,
         \registers[361][6] , \registers[361][5] , \registers[361][4] ,
         \registers[361][3] , \registers[361][2] , \registers[361][1] ,
         \registers[361][0] , \registers[360][7] , \registers[360][6] ,
         \registers[360][5] , \registers[360][4] , \registers[360][3] ,
         \registers[360][2] , \registers[360][1] , \registers[360][0] ,
         \registers[359][7] , \registers[359][6] , \registers[359][5] ,
         \registers[359][4] , \registers[359][3] , \registers[359][2] ,
         \registers[359][1] , \registers[359][0] , \registers[358][7] ,
         \registers[358][6] , \registers[358][5] , \registers[358][4] ,
         \registers[358][3] , \registers[358][2] , \registers[358][1] ,
         \registers[358][0] , \registers[357][7] , \registers[357][6] ,
         \registers[357][5] , \registers[357][4] , \registers[357][3] ,
         \registers[357][2] , \registers[357][1] , \registers[357][0] ,
         \registers[356][7] , \registers[356][6] , \registers[356][5] ,
         \registers[356][4] , \registers[356][3] , \registers[356][2] ,
         \registers[356][1] , \registers[356][0] , \registers[355][7] ,
         \registers[355][6] , \registers[355][5] , \registers[355][4] ,
         \registers[355][3] , \registers[355][2] , \registers[355][1] ,
         \registers[355][0] , \registers[354][7] , \registers[354][6] ,
         \registers[354][5] , \registers[354][4] , \registers[354][3] ,
         \registers[354][2] , \registers[354][1] , \registers[354][0] ,
         \registers[353][7] , \registers[353][6] , \registers[353][5] ,
         \registers[353][4] , \registers[353][3] , \registers[353][2] ,
         \registers[353][1] , \registers[353][0] , \registers[352][7] ,
         \registers[352][6] , \registers[352][5] , \registers[352][4] ,
         \registers[352][3] , \registers[352][2] , \registers[352][1] ,
         \registers[352][0] , \registers[415][7] , \registers[415][6] ,
         \registers[415][5] , \registers[415][4] , \registers[415][3] ,
         \registers[415][2] , \registers[415][1] , \registers[415][0] ,
         \registers[414][7] , \registers[414][6] , \registers[414][5] ,
         \registers[414][4] , \registers[414][3] , \registers[414][2] ,
         \registers[414][1] , \registers[414][0] , \registers[413][7] ,
         \registers[413][6] , \registers[413][5] , \registers[413][4] ,
         \registers[413][3] , \registers[413][2] , \registers[413][1] ,
         \registers[413][0] , \registers[412][7] , \registers[412][6] ,
         \registers[412][5] , \registers[412][4] , \registers[412][3] ,
         \registers[412][2] , \registers[412][1] , \registers[412][0] ,
         \registers[411][7] , \registers[411][6] , \registers[411][5] ,
         \registers[411][4] , \registers[411][3] , \registers[411][2] ,
         \registers[411][1] , \registers[411][0] , \registers[410][7] ,
         \registers[410][6] , \registers[410][5] , \registers[410][4] ,
         \registers[410][3] , \registers[410][2] , \registers[410][1] ,
         \registers[410][0] , \registers[409][7] , \registers[409][6] ,
         \registers[409][5] , \registers[409][4] , \registers[409][3] ,
         \registers[409][2] , \registers[409][1] , \registers[409][0] ,
         \registers[408][7] , \registers[408][6] , \registers[408][5] ,
         \registers[408][4] , \registers[408][3] , \registers[408][2] ,
         \registers[408][1] , \registers[408][0] , \registers[407][7] ,
         \registers[407][6] , \registers[407][5] , \registers[407][4] ,
         \registers[407][3] , \registers[407][2] , \registers[407][1] ,
         \registers[407][0] , \registers[406][7] , \registers[406][6] ,
         \registers[406][5] , \registers[406][4] , \registers[406][3] ,
         \registers[406][2] , \registers[406][1] , \registers[406][0] ,
         \registers[405][7] , \registers[405][6] , \registers[405][5] ,
         \registers[405][4] , \registers[405][3] , \registers[405][2] ,
         \registers[405][1] , \registers[405][0] , \registers[404][7] ,
         \registers[404][6] , \registers[404][5] , \registers[404][4] ,
         \registers[404][3] , \registers[404][2] , \registers[404][1] ,
         \registers[404][0] , \registers[403][7] , \registers[403][6] ,
         \registers[403][5] , \registers[403][4] , \registers[403][3] ,
         \registers[403][2] , \registers[403][1] , \registers[403][0] ,
         \registers[402][7] , \registers[402][6] , \registers[402][5] ,
         \registers[402][4] , \registers[402][3] , \registers[402][2] ,
         \registers[402][1] , \registers[402][0] , \registers[401][7] ,
         \registers[401][6] , \registers[401][5] , \registers[401][4] ,
         \registers[401][3] , \registers[401][2] , \registers[401][1] ,
         \registers[401][0] , \registers[400][7] , \registers[400][6] ,
         \registers[400][5] , \registers[400][4] , \registers[400][3] ,
         \registers[400][2] , \registers[400][1] , \registers[400][0] ,
         \registers[399][7] , \registers[399][6] , \registers[399][5] ,
         \registers[399][4] , \registers[399][3] , \registers[399][2] ,
         \registers[399][1] , \registers[399][0] , \registers[398][7] ,
         \registers[398][6] , \registers[398][5] , \registers[398][4] ,
         \registers[398][3] , \registers[398][2] , \registers[398][1] ,
         \registers[398][0] , \registers[397][7] , \registers[397][6] ,
         \registers[397][5] , \registers[397][4] , \registers[397][3] ,
         \registers[397][2] , \registers[397][1] , \registers[397][0] ,
         \registers[396][7] , \registers[396][6] , \registers[396][5] ,
         \registers[396][4] , \registers[396][3] , \registers[396][2] ,
         \registers[396][1] , \registers[396][0] , \registers[395][7] ,
         \registers[395][6] , \registers[395][5] , \registers[395][4] ,
         \registers[395][3] , \registers[395][2] , \registers[395][1] ,
         \registers[395][0] , \registers[394][7] , \registers[394][6] ,
         \registers[394][5] , \registers[394][4] , \registers[394][3] ,
         \registers[394][2] , \registers[394][1] , \registers[394][0] ,
         \registers[393][7] , \registers[393][6] , \registers[393][5] ,
         \registers[393][4] , \registers[393][3] , \registers[393][2] ,
         \registers[393][1] , \registers[393][0] , \registers[392][7] ,
         \registers[392][6] , \registers[392][5] , \registers[392][4] ,
         \registers[392][3] , \registers[392][2] , \registers[392][1] ,
         \registers[392][0] , \registers[391][7] , \registers[391][6] ,
         \registers[391][5] , \registers[391][4] , \registers[391][3] ,
         \registers[391][2] , \registers[391][1] , \registers[391][0] ,
         \registers[390][7] , \registers[390][6] , \registers[390][5] ,
         \registers[390][4] , \registers[390][3] , \registers[390][2] ,
         \registers[390][1] , \registers[390][0] , \registers[389][7] ,
         \registers[389][6] , \registers[389][5] , \registers[389][4] ,
         \registers[389][3] , \registers[389][2] , \registers[389][1] ,
         \registers[389][0] , \registers[388][7] , \registers[388][6] ,
         \registers[388][5] , \registers[388][4] , \registers[388][3] ,
         \registers[388][2] , \registers[388][1] , \registers[388][0] ,
         \registers[387][7] , \registers[387][6] , \registers[387][5] ,
         \registers[387][4] , \registers[387][3] , \registers[387][2] ,
         \registers[387][1] , \registers[387][0] , \registers[386][7] ,
         \registers[386][6] , \registers[386][5] , \registers[386][4] ,
         \registers[386][3] , \registers[386][2] , \registers[386][1] ,
         \registers[386][0] , \registers[385][7] , \registers[385][6] ,
         \registers[385][5] , \registers[385][4] , \registers[385][3] ,
         \registers[385][2] , \registers[385][1] , \registers[385][0] ,
         \registers[384][7] , \registers[384][6] , \registers[384][5] ,
         \registers[384][4] , \registers[384][3] , \registers[384][2] ,
         \registers[384][1] , \registers[384][0] , \registers[447][7] ,
         \registers[447][6] , \registers[447][5] , \registers[447][4] ,
         \registers[447][3] , \registers[447][2] , \registers[447][1] ,
         \registers[447][0] , \registers[446][7] , \registers[446][6] ,
         \registers[446][5] , \registers[446][4] , \registers[446][3] ,
         \registers[446][2] , \registers[446][1] , \registers[446][0] ,
         \registers[445][7] , \registers[445][6] , \registers[445][5] ,
         \registers[445][4] , \registers[445][3] , \registers[445][2] ,
         \registers[445][1] , \registers[445][0] , \registers[444][7] ,
         \registers[444][6] , \registers[444][5] , \registers[444][4] ,
         \registers[444][3] , \registers[444][2] , \registers[444][1] ,
         \registers[444][0] , \registers[443][7] , \registers[443][6] ,
         \registers[443][5] , \registers[443][4] , \registers[443][3] ,
         \registers[443][2] , \registers[443][1] , \registers[443][0] ,
         \registers[442][7] , \registers[442][6] , \registers[442][5] ,
         \registers[442][4] , \registers[442][3] , \registers[442][2] ,
         \registers[442][1] , \registers[442][0] , \registers[441][7] ,
         \registers[441][6] , \registers[441][5] , \registers[441][4] ,
         \registers[441][3] , \registers[441][2] , \registers[441][1] ,
         \registers[441][0] , \registers[440][7] , \registers[440][6] ,
         \registers[440][5] , \registers[440][4] , \registers[440][3] ,
         \registers[440][2] , \registers[440][1] , \registers[440][0] ,
         \registers[439][7] , \registers[439][6] , \registers[439][5] ,
         \registers[439][4] , \registers[439][3] , \registers[439][2] ,
         \registers[439][1] , \registers[439][0] , \registers[438][7] ,
         \registers[438][6] , \registers[438][5] , \registers[438][4] ,
         \registers[438][3] , \registers[438][2] , \registers[438][1] ,
         \registers[438][0] , \registers[437][7] , \registers[437][6] ,
         \registers[437][5] , \registers[437][4] , \registers[437][3] ,
         \registers[437][2] , \registers[437][1] , \registers[437][0] ,
         \registers[436][7] , \registers[436][6] , \registers[436][5] ,
         \registers[436][4] , \registers[436][3] , \registers[436][2] ,
         \registers[436][1] , \registers[436][0] , \registers[435][7] ,
         \registers[435][6] , \registers[435][5] , \registers[435][4] ,
         \registers[435][3] , \registers[435][2] , \registers[435][1] ,
         \registers[435][0] , \registers[434][7] , \registers[434][6] ,
         \registers[434][5] , \registers[434][4] , \registers[434][3] ,
         \registers[434][2] , \registers[434][1] , \registers[434][0] ,
         \registers[433][7] , \registers[433][6] , \registers[433][5] ,
         \registers[433][4] , \registers[433][3] , \registers[433][2] ,
         \registers[433][1] , \registers[433][0] , \registers[432][7] ,
         \registers[432][6] , \registers[432][5] , \registers[432][4] ,
         \registers[432][3] , \registers[432][2] , \registers[432][1] ,
         \registers[432][0] , \registers[431][7] , \registers[431][6] ,
         \registers[431][5] , \registers[431][4] , \registers[431][3] ,
         \registers[431][2] , \registers[431][1] , \registers[431][0] ,
         \registers[430][7] , \registers[430][6] , \registers[430][5] ,
         \registers[430][4] , \registers[430][3] , \registers[430][2] ,
         \registers[430][1] , \registers[430][0] , \registers[429][7] ,
         \registers[429][6] , \registers[429][5] , \registers[429][4] ,
         \registers[429][3] , \registers[429][2] , \registers[429][1] ,
         \registers[429][0] , \registers[428][7] , \registers[428][6] ,
         \registers[428][5] , \registers[428][4] , \registers[428][3] ,
         \registers[428][2] , \registers[428][1] , \registers[428][0] ,
         \registers[427][7] , \registers[427][6] , \registers[427][5] ,
         \registers[427][4] , \registers[427][3] , \registers[427][2] ,
         \registers[427][1] , \registers[427][0] , \registers[426][7] ,
         \registers[426][6] , \registers[426][5] , \registers[426][4] ,
         \registers[426][3] , \registers[426][2] , \registers[426][1] ,
         \registers[426][0] , \registers[425][7] , \registers[425][6] ,
         \registers[425][5] , \registers[425][4] , \registers[425][3] ,
         \registers[425][2] , \registers[425][1] , \registers[425][0] ,
         \registers[424][7] , \registers[424][6] , \registers[424][5] ,
         \registers[424][4] , \registers[424][3] , \registers[424][2] ,
         \registers[424][1] , \registers[424][0] , \registers[423][7] ,
         \registers[423][6] , \registers[423][5] , \registers[423][4] ,
         \registers[423][3] , \registers[423][2] , \registers[423][1] ,
         \registers[423][0] , \registers[422][7] , \registers[422][6] ,
         \registers[422][5] , \registers[422][4] , \registers[422][3] ,
         \registers[422][2] , \registers[422][1] , \registers[422][0] ,
         \registers[421][7] , \registers[421][6] , \registers[421][5] ,
         \registers[421][4] , \registers[421][3] , \registers[421][2] ,
         \registers[421][1] , \registers[421][0] , \registers[420][7] ,
         \registers[420][6] , \registers[420][5] , \registers[420][4] ,
         \registers[420][3] , \registers[420][2] , \registers[420][1] ,
         \registers[420][0] , \registers[419][7] , \registers[419][6] ,
         \registers[419][5] , \registers[419][4] , \registers[419][3] ,
         \registers[419][2] , \registers[419][1] , \registers[419][0] ,
         \registers[418][7] , \registers[418][6] , \registers[418][5] ,
         \registers[418][4] , \registers[418][3] , \registers[418][2] ,
         \registers[418][1] , \registers[418][0] , \registers[417][7] ,
         \registers[417][6] , \registers[417][5] , \registers[417][4] ,
         \registers[417][3] , \registers[417][2] , \registers[417][1] ,
         \registers[417][0] , \registers[416][7] , \registers[416][6] ,
         \registers[416][5] , \registers[416][4] , \registers[416][3] ,
         \registers[416][2] , \registers[416][1] , \registers[416][0] ,
         \registers[479][7] , \registers[479][6] , \registers[479][5] ,
         \registers[479][4] , \registers[479][3] , \registers[479][2] ,
         \registers[479][1] , \registers[479][0] , \registers[478][7] ,
         \registers[478][6] , \registers[478][5] , \registers[478][4] ,
         \registers[478][3] , \registers[478][2] , \registers[478][1] ,
         \registers[478][0] , \registers[477][7] , \registers[477][6] ,
         \registers[477][5] , \registers[477][4] , \registers[477][3] ,
         \registers[477][2] , \registers[477][1] , \registers[477][0] ,
         \registers[476][7] , \registers[476][6] , \registers[476][5] ,
         \registers[476][4] , \registers[476][3] , \registers[476][2] ,
         \registers[476][1] , \registers[476][0] , \registers[475][7] ,
         \registers[475][6] , \registers[475][5] , \registers[475][4] ,
         \registers[475][3] , \registers[475][2] , \registers[475][1] ,
         \registers[475][0] , \registers[474][7] , \registers[474][6] ,
         \registers[474][5] , \registers[474][4] , \registers[474][3] ,
         \registers[474][2] , \registers[474][1] , \registers[474][0] ,
         \registers[473][7] , \registers[473][6] , \registers[473][5] ,
         \registers[473][4] , \registers[473][3] , \registers[473][2] ,
         \registers[473][1] , \registers[473][0] , \registers[472][7] ,
         \registers[472][6] , \registers[472][5] , \registers[472][4] ,
         \registers[472][3] , \registers[472][2] , \registers[472][1] ,
         \registers[472][0] , \registers[471][7] , \registers[471][6] ,
         \registers[471][5] , \registers[471][4] , \registers[471][3] ,
         \registers[471][2] , \registers[471][1] , \registers[471][0] ,
         \registers[470][7] , \registers[470][6] , \registers[470][5] ,
         \registers[470][4] , \registers[470][3] , \registers[470][2] ,
         \registers[470][1] , \registers[470][0] , \registers[469][7] ,
         \registers[469][6] , \registers[469][5] , \registers[469][4] ,
         \registers[469][3] , \registers[469][2] , \registers[469][1] ,
         \registers[469][0] , \registers[468][7] , \registers[468][6] ,
         \registers[468][5] , \registers[468][4] , \registers[468][3] ,
         \registers[468][2] , \registers[468][1] , \registers[468][0] ,
         \registers[467][7] , \registers[467][6] , \registers[467][5] ,
         \registers[467][4] , \registers[467][3] , \registers[467][2] ,
         \registers[467][1] , \registers[467][0] , \registers[466][7] ,
         \registers[466][6] , \registers[466][5] , \registers[466][4] ,
         \registers[466][3] , \registers[466][2] , \registers[466][1] ,
         \registers[466][0] , \registers[465][7] , \registers[465][6] ,
         \registers[465][5] , \registers[465][4] , \registers[465][3] ,
         \registers[465][2] , \registers[465][1] , \registers[465][0] ,
         \registers[464][7] , \registers[464][6] , \registers[464][5] ,
         \registers[464][4] , \registers[464][3] , \registers[464][2] ,
         \registers[464][1] , \registers[464][0] , \registers[463][7] ,
         \registers[463][6] , \registers[463][5] , \registers[463][4] ,
         \registers[463][3] , \registers[463][2] , \registers[463][1] ,
         \registers[463][0] , \registers[462][7] , \registers[462][6] ,
         \registers[462][5] , \registers[462][4] , \registers[462][3] ,
         \registers[462][2] , \registers[462][1] , \registers[462][0] ,
         \registers[461][7] , \registers[461][6] , \registers[461][5] ,
         \registers[461][4] , \registers[461][3] , \registers[461][2] ,
         \registers[461][1] , \registers[461][0] , \registers[460][7] ,
         \registers[460][6] , \registers[460][5] , \registers[460][4] ,
         \registers[460][3] , \registers[460][2] , \registers[460][1] ,
         \registers[460][0] , \registers[459][7] , \registers[459][6] ,
         \registers[459][5] , \registers[459][4] , \registers[459][3] ,
         \registers[459][2] , \registers[459][1] , \registers[459][0] ,
         \registers[458][7] , \registers[458][6] , \registers[458][5] ,
         \registers[458][4] , \registers[458][3] , \registers[458][2] ,
         \registers[458][1] , \registers[458][0] , \registers[457][7] ,
         \registers[457][6] , \registers[457][5] , \registers[457][4] ,
         \registers[457][3] , \registers[457][2] , \registers[457][1] ,
         \registers[457][0] , \registers[456][7] , \registers[456][6] ,
         \registers[456][5] , \registers[456][4] , \registers[456][3] ,
         \registers[456][2] , \registers[456][1] , \registers[456][0] ,
         \registers[455][7] , \registers[455][6] , \registers[455][5] ,
         \registers[455][4] , \registers[455][3] , \registers[455][2] ,
         \registers[455][1] , \registers[455][0] , \registers[454][7] ,
         \registers[454][6] , \registers[454][5] , \registers[454][4] ,
         \registers[454][3] , \registers[454][2] , \registers[454][1] ,
         \registers[454][0] , \registers[453][7] , \registers[453][6] ,
         \registers[453][5] , \registers[453][4] , \registers[453][3] ,
         \registers[453][2] , \registers[453][1] , \registers[453][0] ,
         \registers[452][7] , \registers[452][6] , \registers[452][5] ,
         \registers[452][4] , \registers[452][3] , \registers[452][2] ,
         \registers[452][1] , \registers[452][0] , \registers[451][7] ,
         \registers[451][6] , \registers[451][5] , \registers[451][4] ,
         \registers[451][3] , \registers[451][2] , \registers[451][1] ,
         \registers[451][0] , \registers[450][7] , \registers[450][6] ,
         \registers[450][5] , \registers[450][4] , \registers[450][3] ,
         \registers[450][2] , \registers[450][1] , \registers[450][0] ,
         \registers[449][7] , \registers[449][6] , \registers[449][5] ,
         \registers[449][4] , \registers[449][3] , \registers[449][2] ,
         \registers[449][1] , \registers[449][0] , \registers[448][7] ,
         \registers[448][6] , \registers[448][5] , \registers[448][4] ,
         \registers[448][3] , \registers[448][2] , \registers[448][1] ,
         \registers[448][0] , \registers[511][7] , \registers[511][6] ,
         \registers[511][5] , \registers[511][4] , \registers[511][3] ,
         \registers[511][2] , \registers[511][1] , \registers[511][0] ,
         \registers[510][7] , \registers[510][6] , \registers[510][5] ,
         \registers[510][4] , \registers[510][3] , \registers[510][2] ,
         \registers[510][1] , \registers[510][0] , \registers[509][7] ,
         \registers[509][6] , \registers[509][5] , \registers[509][4] ,
         \registers[509][3] , \registers[509][2] , \registers[509][1] ,
         \registers[509][0] , \registers[508][7] , \registers[508][6] ,
         \registers[508][5] , \registers[508][4] , \registers[508][3] ,
         \registers[508][2] , \registers[508][1] , \registers[508][0] ,
         \registers[507][7] , \registers[507][6] , \registers[507][5] ,
         \registers[507][4] , \registers[507][3] , \registers[507][2] ,
         \registers[507][1] , \registers[507][0] , \registers[506][7] ,
         \registers[506][6] , \registers[506][5] , \registers[506][4] ,
         \registers[506][3] , \registers[506][2] , \registers[506][1] ,
         \registers[506][0] , \registers[505][7] , \registers[505][6] ,
         \registers[505][5] , \registers[505][4] , \registers[505][3] ,
         \registers[505][2] , \registers[505][1] , \registers[505][0] ,
         \registers[504][7] , \registers[504][6] , \registers[504][5] ,
         \registers[504][4] , \registers[504][3] , \registers[504][2] ,
         \registers[504][1] , \registers[504][0] , \registers[503][7] ,
         \registers[503][6] , \registers[503][5] , \registers[503][4] ,
         \registers[503][3] , \registers[503][2] , \registers[503][1] ,
         \registers[503][0] , \registers[502][7] , \registers[502][6] ,
         \registers[502][5] , \registers[502][4] , \registers[502][3] ,
         \registers[502][2] , \registers[502][1] , \registers[502][0] ,
         \registers[501][7] , \registers[501][6] , \registers[501][5] ,
         \registers[501][4] , \registers[501][3] , \registers[501][2] ,
         \registers[501][1] , \registers[501][0] , \registers[500][7] ,
         \registers[500][6] , \registers[500][5] , \registers[500][4] ,
         \registers[500][3] , \registers[500][2] , \registers[500][1] ,
         \registers[500][0] , \registers[499][7] , \registers[499][6] ,
         \registers[499][5] , \registers[499][4] , \registers[499][3] ,
         \registers[499][2] , \registers[499][1] , \registers[499][0] ,
         \registers[498][7] , \registers[498][6] , \registers[498][5] ,
         \registers[498][4] , \registers[498][3] , \registers[498][2] ,
         \registers[498][1] , \registers[498][0] , \registers[497][7] ,
         \registers[497][6] , \registers[497][5] , \registers[497][4] ,
         \registers[497][3] , \registers[497][2] , \registers[497][1] ,
         \registers[497][0] , \registers[496][7] , \registers[496][6] ,
         \registers[496][5] , \registers[496][4] , \registers[496][3] ,
         \registers[496][2] , \registers[496][1] , \registers[496][0] ,
         \registers[495][7] , \registers[495][6] , \registers[495][5] ,
         \registers[495][4] , \registers[495][3] , \registers[495][2] ,
         \registers[495][1] , \registers[495][0] , \registers[494][7] ,
         \registers[494][6] , \registers[494][5] , \registers[494][4] ,
         \registers[494][3] , \registers[494][2] , \registers[494][1] ,
         \registers[494][0] , \registers[493][7] , \registers[493][6] ,
         \registers[493][5] , \registers[493][4] , \registers[493][3] ,
         \registers[493][2] , \registers[493][1] , \registers[493][0] ,
         \registers[492][7] , \registers[492][6] , \registers[492][5] ,
         \registers[492][4] , \registers[492][3] , \registers[492][2] ,
         \registers[492][1] , \registers[492][0] , \registers[491][7] ,
         \registers[491][6] , \registers[491][5] , \registers[491][4] ,
         \registers[491][3] , \registers[491][2] , \registers[491][1] ,
         \registers[491][0] , \registers[490][7] , \registers[490][6] ,
         \registers[490][5] , \registers[490][4] , \registers[490][3] ,
         \registers[490][2] , \registers[490][1] , \registers[490][0] ,
         \registers[489][7] , \registers[489][6] , \registers[489][5] ,
         \registers[489][4] , \registers[489][3] , \registers[489][2] ,
         \registers[489][1] , \registers[489][0] , \registers[488][7] ,
         \registers[488][6] , \registers[488][5] , \registers[488][4] ,
         \registers[488][3] , \registers[488][2] , \registers[488][1] ,
         \registers[488][0] , \registers[487][7] , \registers[487][6] ,
         \registers[487][5] , \registers[487][4] , \registers[487][3] ,
         \registers[487][2] , \registers[487][1] , \registers[487][0] ,
         \registers[486][7] , \registers[486][6] , \registers[486][5] ,
         \registers[486][4] , \registers[486][3] , \registers[486][2] ,
         \registers[486][1] , \registers[486][0] , \registers[485][7] ,
         \registers[485][6] , \registers[485][5] , \registers[485][4] ,
         \registers[485][3] , \registers[485][2] , \registers[485][1] ,
         \registers[485][0] , \registers[484][7] , \registers[484][6] ,
         \registers[484][5] , \registers[484][4] , \registers[484][3] ,
         \registers[484][2] , \registers[484][1] , \registers[484][0] ,
         \registers[483][7] , \registers[483][6] , \registers[483][5] ,
         \registers[483][4] , \registers[483][3] , \registers[483][2] ,
         \registers[483][1] , \registers[483][0] , \registers[482][7] ,
         \registers[482][6] , \registers[482][5] , \registers[482][4] ,
         \registers[482][3] , \registers[482][2] , \registers[482][1] ,
         \registers[482][0] , \registers[481][7] , \registers[481][6] ,
         \registers[481][5] , \registers[481][4] , \registers[481][3] ,
         \registers[481][2] , \registers[481][1] , \registers[481][0] ,
         \registers[480][7] , \registers[480][6] , \registers[480][5] ,
         \registers[480][4] , \registers[480][3] , \registers[480][2] ,
         \registers[480][1] , \registers[480][0] , \registers[543][7] ,
         \registers[543][6] , \registers[543][5] , \registers[543][4] ,
         \registers[543][3] , \registers[543][2] , \registers[543][1] ,
         \registers[543][0] , \registers[542][7] , \registers[542][6] ,
         \registers[542][5] , \registers[542][4] , \registers[542][3] ,
         \registers[542][2] , \registers[542][1] , \registers[542][0] ,
         \registers[541][7] , \registers[541][6] , \registers[541][5] ,
         \registers[541][4] , \registers[541][3] , \registers[541][2] ,
         \registers[541][1] , \registers[541][0] , \registers[540][7] ,
         \registers[540][6] , \registers[540][5] , \registers[540][4] ,
         \registers[540][3] , \registers[540][2] , \registers[540][1] ,
         \registers[540][0] , \registers[539][7] , \registers[539][6] ,
         \registers[539][5] , \registers[539][4] , \registers[539][3] ,
         \registers[539][2] , \registers[539][1] , \registers[539][0] ,
         \registers[538][7] , \registers[538][6] , \registers[538][5] ,
         \registers[538][4] , \registers[538][3] , \registers[538][2] ,
         \registers[538][1] , \registers[538][0] , \registers[537][7] ,
         \registers[537][6] , \registers[537][5] , \registers[537][4] ,
         \registers[537][3] , \registers[537][2] , \registers[537][1] ,
         \registers[537][0] , \registers[536][7] , \registers[536][6] ,
         \registers[536][5] , \registers[536][4] , \registers[536][3] ,
         \registers[536][2] , \registers[536][1] , \registers[536][0] ,
         \registers[535][7] , \registers[535][6] , \registers[535][5] ,
         \registers[535][4] , \registers[535][3] , \registers[535][2] ,
         \registers[535][1] , \registers[535][0] , \registers[534][7] ,
         \registers[534][6] , \registers[534][5] , \registers[534][4] ,
         \registers[534][3] , \registers[534][2] , \registers[534][1] ,
         \registers[534][0] , \registers[533][7] , \registers[533][6] ,
         \registers[533][5] , \registers[533][4] , \registers[533][3] ,
         \registers[533][2] , \registers[533][1] , \registers[533][0] ,
         \registers[532][7] , \registers[532][6] , \registers[532][5] ,
         \registers[532][4] , \registers[532][3] , \registers[532][2] ,
         \registers[532][1] , \registers[532][0] , \registers[531][7] ,
         \registers[531][6] , \registers[531][5] , \registers[531][4] ,
         \registers[531][3] , \registers[531][2] , \registers[531][1] ,
         \registers[531][0] , \registers[530][7] , \registers[530][6] ,
         \registers[530][5] , \registers[530][4] , \registers[530][3] ,
         \registers[530][2] , \registers[530][1] , \registers[530][0] ,
         \registers[529][7] , \registers[529][6] , \registers[529][5] ,
         \registers[529][4] , \registers[529][3] , \registers[529][2] ,
         \registers[529][1] , \registers[529][0] , \registers[528][7] ,
         \registers[528][6] , \registers[528][5] , \registers[528][4] ,
         \registers[528][3] , \registers[528][2] , \registers[528][1] ,
         \registers[528][0] , \registers[527][7] , \registers[527][6] ,
         \registers[527][5] , \registers[527][4] , \registers[527][3] ,
         \registers[527][2] , \registers[527][1] , \registers[527][0] ,
         \registers[526][7] , \registers[526][6] , \registers[526][5] ,
         \registers[526][4] , \registers[526][3] , \registers[526][2] ,
         \registers[526][1] , \registers[526][0] , \registers[525][7] ,
         \registers[525][6] , \registers[525][5] , \registers[525][4] ,
         \registers[525][3] , \registers[525][2] , \registers[525][1] ,
         \registers[525][0] , \registers[524][7] , \registers[524][6] ,
         \registers[524][5] , \registers[524][4] , \registers[524][3] ,
         \registers[524][2] , \registers[524][1] , \registers[524][0] ,
         \registers[523][7] , \registers[523][6] , \registers[523][5] ,
         \registers[523][4] , \registers[523][3] , \registers[523][2] ,
         \registers[523][1] , \registers[523][0] , \registers[522][7] ,
         \registers[522][6] , \registers[522][5] , \registers[522][4] ,
         \registers[522][3] , \registers[522][2] , \registers[522][1] ,
         \registers[522][0] , \registers[521][7] , \registers[521][6] ,
         \registers[521][5] , \registers[521][4] , \registers[521][3] ,
         \registers[521][2] , \registers[521][1] , \registers[521][0] ,
         \registers[520][7] , \registers[520][6] , \registers[520][5] ,
         \registers[520][4] , \registers[520][3] , \registers[520][2] ,
         \registers[520][1] , \registers[520][0] , \registers[519][7] ,
         \registers[519][6] , \registers[519][5] , \registers[519][4] ,
         \registers[519][3] , \registers[519][2] , \registers[519][1] ,
         \registers[519][0] , \registers[518][7] , \registers[518][6] ,
         \registers[518][5] , \registers[518][4] , \registers[518][3] ,
         \registers[518][2] , \registers[518][1] , \registers[518][0] ,
         \registers[517][7] , \registers[517][6] , \registers[517][5] ,
         \registers[517][4] , \registers[517][3] , \registers[517][2] ,
         \registers[517][1] , \registers[517][0] , \registers[516][7] ,
         \registers[516][6] , \registers[516][5] , \registers[516][4] ,
         \registers[516][3] , \registers[516][2] , \registers[516][1] ,
         \registers[516][0] , \registers[515][7] , \registers[515][6] ,
         \registers[515][5] , \registers[515][4] , \registers[515][3] ,
         \registers[515][2] , \registers[515][1] , \registers[515][0] ,
         \registers[514][7] , \registers[514][6] , \registers[514][5] ,
         \registers[514][4] , \registers[514][3] , \registers[514][2] ,
         \registers[514][1] , \registers[514][0] , \registers[513][7] ,
         \registers[513][6] , \registers[513][5] , \registers[513][4] ,
         \registers[513][3] , \registers[513][2] , \registers[513][1] ,
         \registers[513][0] , \registers[512][7] , \registers[512][6] ,
         \registers[512][5] , \registers[512][4] , \registers[512][3] ,
         \registers[512][2] , \registers[512][1] , \registers[512][0] ,
         \registers[575][7] , \registers[575][6] , \registers[575][5] ,
         \registers[575][4] , \registers[575][3] , \registers[575][2] ,
         \registers[575][1] , \registers[575][0] , \registers[574][7] ,
         \registers[574][6] , \registers[574][5] , \registers[574][4] ,
         \registers[574][3] , \registers[574][2] , \registers[574][1] ,
         \registers[574][0] , \registers[573][7] , \registers[573][6] ,
         \registers[573][5] , \registers[573][4] , \registers[573][3] ,
         \registers[573][2] , \registers[573][1] , \registers[573][0] ,
         \registers[572][7] , \registers[572][6] , \registers[572][5] ,
         \registers[572][4] , \registers[572][3] , \registers[572][2] ,
         \registers[572][1] , \registers[572][0] , \registers[571][7] ,
         \registers[571][6] , \registers[571][5] , \registers[571][4] ,
         \registers[571][3] , \registers[571][2] , \registers[571][1] ,
         \registers[571][0] , \registers[570][7] , \registers[570][6] ,
         \registers[570][5] , \registers[570][4] , \registers[570][3] ,
         \registers[570][2] , \registers[570][1] , \registers[570][0] ,
         \registers[569][7] , \registers[569][6] , \registers[569][5] ,
         \registers[569][4] , \registers[569][3] , \registers[569][2] ,
         \registers[569][1] , \registers[569][0] , \registers[568][7] ,
         \registers[568][6] , \registers[568][5] , \registers[568][4] ,
         \registers[568][3] , \registers[568][2] , \registers[568][1] ,
         \registers[568][0] , \registers[567][7] , \registers[567][6] ,
         \registers[567][5] , \registers[567][4] , \registers[567][3] ,
         \registers[567][2] , \registers[567][1] , \registers[567][0] ,
         \registers[566][7] , \registers[566][6] , \registers[566][5] ,
         \registers[566][4] , \registers[566][3] , \registers[566][2] ,
         \registers[566][1] , \registers[566][0] , \registers[565][7] ,
         \registers[565][6] , \registers[565][5] , \registers[565][4] ,
         \registers[565][3] , \registers[565][2] , \registers[565][1] ,
         \registers[565][0] , \registers[564][7] , \registers[564][6] ,
         \registers[564][5] , \registers[564][4] , \registers[564][3] ,
         \registers[564][2] , \registers[564][1] , \registers[564][0] ,
         \registers[563][7] , \registers[563][6] , \registers[563][5] ,
         \registers[563][4] , \registers[563][3] , \registers[563][2] ,
         \registers[563][1] , \registers[563][0] , \registers[562][7] ,
         \registers[562][6] , \registers[562][5] , \registers[562][4] ,
         \registers[562][3] , \registers[562][2] , \registers[562][1] ,
         \registers[562][0] , \registers[561][7] , \registers[561][6] ,
         \registers[561][5] , \registers[561][4] , \registers[561][3] ,
         \registers[561][2] , \registers[561][1] , \registers[561][0] ,
         \registers[560][7] , \registers[560][6] , \registers[560][5] ,
         \registers[560][4] , \registers[560][3] , \registers[560][2] ,
         \registers[560][1] , \registers[560][0] , \registers[559][7] ,
         \registers[559][6] , \registers[559][5] , \registers[559][4] ,
         \registers[559][3] , \registers[559][2] , \registers[559][1] ,
         \registers[559][0] , \registers[558][7] , \registers[558][6] ,
         \registers[558][5] , \registers[558][4] , \registers[558][3] ,
         \registers[558][2] , \registers[558][1] , \registers[558][0] ,
         \registers[557][7] , \registers[557][6] , \registers[557][5] ,
         \registers[557][4] , \registers[557][3] , \registers[557][2] ,
         \registers[557][1] , \registers[557][0] , \registers[556][7] ,
         \registers[556][6] , \registers[556][5] , \registers[556][4] ,
         \registers[556][3] , \registers[556][2] , \registers[556][1] ,
         \registers[556][0] , \registers[555][7] , \registers[555][6] ,
         \registers[555][5] , \registers[555][4] , \registers[555][3] ,
         \registers[555][2] , \registers[555][1] , \registers[555][0] ,
         \registers[554][7] , \registers[554][6] , \registers[554][5] ,
         \registers[554][4] , \registers[554][3] , \registers[554][2] ,
         \registers[554][1] , \registers[554][0] , \registers[553][7] ,
         \registers[553][6] , \registers[553][5] , \registers[553][4] ,
         \registers[553][3] , \registers[553][2] , \registers[553][1] ,
         \registers[553][0] , \registers[552][7] , \registers[552][6] ,
         \registers[552][5] , \registers[552][4] , \registers[552][3] ,
         \registers[552][2] , \registers[552][1] , \registers[552][0] ,
         \registers[551][7] , \registers[551][6] , \registers[551][5] ,
         \registers[551][4] , \registers[551][3] , \registers[551][2] ,
         \registers[551][1] , \registers[551][0] , \registers[550][7] ,
         \registers[550][6] , \registers[550][5] , \registers[550][4] ,
         \registers[550][3] , \registers[550][2] , \registers[550][1] ,
         \registers[550][0] , \registers[549][7] , \registers[549][6] ,
         \registers[549][5] , \registers[549][4] , \registers[549][3] ,
         \registers[549][2] , \registers[549][1] , \registers[549][0] ,
         \registers[548][7] , \registers[548][6] , \registers[548][5] ,
         \registers[548][4] , \registers[548][3] , \registers[548][2] ,
         \registers[548][1] , \registers[548][0] , \registers[547][7] ,
         \registers[547][6] , \registers[547][5] , \registers[547][4] ,
         \registers[547][3] , \registers[547][2] , \registers[547][1] ,
         \registers[547][0] , \registers[546][7] , \registers[546][6] ,
         \registers[546][5] , \registers[546][4] , \registers[546][3] ,
         \registers[546][2] , \registers[546][1] , \registers[546][0] ,
         \registers[545][7] , \registers[545][6] , \registers[545][5] ,
         \registers[545][4] , \registers[545][3] , \registers[545][2] ,
         \registers[545][1] , \registers[545][0] , \registers[544][7] ,
         \registers[544][6] , \registers[544][5] , \registers[544][4] ,
         \registers[544][3] , \registers[544][2] , \registers[544][1] ,
         \registers[544][0] , \registers[607][7] , \registers[607][6] ,
         \registers[607][5] , \registers[607][4] , \registers[607][3] ,
         \registers[607][2] , \registers[607][1] , \registers[607][0] ,
         \registers[606][7] , \registers[606][6] , \registers[606][5] ,
         \registers[606][4] , \registers[606][3] , \registers[606][2] ,
         \registers[606][1] , \registers[606][0] , \registers[605][7] ,
         \registers[605][6] , \registers[605][5] , \registers[605][4] ,
         \registers[605][3] , \registers[605][2] , \registers[605][1] ,
         \registers[605][0] , \registers[604][7] , \registers[604][6] ,
         \registers[604][5] , \registers[604][4] , \registers[604][3] ,
         \registers[604][2] , \registers[604][1] , \registers[604][0] ,
         \registers[603][7] , \registers[603][6] , \registers[603][5] ,
         \registers[603][4] , \registers[603][3] , \registers[603][2] ,
         \registers[603][1] , \registers[603][0] , \registers[602][7] ,
         \registers[602][6] , \registers[602][5] , \registers[602][4] ,
         \registers[602][3] , \registers[602][2] , \registers[602][1] ,
         \registers[602][0] , \registers[601][7] , \registers[601][6] ,
         \registers[601][5] , \registers[601][4] , \registers[601][3] ,
         \registers[601][2] , \registers[601][1] , \registers[601][0] ,
         \registers[600][7] , \registers[600][6] , \registers[600][5] ,
         \registers[600][4] , \registers[600][3] , \registers[600][2] ,
         \registers[600][1] , \registers[600][0] , \registers[599][7] ,
         \registers[599][6] , \registers[599][5] , \registers[599][4] ,
         \registers[599][3] , \registers[599][2] , \registers[599][1] ,
         \registers[599][0] , \registers[598][7] , \registers[598][6] ,
         \registers[598][5] , \registers[598][4] , \registers[598][3] ,
         \registers[598][2] , \registers[598][1] , \registers[598][0] ,
         \registers[597][7] , \registers[597][6] , \registers[597][5] ,
         \registers[597][4] , \registers[597][3] , \registers[597][2] ,
         \registers[597][1] , \registers[597][0] , \registers[596][7] ,
         \registers[596][6] , \registers[596][5] , \registers[596][4] ,
         \registers[596][3] , \registers[596][2] , \registers[596][1] ,
         \registers[596][0] , \registers[595][7] , \registers[595][6] ,
         \registers[595][5] , \registers[595][4] , \registers[595][3] ,
         \registers[595][2] , \registers[595][1] , \registers[595][0] ,
         \registers[594][7] , \registers[594][6] , \registers[594][5] ,
         \registers[594][4] , \registers[594][3] , \registers[594][2] ,
         \registers[594][1] , \registers[594][0] , \registers[593][7] ,
         \registers[593][6] , \registers[593][5] , \registers[593][4] ,
         \registers[593][3] , \registers[593][2] , \registers[593][1] ,
         \registers[593][0] , \registers[592][7] , \registers[592][6] ,
         \registers[592][5] , \registers[592][4] , \registers[592][3] ,
         \registers[592][2] , \registers[592][1] , \registers[592][0] ,
         \registers[591][7] , \registers[591][6] , \registers[591][5] ,
         \registers[591][4] , \registers[591][3] , \registers[591][2] ,
         \registers[591][1] , \registers[591][0] , \registers[590][7] ,
         \registers[590][6] , \registers[590][5] , \registers[590][4] ,
         \registers[590][3] , \registers[590][2] , \registers[590][1] ,
         \registers[590][0] , \registers[589][7] , \registers[589][6] ,
         \registers[589][5] , \registers[589][4] , \registers[589][3] ,
         \registers[589][2] , \registers[589][1] , \registers[589][0] ,
         \registers[588][7] , \registers[588][6] , \registers[588][5] ,
         \registers[588][4] , \registers[588][3] , \registers[588][2] ,
         \registers[588][1] , \registers[588][0] , \registers[587][7] ,
         \registers[587][6] , \registers[587][5] , \registers[587][4] ,
         \registers[587][3] , \registers[587][2] , \registers[587][1] ,
         \registers[587][0] , \registers[586][7] , \registers[586][6] ,
         \registers[586][5] , \registers[586][4] , \registers[586][3] ,
         \registers[586][2] , \registers[586][1] , \registers[586][0] ,
         \registers[585][7] , \registers[585][6] , \registers[585][5] ,
         \registers[585][4] , \registers[585][3] , \registers[585][2] ,
         \registers[585][1] , \registers[585][0] , \registers[584][7] ,
         \registers[584][6] , \registers[584][5] , \registers[584][4] ,
         \registers[584][3] , \registers[584][2] , \registers[584][1] ,
         \registers[584][0] , \registers[583][7] , \registers[583][6] ,
         \registers[583][5] , \registers[583][4] , \registers[583][3] ,
         \registers[583][2] , \registers[583][1] , \registers[583][0] ,
         \registers[582][7] , \registers[582][6] , \registers[582][5] ,
         \registers[582][4] , \registers[582][3] , \registers[582][2] ,
         \registers[582][1] , \registers[582][0] , \registers[581][7] ,
         \registers[581][6] , \registers[581][5] , \registers[581][4] ,
         \registers[581][3] , \registers[581][2] , \registers[581][1] ,
         \registers[581][0] , \registers[580][7] , \registers[580][6] ,
         \registers[580][5] , \registers[580][4] , \registers[580][3] ,
         \registers[580][2] , \registers[580][1] , \registers[580][0] ,
         \registers[579][7] , \registers[579][6] , \registers[579][5] ,
         \registers[579][4] , \registers[579][3] , \registers[579][2] ,
         \registers[579][1] , \registers[579][0] , \registers[578][7] ,
         \registers[578][6] , \registers[578][5] , \registers[578][4] ,
         \registers[578][3] , \registers[578][2] , \registers[578][1] ,
         \registers[578][0] , \registers[577][7] , \registers[577][6] ,
         \registers[577][5] , \registers[577][4] , \registers[577][3] ,
         \registers[577][2] , \registers[577][1] , \registers[577][0] ,
         \registers[576][7] , \registers[576][6] , \registers[576][5] ,
         \registers[576][4] , \registers[576][3] , \registers[576][2] ,
         \registers[576][1] , \registers[576][0] , \registers[639][7] ,
         \registers[639][6] , \registers[639][5] , \registers[639][4] ,
         \registers[639][3] , \registers[639][2] , \registers[639][1] ,
         \registers[639][0] , \registers[638][7] , \registers[638][6] ,
         \registers[638][5] , \registers[638][4] , \registers[638][3] ,
         \registers[638][2] , \registers[638][1] , \registers[638][0] ,
         \registers[637][7] , \registers[637][6] , \registers[637][5] ,
         \registers[637][4] , \registers[637][3] , \registers[637][2] ,
         \registers[637][1] , \registers[637][0] , \registers[636][7] ,
         \registers[636][6] , \registers[636][5] , \registers[636][4] ,
         \registers[636][3] , \registers[636][2] , \registers[636][1] ,
         \registers[636][0] , \registers[635][7] , \registers[635][6] ,
         \registers[635][5] , \registers[635][4] , \registers[635][3] ,
         \registers[635][2] , \registers[635][1] , \registers[635][0] ,
         \registers[634][7] , \registers[634][6] , \registers[634][5] ,
         \registers[634][4] , \registers[634][3] , \registers[634][2] ,
         \registers[634][1] , \registers[634][0] , \registers[633][7] ,
         \registers[633][6] , \registers[633][5] , \registers[633][4] ,
         \registers[633][3] , \registers[633][2] , \registers[633][1] ,
         \registers[633][0] , \registers[632][7] , \registers[632][6] ,
         \registers[632][5] , \registers[632][4] , \registers[632][3] ,
         \registers[632][2] , \registers[632][1] , \registers[632][0] ,
         \registers[631][7] , \registers[631][6] , \registers[631][5] ,
         \registers[631][4] , \registers[631][3] , \registers[631][2] ,
         \registers[631][1] , \registers[631][0] , \registers[630][7] ,
         \registers[630][6] , \registers[630][5] , \registers[630][4] ,
         \registers[630][3] , \registers[630][2] , \registers[630][1] ,
         \registers[630][0] , \registers[629][7] , \registers[629][6] ,
         \registers[629][5] , \registers[629][4] , \registers[629][3] ,
         \registers[629][2] , \registers[629][1] , \registers[629][0] ,
         \registers[628][7] , \registers[628][6] , \registers[628][5] ,
         \registers[628][4] , \registers[628][3] , \registers[628][2] ,
         \registers[628][1] , \registers[628][0] , \registers[627][7] ,
         \registers[627][6] , \registers[627][5] , \registers[627][4] ,
         \registers[627][3] , \registers[627][2] , \registers[627][1] ,
         \registers[627][0] , \registers[626][7] , \registers[626][6] ,
         \registers[626][5] , \registers[626][4] , \registers[626][3] ,
         \registers[626][2] , \registers[626][1] , \registers[626][0] ,
         \registers[625][7] , \registers[625][6] , \registers[625][5] ,
         \registers[625][4] , \registers[625][3] , \registers[625][2] ,
         \registers[625][1] , \registers[625][0] , \registers[624][7] ,
         \registers[624][6] , \registers[624][5] , \registers[624][4] ,
         \registers[624][3] , \registers[624][2] , \registers[624][1] ,
         \registers[624][0] , \registers[623][7] , \registers[623][6] ,
         \registers[623][5] , \registers[623][4] , \registers[623][3] ,
         \registers[623][2] , \registers[623][1] , \registers[623][0] ,
         \registers[622][7] , \registers[622][6] , \registers[622][5] ,
         \registers[622][4] , \registers[622][3] , \registers[622][2] ,
         \registers[622][1] , \registers[622][0] , \registers[621][7] ,
         \registers[621][6] , \registers[621][5] , \registers[621][4] ,
         \registers[621][3] , \registers[621][2] , \registers[621][1] ,
         \registers[621][0] , \registers[620][7] , \registers[620][6] ,
         \registers[620][5] , \registers[620][4] , \registers[620][3] ,
         \registers[620][2] , \registers[620][1] , \registers[620][0] ,
         \registers[619][7] , \registers[619][6] , \registers[619][5] ,
         \registers[619][4] , \registers[619][3] , \registers[619][2] ,
         \registers[619][1] , \registers[619][0] , \registers[618][7] ,
         \registers[618][6] , \registers[618][5] , \registers[618][4] ,
         \registers[618][3] , \registers[618][2] , \registers[618][1] ,
         \registers[618][0] , \registers[617][7] , \registers[617][6] ,
         \registers[617][5] , \registers[617][4] , \registers[617][3] ,
         \registers[617][2] , \registers[617][1] , \registers[617][0] ,
         \registers[616][7] , \registers[616][6] , \registers[616][5] ,
         \registers[616][4] , \registers[616][3] , \registers[616][2] ,
         \registers[616][1] , \registers[616][0] , \registers[615][7] ,
         \registers[615][6] , \registers[615][5] , \registers[615][4] ,
         \registers[615][3] , \registers[615][2] , \registers[615][1] ,
         \registers[615][0] , \registers[614][7] , \registers[614][6] ,
         \registers[614][5] , \registers[614][4] , \registers[614][3] ,
         \registers[614][2] , \registers[614][1] , \registers[614][0] ,
         \registers[613][7] , \registers[613][6] , \registers[613][5] ,
         \registers[613][4] , \registers[613][3] , \registers[613][2] ,
         \registers[613][1] , \registers[613][0] , \registers[612][7] ,
         \registers[612][6] , \registers[612][5] , \registers[612][4] ,
         \registers[612][3] , \registers[612][2] , \registers[612][1] ,
         \registers[612][0] , \registers[611][7] , \registers[611][6] ,
         \registers[611][5] , \registers[611][4] , \registers[611][3] ,
         \registers[611][2] , \registers[611][1] , \registers[611][0] ,
         \registers[610][7] , \registers[610][6] , \registers[610][5] ,
         \registers[610][4] , \registers[610][3] , \registers[610][2] ,
         \registers[610][1] , \registers[610][0] , \registers[609][7] ,
         \registers[609][6] , \registers[609][5] , \registers[609][4] ,
         \registers[609][3] , \registers[609][2] , \registers[609][1] ,
         \registers[609][0] , \registers[608][7] , \registers[608][6] ,
         \registers[608][5] , \registers[608][4] , \registers[608][3] ,
         \registers[608][2] , \registers[608][1] , \registers[608][0] ,
         \registers[671][7] , \registers[671][6] , \registers[671][5] ,
         \registers[671][4] , \registers[671][3] , \registers[671][2] ,
         \registers[671][1] , \registers[671][0] , \registers[670][7] ,
         \registers[670][6] , \registers[670][5] , \registers[670][4] ,
         \registers[670][3] , \registers[670][2] , \registers[670][1] ,
         \registers[670][0] , \registers[669][7] , \registers[669][6] ,
         \registers[669][5] , \registers[669][4] , \registers[669][3] ,
         \registers[669][2] , \registers[669][1] , \registers[669][0] ,
         \registers[668][7] , \registers[668][6] , \registers[668][5] ,
         \registers[668][4] , \registers[668][3] , \registers[668][2] ,
         \registers[668][1] , \registers[668][0] , \registers[667][7] ,
         \registers[667][6] , \registers[667][5] , \registers[667][4] ,
         \registers[667][3] , \registers[667][2] , \registers[667][1] ,
         \registers[667][0] , \registers[666][7] , \registers[666][6] ,
         \registers[666][5] , \registers[666][4] , \registers[666][3] ,
         \registers[666][2] , \registers[666][1] , \registers[666][0] ,
         \registers[665][7] , \registers[665][6] , \registers[665][5] ,
         \registers[665][4] , \registers[665][3] , \registers[665][2] ,
         \registers[665][1] , \registers[665][0] , \registers[664][7] ,
         \registers[664][6] , \registers[664][5] , \registers[664][4] ,
         \registers[664][3] , \registers[664][2] , \registers[664][1] ,
         \registers[664][0] , \registers[663][7] , \registers[663][6] ,
         \registers[663][5] , \registers[663][4] , \registers[663][3] ,
         \registers[663][2] , \registers[663][1] , \registers[663][0] ,
         \registers[662][7] , \registers[662][6] , \registers[662][5] ,
         \registers[662][4] , \registers[662][3] , \registers[662][2] ,
         \registers[662][1] , \registers[662][0] , \registers[661][7] ,
         \registers[661][6] , \registers[661][5] , \registers[661][4] ,
         \registers[661][3] , \registers[661][2] , \registers[661][1] ,
         \registers[661][0] , \registers[660][7] , \registers[660][6] ,
         \registers[660][5] , \registers[660][4] , \registers[660][3] ,
         \registers[660][2] , \registers[660][1] , \registers[660][0] ,
         \registers[659][7] , \registers[659][6] , \registers[659][5] ,
         \registers[659][4] , \registers[659][3] , \registers[659][2] ,
         \registers[659][1] , \registers[659][0] , \registers[658][7] ,
         \registers[658][6] , \registers[658][5] , \registers[658][4] ,
         \registers[658][3] , \registers[658][2] , \registers[658][1] ,
         \registers[658][0] , \registers[657][7] , \registers[657][6] ,
         \registers[657][5] , \registers[657][4] , \registers[657][3] ,
         \registers[657][2] , \registers[657][1] , \registers[657][0] ,
         \registers[656][7] , \registers[656][6] , \registers[656][5] ,
         \registers[656][4] , \registers[656][3] , \registers[656][2] ,
         \registers[656][1] , \registers[656][0] , \registers[655][7] ,
         \registers[655][6] , \registers[655][5] , \registers[655][4] ,
         \registers[655][3] , \registers[655][2] , \registers[655][1] ,
         \registers[655][0] , \registers[654][7] , \registers[654][6] ,
         \registers[654][5] , \registers[654][4] , \registers[654][3] ,
         \registers[654][2] , \registers[654][1] , \registers[654][0] ,
         \registers[653][7] , \registers[653][6] , \registers[653][5] ,
         \registers[653][4] , \registers[653][3] , \registers[653][2] ,
         \registers[653][1] , \registers[653][0] , \registers[652][7] ,
         \registers[652][6] , \registers[652][5] , \registers[652][4] ,
         \registers[652][3] , \registers[652][2] , \registers[652][1] ,
         \registers[652][0] , \registers[651][7] , \registers[651][6] ,
         \registers[651][5] , \registers[651][4] , \registers[651][3] ,
         \registers[651][2] , \registers[651][1] , \registers[651][0] ,
         \registers[650][7] , \registers[650][6] , \registers[650][5] ,
         \registers[650][4] , \registers[650][3] , \registers[650][2] ,
         \registers[650][1] , \registers[650][0] , \registers[649][7] ,
         \registers[649][6] , \registers[649][5] , \registers[649][4] ,
         \registers[649][3] , \registers[649][2] , \registers[649][1] ,
         \registers[649][0] , \registers[648][7] , \registers[648][6] ,
         \registers[648][5] , \registers[648][4] , \registers[648][3] ,
         \registers[648][2] , \registers[648][1] , \registers[648][0] ,
         \registers[647][7] , \registers[647][6] , \registers[647][5] ,
         \registers[647][4] , \registers[647][3] , \registers[647][2] ,
         \registers[647][1] , \registers[647][0] , \registers[646][7] ,
         \registers[646][6] , \registers[646][5] , \registers[646][4] ,
         \registers[646][3] , \registers[646][2] , \registers[646][1] ,
         \registers[646][0] , \registers[645][7] , \registers[645][6] ,
         \registers[645][5] , \registers[645][4] , \registers[645][3] ,
         \registers[645][2] , \registers[645][1] , \registers[645][0] ,
         \registers[644][7] , \registers[644][6] , \registers[644][5] ,
         \registers[644][4] , \registers[644][3] , \registers[644][2] ,
         \registers[644][1] , \registers[644][0] , \registers[643][7] ,
         \registers[643][6] , \registers[643][5] , \registers[643][4] ,
         \registers[643][3] , \registers[643][2] , \registers[643][1] ,
         \registers[643][0] , \registers[642][7] , \registers[642][6] ,
         \registers[642][5] , \registers[642][4] , \registers[642][3] ,
         \registers[642][2] , \registers[642][1] , \registers[642][0] ,
         \registers[641][7] , \registers[641][6] , \registers[641][5] ,
         \registers[641][4] , \registers[641][3] , \registers[641][2] ,
         \registers[641][1] , \registers[641][0] , \registers[640][7] ,
         \registers[640][6] , \registers[640][5] , \registers[640][4] ,
         \registers[640][3] , \registers[640][2] , \registers[640][1] ,
         \registers[640][0] , \registers[703][7] , \registers[703][6] ,
         \registers[703][5] , \registers[703][4] , \registers[703][3] ,
         \registers[703][2] , \registers[703][1] , \registers[703][0] ,
         \registers[702][7] , \registers[702][6] , \registers[702][5] ,
         \registers[702][4] , \registers[702][3] , \registers[702][2] ,
         \registers[702][1] , \registers[702][0] , \registers[701][7] ,
         \registers[701][6] , \registers[701][5] , \registers[701][4] ,
         \registers[701][3] , \registers[701][2] , \registers[701][1] ,
         \registers[701][0] , \registers[700][7] , \registers[700][6] ,
         \registers[700][5] , \registers[700][4] , \registers[700][3] ,
         \registers[700][2] , \registers[700][1] , \registers[700][0] ,
         \registers[699][7] , \registers[699][6] , \registers[699][5] ,
         \registers[699][4] , \registers[699][3] , \registers[699][2] ,
         \registers[699][1] , \registers[699][0] , \registers[698][7] ,
         \registers[698][6] , \registers[698][5] , \registers[698][4] ,
         \registers[698][3] , \registers[698][2] , \registers[698][1] ,
         \registers[698][0] , \registers[697][7] , \registers[697][6] ,
         \registers[697][5] , \registers[697][4] , \registers[697][3] ,
         \registers[697][2] , \registers[697][1] , \registers[697][0] ,
         \registers[696][7] , \registers[696][6] , \registers[696][5] ,
         \registers[696][4] , \registers[696][3] , \registers[696][2] ,
         \registers[696][1] , \registers[696][0] , \registers[695][7] ,
         \registers[695][6] , \registers[695][5] , \registers[695][4] ,
         \registers[695][3] , \registers[695][2] , \registers[695][1] ,
         \registers[695][0] , \registers[694][7] , \registers[694][6] ,
         \registers[694][5] , \registers[694][4] , \registers[694][3] ,
         \registers[694][2] , \registers[694][1] , \registers[694][0] ,
         \registers[693][7] , \registers[693][6] , \registers[693][5] ,
         \registers[693][4] , \registers[693][3] , \registers[693][2] ,
         \registers[693][1] , \registers[693][0] , \registers[692][7] ,
         \registers[692][6] , \registers[692][5] , \registers[692][4] ,
         \registers[692][3] , \registers[692][2] , \registers[692][1] ,
         \registers[692][0] , \registers[691][7] , \registers[691][6] ,
         \registers[691][5] , \registers[691][4] , \registers[691][3] ,
         \registers[691][2] , \registers[691][1] , \registers[691][0] ,
         \registers[690][7] , \registers[690][6] , \registers[690][5] ,
         \registers[690][4] , \registers[690][3] , \registers[690][2] ,
         \registers[690][1] , \registers[690][0] , \registers[689][7] ,
         \registers[689][6] , \registers[689][5] , \registers[689][4] ,
         \registers[689][3] , \registers[689][2] , \registers[689][1] ,
         \registers[689][0] , \registers[688][7] , \registers[688][6] ,
         \registers[688][5] , \registers[688][4] , \registers[688][3] ,
         \registers[688][2] , \registers[688][1] , \registers[688][0] ,
         \registers[687][7] , \registers[687][6] , \registers[687][5] ,
         \registers[687][4] , \registers[687][3] , \registers[687][2] ,
         \registers[687][1] , \registers[687][0] , \registers[686][7] ,
         \registers[686][6] , \registers[686][5] , \registers[686][4] ,
         \registers[686][3] , \registers[686][2] , \registers[686][1] ,
         \registers[686][0] , \registers[685][7] , \registers[685][6] ,
         \registers[685][5] , \registers[685][4] , \registers[685][3] ,
         \registers[685][2] , \registers[685][1] , \registers[685][0] ,
         \registers[684][7] , \registers[684][6] , \registers[684][5] ,
         \registers[684][4] , \registers[684][3] , \registers[684][2] ,
         \registers[684][1] , \registers[684][0] , \registers[683][7] ,
         \registers[683][6] , \registers[683][5] , \registers[683][4] ,
         \registers[683][3] , \registers[683][2] , \registers[683][1] ,
         \registers[683][0] , \registers[682][7] , \registers[682][6] ,
         \registers[682][5] , \registers[682][4] , \registers[682][3] ,
         \registers[682][2] , \registers[682][1] , \registers[682][0] ,
         \registers[681][7] , \registers[681][6] , \registers[681][5] ,
         \registers[681][4] , \registers[681][3] , \registers[681][2] ,
         \registers[681][1] , \registers[681][0] , \registers[680][7] ,
         \registers[680][6] , \registers[680][5] , \registers[680][4] ,
         \registers[680][3] , \registers[680][2] , \registers[680][1] ,
         \registers[680][0] , \registers[679][7] , \registers[679][6] ,
         \registers[679][5] , \registers[679][4] , \registers[679][3] ,
         \registers[679][2] , \registers[679][1] , \registers[679][0] ,
         \registers[678][7] , \registers[678][6] , \registers[678][5] ,
         \registers[678][4] , \registers[678][3] , \registers[678][2] ,
         \registers[678][1] , \registers[678][0] , \registers[677][7] ,
         \registers[677][6] , \registers[677][5] , \registers[677][4] ,
         \registers[677][3] , \registers[677][2] , \registers[677][1] ,
         \registers[677][0] , \registers[676][7] , \registers[676][6] ,
         \registers[676][5] , \registers[676][4] , \registers[676][3] ,
         \registers[676][2] , \registers[676][1] , \registers[676][0] ,
         \registers[675][7] , \registers[675][6] , \registers[675][5] ,
         \registers[675][4] , \registers[675][3] , \registers[675][2] ,
         \registers[675][1] , \registers[675][0] , \registers[674][7] ,
         \registers[674][6] , \registers[674][5] , \registers[674][4] ,
         \registers[674][3] , \registers[674][2] , \registers[674][1] ,
         \registers[674][0] , \registers[673][7] , \registers[673][6] ,
         \registers[673][5] , \registers[673][4] , \registers[673][3] ,
         \registers[673][2] , \registers[673][1] , \registers[673][0] ,
         \registers[672][7] , \registers[672][6] , \registers[672][5] ,
         \registers[672][4] , \registers[672][3] , \registers[672][2] ,
         \registers[672][1] , \registers[672][0] , \registers[735][7] ,
         \registers[735][6] , \registers[735][5] , \registers[735][4] ,
         \registers[735][3] , \registers[735][2] , \registers[735][1] ,
         \registers[735][0] , \registers[734][7] , \registers[734][6] ,
         \registers[734][5] , \registers[734][4] , \registers[734][3] ,
         \registers[734][2] , \registers[734][1] , \registers[734][0] ,
         \registers[733][7] , \registers[733][6] , \registers[733][5] ,
         \registers[733][4] , \registers[733][3] , \registers[733][2] ,
         \registers[733][1] , \registers[733][0] , \registers[732][7] ,
         \registers[732][6] , \registers[732][5] , \registers[732][4] ,
         \registers[732][3] , \registers[732][2] , \registers[732][1] ,
         \registers[732][0] , \registers[731][7] , \registers[731][6] ,
         \registers[731][5] , \registers[731][4] , \registers[731][3] ,
         \registers[731][2] , \registers[731][1] , \registers[731][0] ,
         \registers[730][7] , \registers[730][6] , \registers[730][5] ,
         \registers[730][4] , \registers[730][3] , \registers[730][2] ,
         \registers[730][1] , \registers[730][0] , \registers[729][7] ,
         \registers[729][6] , \registers[729][5] , \registers[729][4] ,
         \registers[729][3] , \registers[729][2] , \registers[729][1] ,
         \registers[729][0] , \registers[728][7] , \registers[728][6] ,
         \registers[728][5] , \registers[728][4] , \registers[728][3] ,
         \registers[728][2] , \registers[728][1] , \registers[728][0] ,
         \registers[727][7] , \registers[727][6] , \registers[727][5] ,
         \registers[727][4] , \registers[727][3] , \registers[727][2] ,
         \registers[727][1] , \registers[727][0] , \registers[726][7] ,
         \registers[726][6] , \registers[726][5] , \registers[726][4] ,
         \registers[726][3] , \registers[726][2] , \registers[726][1] ,
         \registers[726][0] , \registers[725][7] , \registers[725][6] ,
         \registers[725][5] , \registers[725][4] , \registers[725][3] ,
         \registers[725][2] , \registers[725][1] , \registers[725][0] ,
         \registers[724][7] , \registers[724][6] , \registers[724][5] ,
         \registers[724][4] , \registers[724][3] , \registers[724][2] ,
         \registers[724][1] , \registers[724][0] , \registers[723][7] ,
         \registers[723][6] , \registers[723][5] , \registers[723][4] ,
         \registers[723][3] , \registers[723][2] , \registers[723][1] ,
         \registers[723][0] , \registers[722][7] , \registers[722][6] ,
         \registers[722][5] , \registers[722][4] , \registers[722][3] ,
         \registers[722][2] , \registers[722][1] , \registers[722][0] ,
         \registers[721][7] , \registers[721][6] , \registers[721][5] ,
         \registers[721][4] , \registers[721][3] , \registers[721][2] ,
         \registers[721][1] , \registers[721][0] , \registers[720][7] ,
         \registers[720][6] , \registers[720][5] , \registers[720][4] ,
         \registers[720][3] , \registers[720][2] , \registers[720][1] ,
         \registers[720][0] , \registers[719][7] , \registers[719][6] ,
         \registers[719][5] , \registers[719][4] , \registers[719][3] ,
         \registers[719][2] , \registers[719][1] , \registers[719][0] ,
         \registers[718][7] , \registers[718][6] , \registers[718][5] ,
         \registers[718][4] , \registers[718][3] , \registers[718][2] ,
         \registers[718][1] , \registers[718][0] , \registers[717][7] ,
         \registers[717][6] , \registers[717][5] , \registers[717][4] ,
         \registers[717][3] , \registers[717][2] , \registers[717][1] ,
         \registers[717][0] , \registers[716][7] , \registers[716][6] ,
         \registers[716][5] , \registers[716][4] , \registers[716][3] ,
         \registers[716][2] , \registers[716][1] , \registers[716][0] ,
         \registers[715][7] , \registers[715][6] , \registers[715][5] ,
         \registers[715][4] , \registers[715][3] , \registers[715][2] ,
         \registers[715][1] , \registers[715][0] , \registers[714][7] ,
         \registers[714][6] , \registers[714][5] , \registers[714][4] ,
         \registers[714][3] , \registers[714][2] , \registers[714][1] ,
         \registers[714][0] , \registers[713][7] , \registers[713][6] ,
         \registers[713][5] , \registers[713][4] , \registers[713][3] ,
         \registers[713][2] , \registers[713][1] , \registers[713][0] ,
         \registers[712][7] , \registers[712][6] , \registers[712][5] ,
         \registers[712][4] , \registers[712][3] , \registers[712][2] ,
         \registers[712][1] , \registers[712][0] , \registers[711][7] ,
         \registers[711][6] , \registers[711][5] , \registers[711][4] ,
         \registers[711][3] , \registers[711][2] , \registers[711][1] ,
         \registers[711][0] , \registers[710][7] , \registers[710][6] ,
         \registers[710][5] , \registers[710][4] , \registers[710][3] ,
         \registers[710][2] , \registers[710][1] , \registers[710][0] ,
         \registers[709][7] , \registers[709][6] , \registers[709][5] ,
         \registers[709][4] , \registers[709][3] , \registers[709][2] ,
         \registers[709][1] , \registers[709][0] , \registers[708][7] ,
         \registers[708][6] , \registers[708][5] , \registers[708][4] ,
         \registers[708][3] , \registers[708][2] , \registers[708][1] ,
         \registers[708][0] , \registers[707][7] , \registers[707][6] ,
         \registers[707][5] , \registers[707][4] , \registers[707][3] ,
         \registers[707][2] , \registers[707][1] , \registers[707][0] ,
         \registers[706][7] , \registers[706][6] , \registers[706][5] ,
         \registers[706][4] , \registers[706][3] , \registers[706][2] ,
         \registers[706][1] , \registers[706][0] , \registers[705][7] ,
         \registers[705][6] , \registers[705][5] , \registers[705][4] ,
         \registers[705][3] , \registers[705][2] , \registers[705][1] ,
         \registers[705][0] , \registers[704][7] , \registers[704][6] ,
         \registers[704][5] , \registers[704][4] , \registers[704][3] ,
         \registers[704][2] , \registers[704][1] , \registers[704][0] ,
         \registers[767][7] , \registers[767][6] , \registers[767][5] ,
         \registers[767][4] , \registers[767][3] , \registers[767][2] ,
         \registers[767][1] , \registers[767][0] , \registers[766][7] ,
         \registers[766][6] , \registers[766][5] , \registers[766][4] ,
         \registers[766][3] , \registers[766][2] , \registers[766][1] ,
         \registers[766][0] , \registers[765][7] , \registers[765][6] ,
         \registers[765][5] , \registers[765][4] , \registers[765][3] ,
         \registers[765][2] , \registers[765][1] , \registers[765][0] ,
         \registers[764][7] , \registers[764][6] , \registers[764][5] ,
         \registers[764][4] , \registers[764][3] , \registers[764][2] ,
         \registers[764][1] , \registers[764][0] , \registers[763][7] ,
         \registers[763][6] , \registers[763][5] , \registers[763][4] ,
         \registers[763][3] , \registers[763][2] , \registers[763][1] ,
         \registers[763][0] , \registers[762][7] , \registers[762][6] ,
         \registers[762][5] , \registers[762][4] , \registers[762][3] ,
         \registers[762][2] , \registers[762][1] , \registers[762][0] ,
         \registers[761][7] , \registers[761][6] , \registers[761][5] ,
         \registers[761][4] , \registers[761][3] , \registers[761][2] ,
         \registers[761][1] , \registers[761][0] , \registers[760][7] ,
         \registers[760][6] , \registers[760][5] , \registers[760][4] ,
         \registers[760][3] , \registers[760][2] , \registers[760][1] ,
         \registers[760][0] , \registers[759][7] , \registers[759][6] ,
         \registers[759][5] , \registers[759][4] , \registers[759][3] ,
         \registers[759][2] , \registers[759][1] , \registers[759][0] ,
         \registers[758][7] , \registers[758][6] , \registers[758][5] ,
         \registers[758][4] , \registers[758][3] , \registers[758][2] ,
         \registers[758][1] , \registers[758][0] , \registers[757][7] ,
         \registers[757][6] , \registers[757][5] , \registers[757][4] ,
         \registers[757][3] , \registers[757][2] , \registers[757][1] ,
         \registers[757][0] , \registers[756][7] , \registers[756][6] ,
         \registers[756][5] , \registers[756][4] , \registers[756][3] ,
         \registers[756][2] , \registers[756][1] , \registers[756][0] ,
         \registers[755][7] , \registers[755][6] , \registers[755][5] ,
         \registers[755][4] , \registers[755][3] , \registers[755][2] ,
         \registers[755][1] , \registers[755][0] , \registers[754][7] ,
         \registers[754][6] , \registers[754][5] , \registers[754][4] ,
         \registers[754][3] , \registers[754][2] , \registers[754][1] ,
         \registers[754][0] , \registers[753][7] , \registers[753][6] ,
         \registers[753][5] , \registers[753][4] , \registers[753][3] ,
         \registers[753][2] , \registers[753][1] , \registers[753][0] ,
         \registers[752][7] , \registers[752][6] , \registers[752][5] ,
         \registers[752][4] , \registers[752][3] , \registers[752][2] ,
         \registers[752][1] , \registers[752][0] , \registers[751][7] ,
         \registers[751][6] , \registers[751][5] , \registers[751][4] ,
         \registers[751][3] , \registers[751][2] , \registers[751][1] ,
         \registers[751][0] , \registers[750][7] , \registers[750][6] ,
         \registers[750][5] , \registers[750][4] , \registers[750][3] ,
         \registers[750][2] , \registers[750][1] , \registers[750][0] ,
         \registers[749][7] , \registers[749][6] , \registers[749][5] ,
         \registers[749][4] , \registers[749][3] , \registers[749][2] ,
         \registers[749][1] , \registers[749][0] , \registers[748][7] ,
         \registers[748][6] , \registers[748][5] , \registers[748][4] ,
         \registers[748][3] , \registers[748][2] , \registers[748][1] ,
         \registers[748][0] , \registers[747][7] , \registers[747][6] ,
         \registers[747][5] , \registers[747][4] , \registers[747][3] ,
         \registers[747][2] , \registers[747][1] , \registers[747][0] ,
         \registers[746][7] , \registers[746][6] , \registers[746][5] ,
         \registers[746][4] , \registers[746][3] , \registers[746][2] ,
         \registers[746][1] , \registers[746][0] , \registers[745][7] ,
         \registers[745][6] , \registers[745][5] , \registers[745][4] ,
         \registers[745][3] , \registers[745][2] , \registers[745][1] ,
         \registers[745][0] , \registers[744][7] , \registers[744][6] ,
         \registers[744][5] , \registers[744][4] , \registers[744][3] ,
         \registers[744][2] , \registers[744][1] , \registers[744][0] ,
         \registers[743][7] , \registers[743][6] , \registers[743][5] ,
         \registers[743][4] , \registers[743][3] , \registers[743][2] ,
         \registers[743][1] , \registers[743][0] , \registers[742][7] ,
         \registers[742][6] , \registers[742][5] , \registers[742][4] ,
         \registers[742][3] , \registers[742][2] , \registers[742][1] ,
         \registers[742][0] , \registers[741][7] , \registers[741][6] ,
         \registers[741][5] , \registers[741][4] , \registers[741][3] ,
         \registers[741][2] , \registers[741][1] , \registers[741][0] ,
         \registers[740][7] , \registers[740][6] , \registers[740][5] ,
         \registers[740][4] , \registers[740][3] , \registers[740][2] ,
         \registers[740][1] , \registers[740][0] , \registers[739][7] ,
         \registers[739][6] , \registers[739][5] , \registers[739][4] ,
         \registers[739][3] , \registers[739][2] , \registers[739][1] ,
         \registers[739][0] , \registers[738][7] , \registers[738][6] ,
         \registers[738][5] , \registers[738][4] , \registers[738][3] ,
         \registers[738][2] , \registers[738][1] , \registers[738][0] ,
         \registers[737][7] , \registers[737][6] , \registers[737][5] ,
         \registers[737][4] , \registers[737][3] , \registers[737][2] ,
         \registers[737][1] , \registers[737][0] , \registers[736][7] ,
         \registers[736][6] , \registers[736][5] , \registers[736][4] ,
         \registers[736][3] , \registers[736][2] , \registers[736][1] ,
         \registers[736][0] , \registers[799][7] , \registers[799][6] ,
         \registers[799][5] , \registers[799][4] , \registers[799][3] ,
         \registers[799][2] , \registers[799][1] , \registers[799][0] ,
         \registers[798][7] , \registers[798][6] , \registers[798][5] ,
         \registers[798][4] , \registers[798][3] , \registers[798][2] ,
         \registers[798][1] , \registers[798][0] , \registers[797][7] ,
         \registers[797][6] , \registers[797][5] , \registers[797][4] ,
         \registers[797][3] , \registers[797][2] , \registers[797][1] ,
         \registers[797][0] , \registers[796][7] , \registers[796][6] ,
         \registers[796][5] , \registers[796][4] , \registers[796][3] ,
         \registers[796][2] , \registers[796][1] , \registers[796][0] ,
         \registers[795][7] , \registers[795][6] , \registers[795][5] ,
         \registers[795][4] , \registers[795][3] , \registers[795][2] ,
         \registers[795][1] , \registers[795][0] , \registers[794][7] ,
         \registers[794][6] , \registers[794][5] , \registers[794][4] ,
         \registers[794][3] , \registers[794][2] , \registers[794][1] ,
         \registers[794][0] , \registers[793][7] , \registers[793][6] ,
         \registers[793][5] , \registers[793][4] , \registers[793][3] ,
         \registers[793][2] , \registers[793][1] , \registers[793][0] ,
         \registers[792][7] , \registers[792][6] , \registers[792][5] ,
         \registers[792][4] , \registers[792][3] , \registers[792][2] ,
         \registers[792][1] , \registers[792][0] , \registers[791][7] ,
         \registers[791][6] , \registers[791][5] , \registers[791][4] ,
         \registers[791][3] , \registers[791][2] , \registers[791][1] ,
         \registers[791][0] , \registers[790][7] , \registers[790][6] ,
         \registers[790][5] , \registers[790][4] , \registers[790][3] ,
         \registers[790][2] , \registers[790][1] , \registers[790][0] ,
         \registers[789][7] , \registers[789][6] , \registers[789][5] ,
         \registers[789][4] , \registers[789][3] , \registers[789][2] ,
         \registers[789][1] , \registers[789][0] , \registers[788][7] ,
         \registers[788][6] , \registers[788][5] , \registers[788][4] ,
         \registers[788][3] , \registers[788][2] , \registers[788][1] ,
         \registers[788][0] , \registers[787][7] , \registers[787][6] ,
         \registers[787][5] , \registers[787][4] , \registers[787][3] ,
         \registers[787][2] , \registers[787][1] , \registers[787][0] ,
         \registers[786][7] , \registers[786][6] , \registers[786][5] ,
         \registers[786][4] , \registers[786][3] , \registers[786][2] ,
         \registers[786][1] , \registers[786][0] , \registers[785][7] ,
         \registers[785][6] , \registers[785][5] , \registers[785][4] ,
         \registers[785][3] , \registers[785][2] , \registers[785][1] ,
         \registers[785][0] , \registers[784][7] , \registers[784][6] ,
         \registers[784][5] , \registers[784][4] , \registers[784][3] ,
         \registers[784][2] , \registers[784][1] , \registers[784][0] ,
         \registers[783][7] , \registers[783][6] , \registers[783][5] ,
         \registers[783][4] , \registers[783][3] , \registers[783][2] ,
         \registers[783][1] , \registers[783][0] , \registers[782][7] ,
         \registers[782][6] , \registers[782][5] , \registers[782][4] ,
         \registers[782][3] , \registers[782][2] , \registers[782][1] ,
         \registers[782][0] , \registers[781][7] , \registers[781][6] ,
         \registers[781][5] , \registers[781][4] , \registers[781][3] ,
         \registers[781][2] , \registers[781][1] , \registers[781][0] ,
         \registers[780][7] , \registers[780][6] , \registers[780][5] ,
         \registers[780][4] , \registers[780][3] , \registers[780][2] ,
         \registers[780][1] , \registers[780][0] , \registers[779][7] ,
         \registers[779][6] , \registers[779][5] , \registers[779][4] ,
         \registers[779][3] , \registers[779][2] , \registers[779][1] ,
         \registers[779][0] , \registers[778][7] , \registers[778][6] ,
         \registers[778][5] , \registers[778][4] , \registers[778][3] ,
         \registers[778][2] , \registers[778][1] , \registers[778][0] ,
         \registers[777][7] , \registers[777][6] , \registers[777][5] ,
         \registers[777][4] , \registers[777][3] , \registers[777][2] ,
         \registers[777][1] , \registers[777][0] , \registers[776][7] ,
         \registers[776][6] , \registers[776][5] , \registers[776][4] ,
         \registers[776][3] , \registers[776][2] , \registers[776][1] ,
         \registers[776][0] , \registers[775][7] , \registers[775][6] ,
         \registers[775][5] , \registers[775][4] , \registers[775][3] ,
         \registers[775][2] , \registers[775][1] , \registers[775][0] ,
         \registers[774][7] , \registers[774][6] , \registers[774][5] ,
         \registers[774][4] , \registers[774][3] , \registers[774][2] ,
         \registers[774][1] , \registers[774][0] , \registers[773][7] ,
         \registers[773][6] , \registers[773][5] , \registers[773][4] ,
         \registers[773][3] , \registers[773][2] , \registers[773][1] ,
         \registers[773][0] , \registers[772][7] , \registers[772][6] ,
         \registers[772][5] , \registers[772][4] , \registers[772][3] ,
         \registers[772][2] , \registers[772][1] , \registers[772][0] ,
         \registers[771][7] , \registers[771][6] , \registers[771][5] ,
         \registers[771][4] , \registers[771][3] , \registers[771][2] ,
         \registers[771][1] , \registers[771][0] , \registers[770][7] ,
         \registers[770][6] , \registers[770][5] , \registers[770][4] ,
         \registers[770][3] , \registers[770][2] , \registers[770][1] ,
         \registers[770][0] , \registers[769][7] , \registers[769][6] ,
         \registers[769][5] , \registers[769][4] , \registers[769][3] ,
         \registers[769][2] , \registers[769][1] , \registers[769][0] ,
         \registers[768][7] , \registers[768][6] , \registers[768][5] ,
         \registers[768][4] , \registers[768][3] , \registers[768][2] ,
         \registers[768][1] , \registers[768][0] , \registers[831][7] ,
         \registers[831][6] , \registers[831][5] , \registers[831][4] ,
         \registers[831][3] , \registers[831][2] , \registers[831][1] ,
         \registers[831][0] , \registers[830][7] , \registers[830][6] ,
         \registers[830][5] , \registers[830][4] , \registers[830][3] ,
         \registers[830][2] , \registers[830][1] , \registers[830][0] ,
         \registers[829][7] , \registers[829][6] , \registers[829][5] ,
         \registers[829][4] , \registers[829][3] , \registers[829][2] ,
         \registers[829][1] , \registers[829][0] , \registers[828][7] ,
         \registers[828][6] , \registers[828][5] , \registers[828][4] ,
         \registers[828][3] , \registers[828][2] , \registers[828][1] ,
         \registers[828][0] , \registers[827][7] , \registers[827][6] ,
         \registers[827][5] , \registers[827][4] , \registers[827][3] ,
         \registers[827][2] , \registers[827][1] , \registers[827][0] ,
         \registers[826][7] , \registers[826][6] , \registers[826][5] ,
         \registers[826][4] , \registers[826][3] , \registers[826][2] ,
         \registers[826][1] , \registers[826][0] , \registers[825][7] ,
         \registers[825][6] , \registers[825][5] , \registers[825][4] ,
         \registers[825][3] , \registers[825][2] , \registers[825][1] ,
         \registers[825][0] , \registers[824][7] , \registers[824][6] ,
         \registers[824][5] , \registers[824][4] , \registers[824][3] ,
         \registers[824][2] , \registers[824][1] , \registers[824][0] ,
         \registers[823][7] , \registers[823][6] , \registers[823][5] ,
         \registers[823][4] , \registers[823][3] , \registers[823][2] ,
         \registers[823][1] , \registers[823][0] , \registers[822][7] ,
         \registers[822][6] , \registers[822][5] , \registers[822][4] ,
         \registers[822][3] , \registers[822][2] , \registers[822][1] ,
         \registers[822][0] , \registers[821][7] , \registers[821][6] ,
         \registers[821][5] , \registers[821][4] , \registers[821][3] ,
         \registers[821][2] , \registers[821][1] , \registers[821][0] ,
         \registers[820][7] , \registers[820][6] , \registers[820][5] ,
         \registers[820][4] , \registers[820][3] , \registers[820][2] ,
         \registers[820][1] , \registers[820][0] , \registers[819][7] ,
         \registers[819][6] , \registers[819][5] , \registers[819][4] ,
         \registers[819][3] , \registers[819][2] , \registers[819][1] ,
         \registers[819][0] , \registers[818][7] , \registers[818][6] ,
         \registers[818][5] , \registers[818][4] , \registers[818][3] ,
         \registers[818][2] , \registers[818][1] , \registers[818][0] ,
         \registers[817][7] , \registers[817][6] , \registers[817][5] ,
         \registers[817][4] , \registers[817][3] , \registers[817][2] ,
         \registers[817][1] , \registers[817][0] , \registers[816][7] ,
         \registers[816][6] , \registers[816][5] , \registers[816][4] ,
         \registers[816][3] , \registers[816][2] , \registers[816][1] ,
         \registers[816][0] , \registers[815][7] , \registers[815][6] ,
         \registers[815][5] , \registers[815][4] , \registers[815][3] ,
         \registers[815][2] , \registers[815][1] , \registers[815][0] ,
         \registers[814][7] , \registers[814][6] , \registers[814][5] ,
         \registers[814][4] , \registers[814][3] , \registers[814][2] ,
         \registers[814][1] , \registers[814][0] , \registers[813][7] ,
         \registers[813][6] , \registers[813][5] , \registers[813][4] ,
         \registers[813][3] , \registers[813][2] , \registers[813][1] ,
         \registers[813][0] , \registers[812][7] , \registers[812][6] ,
         \registers[812][5] , \registers[812][4] , \registers[812][3] ,
         \registers[812][2] , \registers[812][1] , \registers[812][0] ,
         \registers[811][7] , \registers[811][6] , \registers[811][5] ,
         \registers[811][4] , \registers[811][3] , \registers[811][2] ,
         \registers[811][1] , \registers[811][0] , \registers[810][7] ,
         \registers[810][6] , \registers[810][5] , \registers[810][4] ,
         \registers[810][3] , \registers[810][2] , \registers[810][1] ,
         \registers[810][0] , \registers[809][7] , \registers[809][6] ,
         \registers[809][5] , \registers[809][4] , \registers[809][3] ,
         \registers[809][2] , \registers[809][1] , \registers[809][0] ,
         \registers[808][7] , \registers[808][6] , \registers[808][5] ,
         \registers[808][4] , \registers[808][3] , \registers[808][2] ,
         \registers[808][1] , \registers[808][0] , \registers[807][7] ,
         \registers[807][6] , \registers[807][5] , \registers[807][4] ,
         \registers[807][3] , \registers[807][2] , \registers[807][1] ,
         \registers[807][0] , \registers[806][7] , \registers[806][6] ,
         \registers[806][5] , \registers[806][4] , \registers[806][3] ,
         \registers[806][2] , \registers[806][1] , \registers[806][0] ,
         \registers[805][7] , \registers[805][6] , \registers[805][5] ,
         \registers[805][4] , \registers[805][3] , \registers[805][2] ,
         \registers[805][1] , \registers[805][0] , \registers[804][7] ,
         \registers[804][6] , \registers[804][5] , \registers[804][4] ,
         \registers[804][3] , \registers[804][2] , \registers[804][1] ,
         \registers[804][0] , \registers[803][7] , \registers[803][6] ,
         \registers[803][5] , \registers[803][4] , \registers[803][3] ,
         \registers[803][2] , \registers[803][1] , \registers[803][0] ,
         \registers[802][7] , \registers[802][6] , \registers[802][5] ,
         \registers[802][4] , \registers[802][3] , \registers[802][2] ,
         \registers[802][1] , \registers[802][0] , \registers[801][7] ,
         \registers[801][6] , \registers[801][5] , \registers[801][4] ,
         \registers[801][3] , \registers[801][2] , \registers[801][1] ,
         \registers[801][0] , \registers[800][7] , \registers[800][6] ,
         \registers[800][5] , \registers[800][4] , \registers[800][3] ,
         \registers[800][2] , \registers[800][1] , \registers[800][0] ,
         \registers[863][7] , \registers[863][6] , \registers[863][5] ,
         \registers[863][4] , \registers[863][3] , \registers[863][2] ,
         \registers[863][1] , \registers[863][0] , \registers[862][7] ,
         \registers[862][6] , \registers[862][5] , \registers[862][4] ,
         \registers[862][3] , \registers[862][2] , \registers[862][1] ,
         \registers[862][0] , \registers[861][7] , \registers[861][6] ,
         \registers[861][5] , \registers[861][4] , \registers[861][3] ,
         \registers[861][2] , \registers[861][1] , \registers[861][0] ,
         \registers[860][7] , \registers[860][6] , \registers[860][5] ,
         \registers[860][4] , \registers[860][3] , \registers[860][2] ,
         \registers[860][1] , \registers[860][0] , \registers[859][7] ,
         \registers[859][6] , \registers[859][5] , \registers[859][4] ,
         \registers[859][3] , \registers[859][2] , \registers[859][1] ,
         \registers[859][0] , \registers[858][7] , \registers[858][6] ,
         \registers[858][5] , \registers[858][4] , \registers[858][3] ,
         \registers[858][2] , \registers[858][1] , \registers[858][0] ,
         \registers[857][7] , \registers[857][6] , \registers[857][5] ,
         \registers[857][4] , \registers[857][3] , \registers[857][2] ,
         \registers[857][1] , \registers[857][0] , \registers[856][7] ,
         \registers[856][6] , \registers[856][5] , \registers[856][4] ,
         \registers[856][3] , \registers[856][2] , \registers[856][1] ,
         \registers[856][0] , \registers[855][7] , \registers[855][6] ,
         \registers[855][5] , \registers[855][4] , \registers[855][3] ,
         \registers[855][2] , \registers[855][1] , \registers[855][0] ,
         \registers[854][7] , \registers[854][6] , \registers[854][5] ,
         \registers[854][4] , \registers[854][3] , \registers[854][2] ,
         \registers[854][1] , \registers[854][0] , \registers[853][7] ,
         \registers[853][6] , \registers[853][5] , \registers[853][4] ,
         \registers[853][3] , \registers[853][2] , \registers[853][1] ,
         \registers[853][0] , \registers[852][7] , \registers[852][6] ,
         \registers[852][5] , \registers[852][4] , \registers[852][3] ,
         \registers[852][2] , \registers[852][1] , \registers[852][0] ,
         \registers[851][7] , \registers[851][6] , \registers[851][5] ,
         \registers[851][4] , \registers[851][3] , \registers[851][2] ,
         \registers[851][1] , \registers[851][0] , \registers[850][7] ,
         \registers[850][6] , \registers[850][5] , \registers[850][4] ,
         \registers[850][3] , \registers[850][2] , \registers[850][1] ,
         \registers[850][0] , \registers[849][7] , \registers[849][6] ,
         \registers[849][5] , \registers[849][4] , \registers[849][3] ,
         \registers[849][2] , \registers[849][1] , \registers[849][0] ,
         \registers[848][7] , \registers[848][6] , \registers[848][5] ,
         \registers[848][4] , \registers[848][3] , \registers[848][2] ,
         \registers[848][1] , \registers[848][0] , \registers[847][7] ,
         \registers[847][6] , \registers[847][5] , \registers[847][4] ,
         \registers[847][3] , \registers[847][2] , \registers[847][1] ,
         \registers[847][0] , \registers[846][7] , \registers[846][6] ,
         \registers[846][5] , \registers[846][4] , \registers[846][3] ,
         \registers[846][2] , \registers[846][1] , \registers[846][0] ,
         \registers[845][7] , \registers[845][6] , \registers[845][5] ,
         \registers[845][4] , \registers[845][3] , \registers[845][2] ,
         \registers[845][1] , \registers[845][0] , \registers[844][7] ,
         \registers[844][6] , \registers[844][5] , \registers[844][4] ,
         \registers[844][3] , \registers[844][2] , \registers[844][1] ,
         \registers[844][0] , \registers[843][7] , \registers[843][6] ,
         \registers[843][5] , \registers[843][4] , \registers[843][3] ,
         \registers[843][2] , \registers[843][1] , \registers[843][0] ,
         \registers[842][7] , \registers[842][6] , \registers[842][5] ,
         \registers[842][4] , \registers[842][3] , \registers[842][2] ,
         \registers[842][1] , \registers[842][0] , \registers[841][7] ,
         \registers[841][6] , \registers[841][5] , \registers[841][4] ,
         \registers[841][3] , \registers[841][2] , \registers[841][1] ,
         \registers[841][0] , \registers[840][7] , \registers[840][6] ,
         \registers[840][5] , \registers[840][4] , \registers[840][3] ,
         \registers[840][2] , \registers[840][1] , \registers[840][0] ,
         \registers[839][7] , \registers[839][6] , \registers[839][5] ,
         \registers[839][4] , \registers[839][3] , \registers[839][2] ,
         \registers[839][1] , \registers[839][0] , \registers[838][7] ,
         \registers[838][6] , \registers[838][5] , \registers[838][4] ,
         \registers[838][3] , \registers[838][2] , \registers[838][1] ,
         \registers[838][0] , \registers[837][7] , \registers[837][6] ,
         \registers[837][5] , \registers[837][4] , \registers[837][3] ,
         \registers[837][2] , \registers[837][1] , \registers[837][0] ,
         \registers[836][7] , \registers[836][6] , \registers[836][5] ,
         \registers[836][4] , \registers[836][3] , \registers[836][2] ,
         \registers[836][1] , \registers[836][0] , \registers[835][7] ,
         \registers[835][6] , \registers[835][5] , \registers[835][4] ,
         \registers[835][3] , \registers[835][2] , \registers[835][1] ,
         \registers[835][0] , \registers[834][7] , \registers[834][6] ,
         \registers[834][5] , \registers[834][4] , \registers[834][3] ,
         \registers[834][2] , \registers[834][1] , \registers[834][0] ,
         \registers[833][7] , \registers[833][6] , \registers[833][5] ,
         \registers[833][4] , \registers[833][3] , \registers[833][2] ,
         \registers[833][1] , \registers[833][0] , \registers[832][7] ,
         \registers[832][6] , \registers[832][5] , \registers[832][4] ,
         \registers[832][3] , \registers[832][2] , \registers[832][1] ,
         \registers[832][0] , \registers[895][7] , \registers[895][6] ,
         \registers[895][5] , \registers[895][4] , \registers[895][3] ,
         \registers[895][2] , \registers[895][1] , \registers[895][0] ,
         \registers[894][7] , \registers[894][6] , \registers[894][5] ,
         \registers[894][4] , \registers[894][3] , \registers[894][2] ,
         \registers[894][1] , \registers[894][0] , \registers[893][7] ,
         \registers[893][6] , \registers[893][5] , \registers[893][4] ,
         \registers[893][3] , \registers[893][2] , \registers[893][1] ,
         \registers[893][0] , \registers[892][7] , \registers[892][6] ,
         \registers[892][5] , \registers[892][4] , \registers[892][3] ,
         \registers[892][2] , \registers[892][1] , \registers[892][0] ,
         \registers[891][7] , \registers[891][6] , \registers[891][5] ,
         \registers[891][4] , \registers[891][3] , \registers[891][2] ,
         \registers[891][1] , \registers[891][0] , \registers[890][7] ,
         \registers[890][6] , \registers[890][5] , \registers[890][4] ,
         \registers[890][3] , \registers[890][2] , \registers[890][1] ,
         \registers[890][0] , \registers[889][7] , \registers[889][6] ,
         \registers[889][5] , \registers[889][4] , \registers[889][3] ,
         \registers[889][2] , \registers[889][1] , \registers[889][0] ,
         \registers[888][7] , \registers[888][6] , \registers[888][5] ,
         \registers[888][4] , \registers[888][3] , \registers[888][2] ,
         \registers[888][1] , \registers[888][0] , \registers[887][7] ,
         \registers[887][6] , \registers[887][5] , \registers[887][4] ,
         \registers[887][3] , \registers[887][2] , \registers[887][1] ,
         \registers[887][0] , \registers[886][7] , \registers[886][6] ,
         \registers[886][5] , \registers[886][4] , \registers[886][3] ,
         \registers[886][2] , \registers[886][1] , \registers[886][0] ,
         \registers[885][7] , \registers[885][6] , \registers[885][5] ,
         \registers[885][4] , \registers[885][3] , \registers[885][2] ,
         \registers[885][1] , \registers[885][0] , \registers[884][7] ,
         \registers[884][6] , \registers[884][5] , \registers[884][4] ,
         \registers[884][3] , \registers[884][2] , \registers[884][1] ,
         \registers[884][0] , \registers[883][7] , \registers[883][6] ,
         \registers[883][5] , \registers[883][4] , \registers[883][3] ,
         \registers[883][2] , \registers[883][1] , \registers[883][0] ,
         \registers[882][7] , \registers[882][6] , \registers[882][5] ,
         \registers[882][4] , \registers[882][3] , \registers[882][2] ,
         \registers[882][1] , \registers[882][0] , \registers[881][7] ,
         \registers[881][6] , \registers[881][5] , \registers[881][4] ,
         \registers[881][3] , \registers[881][2] , \registers[881][1] ,
         \registers[881][0] , \registers[880][7] , \registers[880][6] ,
         \registers[880][5] , \registers[880][4] , \registers[880][3] ,
         \registers[880][2] , \registers[880][1] , \registers[880][0] ,
         \registers[879][7] , \registers[879][6] , \registers[879][5] ,
         \registers[879][4] , \registers[879][3] , \registers[879][2] ,
         \registers[879][1] , \registers[879][0] , \registers[878][7] ,
         \registers[878][6] , \registers[878][5] , \registers[878][4] ,
         \registers[878][3] , \registers[878][2] , \registers[878][1] ,
         \registers[878][0] , \registers[877][7] , \registers[877][6] ,
         \registers[877][5] , \registers[877][4] , \registers[877][3] ,
         \registers[877][2] , \registers[877][1] , \registers[877][0] ,
         \registers[876][7] , \registers[876][6] , \registers[876][5] ,
         \registers[876][4] , \registers[876][3] , \registers[876][2] ,
         \registers[876][1] , \registers[876][0] , \registers[875][7] ,
         \registers[875][6] , \registers[875][5] , \registers[875][4] ,
         \registers[875][3] , \registers[875][2] , \registers[875][1] ,
         \registers[875][0] , \registers[874][7] , \registers[874][6] ,
         \registers[874][5] , \registers[874][4] , \registers[874][3] ,
         \registers[874][2] , \registers[874][1] , \registers[874][0] ,
         \registers[873][7] , \registers[873][6] , \registers[873][5] ,
         \registers[873][4] , \registers[873][3] , \registers[873][2] ,
         \registers[873][1] , \registers[873][0] , \registers[872][7] ,
         \registers[872][6] , \registers[872][5] , \registers[872][4] ,
         \registers[872][3] , \registers[872][2] , \registers[872][1] ,
         \registers[872][0] , \registers[871][7] , \registers[871][6] ,
         \registers[871][5] , \registers[871][4] , \registers[871][3] ,
         \registers[871][2] , \registers[871][1] , \registers[871][0] ,
         \registers[870][7] , \registers[870][6] , \registers[870][5] ,
         \registers[870][4] , \registers[870][3] , \registers[870][2] ,
         \registers[870][1] , \registers[870][0] , \registers[869][7] ,
         \registers[869][6] , \registers[869][5] , \registers[869][4] ,
         \registers[869][3] , \registers[869][2] , \registers[869][1] ,
         \registers[869][0] , \registers[868][7] , \registers[868][6] ,
         \registers[868][5] , \registers[868][4] , \registers[868][3] ,
         \registers[868][2] , \registers[868][1] , \registers[868][0] ,
         \registers[867][7] , \registers[867][6] , \registers[867][5] ,
         \registers[867][4] , \registers[867][3] , \registers[867][2] ,
         \registers[867][1] , \registers[867][0] , \registers[866][7] ,
         \registers[866][6] , \registers[866][5] , \registers[866][4] ,
         \registers[866][3] , \registers[866][2] , \registers[866][1] ,
         \registers[866][0] , \registers[865][7] , \registers[865][6] ,
         \registers[865][5] , \registers[865][4] , \registers[865][3] ,
         \registers[865][2] , \registers[865][1] , \registers[865][0] ,
         \registers[864][7] , \registers[864][6] , \registers[864][5] ,
         \registers[864][4] , \registers[864][3] , \registers[864][2] ,
         \registers[864][1] , \registers[864][0] , \registers[927][7] ,
         \registers[927][6] , \registers[927][5] , \registers[927][4] ,
         \registers[927][3] , \registers[927][2] , \registers[927][1] ,
         \registers[927][0] , \registers[926][7] , \registers[926][6] ,
         \registers[926][5] , \registers[926][4] , \registers[926][3] ,
         \registers[926][2] , \registers[926][1] , \registers[926][0] ,
         \registers[925][7] , \registers[925][6] , \registers[925][5] ,
         \registers[925][4] , \registers[925][3] , \registers[925][2] ,
         \registers[925][1] , \registers[925][0] , \registers[924][7] ,
         \registers[924][6] , \registers[924][5] , \registers[924][4] ,
         \registers[924][3] , \registers[924][2] , \registers[924][1] ,
         \registers[924][0] , \registers[923][7] , \registers[923][6] ,
         \registers[923][5] , \registers[923][4] , \registers[923][3] ,
         \registers[923][2] , \registers[923][1] , \registers[923][0] ,
         \registers[922][7] , \registers[922][6] , \registers[922][5] ,
         \registers[922][4] , \registers[922][3] , \registers[922][2] ,
         \registers[922][1] , \registers[922][0] , \registers[921][7] ,
         \registers[921][6] , \registers[921][5] , \registers[921][4] ,
         \registers[921][3] , \registers[921][2] , \registers[921][1] ,
         \registers[921][0] , \registers[920][7] , \registers[920][6] ,
         \registers[920][5] , \registers[920][4] , \registers[920][3] ,
         \registers[920][2] , \registers[920][1] , \registers[920][0] ,
         \registers[919][7] , \registers[919][6] , \registers[919][5] ,
         \registers[919][4] , \registers[919][3] , \registers[919][2] ,
         \registers[919][1] , \registers[919][0] , \registers[918][7] ,
         \registers[918][6] , \registers[918][5] , \registers[918][4] ,
         \registers[918][3] , \registers[918][2] , \registers[918][1] ,
         \registers[918][0] , \registers[917][7] , \registers[917][6] ,
         \registers[917][5] , \registers[917][4] , \registers[917][3] ,
         \registers[917][2] , \registers[917][1] , \registers[917][0] ,
         \registers[916][7] , \registers[916][6] , \registers[916][5] ,
         \registers[916][4] , \registers[916][3] , \registers[916][2] ,
         \registers[916][1] , \registers[916][0] , \registers[915][7] ,
         \registers[915][6] , \registers[915][5] , \registers[915][4] ,
         \registers[915][3] , \registers[915][2] , \registers[915][1] ,
         \registers[915][0] , \registers[914][7] , \registers[914][6] ,
         \registers[914][5] , \registers[914][4] , \registers[914][3] ,
         \registers[914][2] , \registers[914][1] , \registers[914][0] ,
         \registers[913][7] , \registers[913][6] , \registers[913][5] ,
         \registers[913][4] , \registers[913][3] , \registers[913][2] ,
         \registers[913][1] , \registers[913][0] , \registers[912][7] ,
         \registers[912][6] , \registers[912][5] , \registers[912][4] ,
         \registers[912][3] , \registers[912][2] , \registers[912][1] ,
         \registers[912][0] , \registers[911][7] , \registers[911][6] ,
         \registers[911][5] , \registers[911][4] , \registers[911][3] ,
         \registers[911][2] , \registers[911][1] , \registers[911][0] ,
         \registers[910][7] , \registers[910][6] , \registers[910][5] ,
         \registers[910][4] , \registers[910][3] , \registers[910][2] ,
         \registers[910][1] , \registers[910][0] , \registers[909][7] ,
         \registers[909][6] , \registers[909][5] , \registers[909][4] ,
         \registers[909][3] , \registers[909][2] , \registers[909][1] ,
         \registers[909][0] , \registers[908][7] , \registers[908][6] ,
         \registers[908][5] , \registers[908][4] , \registers[908][3] ,
         \registers[908][2] , \registers[908][1] , \registers[908][0] ,
         \registers[907][7] , \registers[907][6] , \registers[907][5] ,
         \registers[907][4] , \registers[907][3] , \registers[907][2] ,
         \registers[907][1] , \registers[907][0] , \registers[906][7] ,
         \registers[906][6] , \registers[906][5] , \registers[906][4] ,
         \registers[906][3] , \registers[906][2] , \registers[906][1] ,
         \registers[906][0] , \registers[905][7] , \registers[905][6] ,
         \registers[905][5] , \registers[905][4] , \registers[905][3] ,
         \registers[905][2] , \registers[905][1] , \registers[905][0] ,
         \registers[904][7] , \registers[904][6] , \registers[904][5] ,
         \registers[904][4] , \registers[904][3] , \registers[904][2] ,
         \registers[904][1] , \registers[904][0] , \registers[903][7] ,
         \registers[903][6] , \registers[903][5] , \registers[903][4] ,
         \registers[903][3] , \registers[903][2] , \registers[903][1] ,
         \registers[903][0] , \registers[902][7] , \registers[902][6] ,
         \registers[902][5] , \registers[902][4] , \registers[902][3] ,
         \registers[902][2] , \registers[902][1] , \registers[902][0] ,
         \registers[901][7] , \registers[901][6] , \registers[901][5] ,
         \registers[901][4] , \registers[901][3] , \registers[901][2] ,
         \registers[901][1] , \registers[901][0] , \registers[900][7] ,
         \registers[900][6] , \registers[900][5] , \registers[900][4] ,
         \registers[900][3] , \registers[900][2] , \registers[900][1] ,
         \registers[900][0] , \registers[899][7] , \registers[899][6] ,
         \registers[899][5] , \registers[899][4] , \registers[899][3] ,
         \registers[899][2] , \registers[899][1] , \registers[899][0] ,
         \registers[898][7] , \registers[898][6] , \registers[898][5] ,
         \registers[898][4] , \registers[898][3] , \registers[898][2] ,
         \registers[898][1] , \registers[898][0] , \registers[897][7] ,
         \registers[897][6] , \registers[897][5] , \registers[897][4] ,
         \registers[897][3] , \registers[897][2] , \registers[897][1] ,
         \registers[897][0] , \registers[896][7] , \registers[896][6] ,
         \registers[896][5] , \registers[896][4] , \registers[896][3] ,
         \registers[896][2] , \registers[896][1] , \registers[896][0] ,
         \registers[959][7] , \registers[959][6] , \registers[959][5] ,
         \registers[959][4] , \registers[959][3] , \registers[959][2] ,
         \registers[959][1] , \registers[959][0] , \registers[958][7] ,
         \registers[958][6] , \registers[958][5] , \registers[958][4] ,
         \registers[958][3] , \registers[958][2] , \registers[958][1] ,
         \registers[958][0] , \registers[957][7] , \registers[957][6] ,
         \registers[957][5] , \registers[957][4] , \registers[957][3] ,
         \registers[957][2] , \registers[957][1] , \registers[957][0] ,
         \registers[956][7] , \registers[956][6] , \registers[956][5] ,
         \registers[956][4] , \registers[956][3] , \registers[956][2] ,
         \registers[956][1] , \registers[956][0] , \registers[955][7] ,
         \registers[955][6] , \registers[955][5] , \registers[955][4] ,
         \registers[955][3] , \registers[955][2] , \registers[955][1] ,
         \registers[955][0] , \registers[954][7] , \registers[954][6] ,
         \registers[954][5] , \registers[954][4] , \registers[954][3] ,
         \registers[954][2] , \registers[954][1] , \registers[954][0] ,
         \registers[953][7] , \registers[953][6] , \registers[953][5] ,
         \registers[953][4] , \registers[953][3] , \registers[953][2] ,
         \registers[953][1] , \registers[953][0] , \registers[952][7] ,
         \registers[952][6] , \registers[952][5] , \registers[952][4] ,
         \registers[952][3] , \registers[952][2] , \registers[952][1] ,
         \registers[952][0] , \registers[951][7] , \registers[951][6] ,
         \registers[951][5] , \registers[951][4] , \registers[951][3] ,
         \registers[951][2] , \registers[951][1] , \registers[951][0] ,
         \registers[950][7] , \registers[950][6] , \registers[950][5] ,
         \registers[950][4] , \registers[950][3] , \registers[950][2] ,
         \registers[950][1] , \registers[950][0] , \registers[949][7] ,
         \registers[949][6] , \registers[949][5] , \registers[949][4] ,
         \registers[949][3] , \registers[949][2] , \registers[949][1] ,
         \registers[949][0] , \registers[948][7] , \registers[948][6] ,
         \registers[948][5] , \registers[948][4] , \registers[948][3] ,
         \registers[948][2] , \registers[948][1] , \registers[948][0] ,
         \registers[947][7] , \registers[947][6] , \registers[947][5] ,
         \registers[947][4] , \registers[947][3] , \registers[947][2] ,
         \registers[947][1] , \registers[947][0] , \registers[946][7] ,
         \registers[946][6] , \registers[946][5] , \registers[946][4] ,
         \registers[946][3] , \registers[946][2] , \registers[946][1] ,
         \registers[946][0] , \registers[945][7] , \registers[945][6] ,
         \registers[945][5] , \registers[945][4] , \registers[945][3] ,
         \registers[945][2] , \registers[945][1] , \registers[945][0] ,
         \registers[944][7] , \registers[944][6] , \registers[944][5] ,
         \registers[944][4] , \registers[944][3] , \registers[944][2] ,
         \registers[944][1] , \registers[944][0] , \registers[943][7] ,
         \registers[943][6] , \registers[943][5] , \registers[943][4] ,
         \registers[943][3] , \registers[943][2] , \registers[943][1] ,
         \registers[943][0] , \registers[942][7] , \registers[942][6] ,
         \registers[942][5] , \registers[942][4] , \registers[942][3] ,
         \registers[942][2] , \registers[942][1] , \registers[942][0] ,
         \registers[941][7] , \registers[941][6] , \registers[941][5] ,
         \registers[941][4] , \registers[941][3] , \registers[941][2] ,
         \registers[941][1] , \registers[941][0] , \registers[940][7] ,
         \registers[940][6] , \registers[940][5] , \registers[940][4] ,
         \registers[940][3] , \registers[940][2] , \registers[940][1] ,
         \registers[940][0] , \registers[939][7] , \registers[939][6] ,
         \registers[939][5] , \registers[939][4] , \registers[939][3] ,
         \registers[939][2] , \registers[939][1] , \registers[939][0] ,
         \registers[938][7] , \registers[938][6] , \registers[938][5] ,
         \registers[938][4] , \registers[938][3] , \registers[938][2] ,
         \registers[938][1] , \registers[938][0] , \registers[937][7] ,
         \registers[937][6] , \registers[937][5] , \registers[937][4] ,
         \registers[937][3] , \registers[937][2] , \registers[937][1] ,
         \registers[937][0] , \registers[936][7] , \registers[936][6] ,
         \registers[936][5] , \registers[936][4] , \registers[936][3] ,
         \registers[936][2] , \registers[936][1] , \registers[936][0] ,
         \registers[935][7] , \registers[935][6] , \registers[935][5] ,
         \registers[935][4] , \registers[935][3] , \registers[935][2] ,
         \registers[935][1] , \registers[935][0] , \registers[934][7] ,
         \registers[934][6] , \registers[934][5] , \registers[934][4] ,
         \registers[934][3] , \registers[934][2] , \registers[934][1] ,
         \registers[934][0] , \registers[933][7] , \registers[933][6] ,
         \registers[933][5] , \registers[933][4] , \registers[933][3] ,
         \registers[933][2] , \registers[933][1] , \registers[933][0] ,
         \registers[932][7] , \registers[932][6] , \registers[932][5] ,
         \registers[932][4] , \registers[932][3] , \registers[932][2] ,
         \registers[932][1] , \registers[932][0] , \registers[931][7] ,
         \registers[931][6] , \registers[931][5] , \registers[931][4] ,
         \registers[931][3] , \registers[931][2] , \registers[931][1] ,
         \registers[931][0] , \registers[930][7] , \registers[930][6] ,
         \registers[930][5] , \registers[930][4] , \registers[930][3] ,
         \registers[930][2] , \registers[930][1] , \registers[930][0] ,
         \registers[929][7] , \registers[929][6] , \registers[929][5] ,
         \registers[929][4] , \registers[929][3] , \registers[929][2] ,
         \registers[929][1] , \registers[929][0] , \registers[928][7] ,
         \registers[928][6] , \registers[928][5] , \registers[928][4] ,
         \registers[928][3] , \registers[928][2] , \registers[928][1] ,
         \registers[928][0] , \registers[991][7] , \registers[991][6] ,
         \registers[991][5] , \registers[991][4] , \registers[991][3] ,
         \registers[991][2] , \registers[991][1] , \registers[991][0] ,
         \registers[990][7] , \registers[990][6] , \registers[990][5] ,
         \registers[990][4] , \registers[990][3] , \registers[990][2] ,
         \registers[990][1] , \registers[990][0] , \registers[989][7] ,
         \registers[989][6] , \registers[989][5] , \registers[989][4] ,
         \registers[989][3] , \registers[989][2] , \registers[989][1] ,
         \registers[989][0] , \registers[988][7] , \registers[988][6] ,
         \registers[988][5] , \registers[988][4] , \registers[988][3] ,
         \registers[988][2] , \registers[988][1] , \registers[988][0] ,
         \registers[987][7] , \registers[987][6] , \registers[987][5] ,
         \registers[987][4] , \registers[987][3] , \registers[987][2] ,
         \registers[987][1] , \registers[987][0] , \registers[986][7] ,
         \registers[986][6] , \registers[986][5] , \registers[986][4] ,
         \registers[986][3] , \registers[986][2] , \registers[986][1] ,
         \registers[986][0] , \registers[985][7] , \registers[985][6] ,
         \registers[985][5] , \registers[985][4] , \registers[985][3] ,
         \registers[985][2] , \registers[985][1] , \registers[985][0] ,
         \registers[984][7] , \registers[984][6] , \registers[984][5] ,
         \registers[984][4] , \registers[984][3] , \registers[984][2] ,
         \registers[984][1] , \registers[984][0] , \registers[983][7] ,
         \registers[983][6] , \registers[983][5] , \registers[983][4] ,
         \registers[983][3] , \registers[983][2] , \registers[983][1] ,
         \registers[983][0] , \registers[982][7] , \registers[982][6] ,
         \registers[982][5] , \registers[982][4] , \registers[982][3] ,
         \registers[982][2] , \registers[982][1] , \registers[982][0] ,
         \registers[981][7] , \registers[981][6] , \registers[981][5] ,
         \registers[981][4] , \registers[981][3] , \registers[981][2] ,
         \registers[981][1] , \registers[981][0] , \registers[980][7] ,
         \registers[980][6] , \registers[980][5] , \registers[980][4] ,
         \registers[980][3] , \registers[980][2] , \registers[980][1] ,
         \registers[980][0] , \registers[979][7] , \registers[979][6] ,
         \registers[979][5] , \registers[979][4] , \registers[979][3] ,
         \registers[979][2] , \registers[979][1] , \registers[979][0] ,
         \registers[978][7] , \registers[978][6] , \registers[978][5] ,
         \registers[978][4] , \registers[978][3] , \registers[978][2] ,
         \registers[978][1] , \registers[978][0] , \registers[977][7] ,
         \registers[977][6] , \registers[977][5] , \registers[977][4] ,
         \registers[977][3] , \registers[977][2] , \registers[977][1] ,
         \registers[977][0] , \registers[976][7] , \registers[976][6] ,
         \registers[976][5] , \registers[976][4] , \registers[976][3] ,
         \registers[976][2] , \registers[976][1] , \registers[976][0] ,
         \registers[975][7] , \registers[975][6] , \registers[975][5] ,
         \registers[975][4] , \registers[975][3] , \registers[975][2] ,
         \registers[975][1] , \registers[975][0] , \registers[974][7] ,
         \registers[974][6] , \registers[974][5] , \registers[974][4] ,
         \registers[974][3] , \registers[974][2] , \registers[974][1] ,
         \registers[974][0] , \registers[973][7] , \registers[973][6] ,
         \registers[973][5] , \registers[973][4] , \registers[973][3] ,
         \registers[973][2] , \registers[973][1] , \registers[973][0] ,
         \registers[972][7] , \registers[972][6] , \registers[972][5] ,
         \registers[972][4] , \registers[972][3] , \registers[972][2] ,
         \registers[972][1] , \registers[972][0] , \registers[971][7] ,
         \registers[971][6] , \registers[971][5] , \registers[971][4] ,
         \registers[971][3] , \registers[971][2] , \registers[971][1] ,
         \registers[971][0] , \registers[970][7] , \registers[970][6] ,
         \registers[970][5] , \registers[970][4] , \registers[970][3] ,
         \registers[970][2] , \registers[970][1] , \registers[970][0] ,
         \registers[969][7] , \registers[969][6] , \registers[969][5] ,
         \registers[969][4] , \registers[969][3] , \registers[969][2] ,
         \registers[969][1] , \registers[969][0] , \registers[968][7] ,
         \registers[968][6] , \registers[968][5] , \registers[968][4] ,
         \registers[968][3] , \registers[968][2] , \registers[968][1] ,
         \registers[968][0] , \registers[967][7] , \registers[967][6] ,
         \registers[967][5] , \registers[967][4] , \registers[967][3] ,
         \registers[967][2] , \registers[967][1] , \registers[967][0] ,
         \registers[966][7] , \registers[966][6] , \registers[966][5] ,
         \registers[966][4] , \registers[966][3] , \registers[966][2] ,
         \registers[966][1] , \registers[966][0] , \registers[965][7] ,
         \registers[965][6] , \registers[965][5] , \registers[965][4] ,
         \registers[965][3] , \registers[965][2] , \registers[965][1] ,
         \registers[965][0] , \registers[964][7] , \registers[964][6] ,
         \registers[964][5] , \registers[964][4] , \registers[964][3] ,
         \registers[964][2] , \registers[964][1] , \registers[964][0] ,
         \registers[963][7] , \registers[963][6] , \registers[963][5] ,
         \registers[963][4] , \registers[963][3] , \registers[963][2] ,
         \registers[963][1] , \registers[963][0] , \registers[962][7] ,
         \registers[962][6] , \registers[962][5] , \registers[962][4] ,
         \registers[962][3] , \registers[962][2] , \registers[962][1] ,
         \registers[962][0] , \registers[961][7] , \registers[961][6] ,
         \registers[961][5] , \registers[961][4] , \registers[961][3] ,
         \registers[961][2] , \registers[961][1] , \registers[961][0] ,
         \registers[960][7] , \registers[960][6] , \registers[960][5] ,
         \registers[960][4] , \registers[960][3] , \registers[960][2] ,
         \registers[960][1] , \registers[960][0] , \registers[1023][7] ,
         \registers[1023][6] , \registers[1023][5] , \registers[1023][4] ,
         \registers[1023][3] , \registers[1023][2] , \registers[1023][1] ,
         \registers[1023][0] , \registers[1022][7] , \registers[1022][6] ,
         \registers[1022][5] , \registers[1022][4] , \registers[1022][3] ,
         \registers[1022][2] , \registers[1022][1] , \registers[1022][0] ,
         \registers[1021][7] , \registers[1021][6] , \registers[1021][5] ,
         \registers[1021][4] , \registers[1021][3] , \registers[1021][2] ,
         \registers[1021][1] , \registers[1021][0] , \registers[1020][7] ,
         \registers[1020][6] , \registers[1020][5] , \registers[1020][4] ,
         \registers[1020][3] , \registers[1020][2] , \registers[1020][1] ,
         \registers[1020][0] , \registers[1019][7] , \registers[1019][6] ,
         \registers[1019][5] , \registers[1019][4] , \registers[1019][3] ,
         \registers[1019][2] , \registers[1019][1] , \registers[1019][0] ,
         \registers[1018][7] , \registers[1018][6] , \registers[1018][5] ,
         \registers[1018][4] , \registers[1018][3] , \registers[1018][2] ,
         \registers[1018][1] , \registers[1018][0] , \registers[1017][7] ,
         \registers[1017][6] , \registers[1017][5] , \registers[1017][4] ,
         \registers[1017][3] , \registers[1017][2] , \registers[1017][1] ,
         \registers[1017][0] , \registers[1016][7] , \registers[1016][6] ,
         \registers[1016][5] , \registers[1016][4] , \registers[1016][3] ,
         \registers[1016][2] , \registers[1016][1] , \registers[1016][0] ,
         \registers[1015][7] , \registers[1015][6] , \registers[1015][5] ,
         \registers[1015][4] , \registers[1015][3] , \registers[1015][2] ,
         \registers[1015][1] , \registers[1015][0] , \registers[1014][7] ,
         \registers[1014][6] , \registers[1014][5] , \registers[1014][4] ,
         \registers[1014][3] , \registers[1014][2] , \registers[1014][1] ,
         \registers[1014][0] , \registers[1013][7] , \registers[1013][6] ,
         \registers[1013][5] , \registers[1013][4] , \registers[1013][3] ,
         \registers[1013][2] , \registers[1013][1] , \registers[1013][0] ,
         \registers[1012][7] , \registers[1012][6] , \registers[1012][5] ,
         \registers[1012][4] , \registers[1012][3] , \registers[1012][2] ,
         \registers[1012][1] , \registers[1012][0] , \registers[1011][7] ,
         \registers[1011][6] , \registers[1011][5] , \registers[1011][4] ,
         \registers[1011][3] , \registers[1011][2] , \registers[1011][1] ,
         \registers[1011][0] , \registers[1010][7] , \registers[1010][6] ,
         \registers[1010][5] , \registers[1010][4] , \registers[1010][3] ,
         \registers[1010][2] , \registers[1010][1] , \registers[1010][0] ,
         \registers[1009][7] , \registers[1009][6] , \registers[1009][5] ,
         \registers[1009][4] , \registers[1009][3] , \registers[1009][2] ,
         \registers[1009][1] , \registers[1009][0] , \registers[1008][7] ,
         \registers[1008][6] , \registers[1008][5] , \registers[1008][4] ,
         \registers[1008][3] , \registers[1008][2] , \registers[1008][1] ,
         \registers[1008][0] , \registers[1007][7] , \registers[1007][6] ,
         \registers[1007][5] , \registers[1007][4] , \registers[1007][3] ,
         \registers[1007][2] , \registers[1007][1] , \registers[1007][0] ,
         \registers[1006][7] , \registers[1006][6] , \registers[1006][5] ,
         \registers[1006][4] , \registers[1006][3] , \registers[1006][2] ,
         \registers[1006][1] , \registers[1006][0] , \registers[1005][7] ,
         \registers[1005][6] , \registers[1005][5] , \registers[1005][4] ,
         \registers[1005][3] , \registers[1005][2] , \registers[1005][1] ,
         \registers[1005][0] , \registers[1004][7] , \registers[1004][6] ,
         \registers[1004][5] , \registers[1004][4] , \registers[1004][3] ,
         \registers[1004][2] , \registers[1004][1] , \registers[1004][0] ,
         \registers[1003][7] , \registers[1003][6] , \registers[1003][5] ,
         \registers[1003][4] , \registers[1003][3] , \registers[1003][2] ,
         \registers[1003][1] , \registers[1003][0] , \registers[1002][7] ,
         \registers[1002][6] , \registers[1002][5] , \registers[1002][4] ,
         \registers[1002][3] , \registers[1002][2] , \registers[1002][1] ,
         \registers[1002][0] , \registers[1001][7] , \registers[1001][6] ,
         \registers[1001][5] , \registers[1001][4] , \registers[1001][3] ,
         \registers[1001][2] , \registers[1001][1] , \registers[1001][0] ,
         \registers[1000][7] , \registers[1000][6] , \registers[1000][5] ,
         \registers[1000][4] , \registers[1000][3] , \registers[1000][2] ,
         \registers[1000][1] , \registers[1000][0] , \registers[999][7] ,
         \registers[999][6] , \registers[999][5] , \registers[999][4] ,
         \registers[999][3] , \registers[999][2] , \registers[999][1] ,
         \registers[999][0] , \registers[998][7] , \registers[998][6] ,
         \registers[998][5] , \registers[998][4] , \registers[998][3] ,
         \registers[998][2] , \registers[998][1] , \registers[998][0] ,
         \registers[997][7] , \registers[997][6] , \registers[997][5] ,
         \registers[997][4] , \registers[997][3] , \registers[997][2] ,
         \registers[997][1] , \registers[997][0] , \registers[996][7] ,
         \registers[996][6] , \registers[996][5] , \registers[996][4] ,
         \registers[996][3] , \registers[996][2] , \registers[996][1] ,
         \registers[996][0] , \registers[995][7] , \registers[995][6] ,
         \registers[995][5] , \registers[995][4] , \registers[995][3] ,
         \registers[995][2] , \registers[995][1] , \registers[995][0] ,
         \registers[994][7] , \registers[994][6] , \registers[994][5] ,
         \registers[994][4] , \registers[994][3] , \registers[994][2] ,
         \registers[994][1] , \registers[994][0] , \registers[993][7] ,
         \registers[993][6] , \registers[993][5] , \registers[993][4] ,
         \registers[993][3] , \registers[993][2] , \registers[993][1] ,
         \registers[993][0] , \registers[992][7] , \registers[992][6] ,
         \registers[992][5] , \registers[992][4] , \registers[992][3] ,
         \registers[992][2] , \registers[992][1] , \registers[992][0] , N108,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, StartBit, N1195, N1197, N1198, N1199, N1200,
         N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210,
         N1211, N1212, N1213, N1214, N1215, N1216, N1227, N1228, N1229, N1230,
         N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240,
         N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1308, N1309, N1310,
         N1311, N1312, N1313, N1314, N1315, N1349, N1350, N1351, N1352, N1353,
         N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363,
         N1364, N1365, N1366, N1367, N1387, N1388, N1389, N1390, N1391, N1392,
         N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402,
         N1403, N1404, N1405, N1406, N1407, N1408, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1196, n1197,
         n1199, n1200, n1203, n1206, n1208, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1271, n1272, n1274, n1276, n1278, n1280,
         n1282, n1284, n1286, n1288, n1290, n1292, n1294, n1296, n1298, n1300,
         n1302, n1304, n1306, n1308, n1310, n1312, n1314, n1316, n1318, n1320,
         n1322, n1324, n1326, n1328, n1330, n1332, n1334, n1366, n1367, n1369,
         n1401, n1403, n1435, n1437, n1469, n1471, n1503, n1505, n1537, n1539,
         n1571, n1573, n1605, n1606, n1608, n1641, n1674, n1707, n1740, n1773,
         n1806, n1839, n1871, n1873, n1906, n1939, n1972, n2005, n2038, n2071,
         n2104, n2136, n2138, n2171, n2204, n2237, n2270, n2303, n2336, n2337,
         n2338, n2340, n2342, n2344, n2346, n2348, n2350, n2352, n2354, n2363,
         n2372, n2381, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, N1287, N1286, N1285, N1284,
         N1283, N1282, N1281, N1280, N1279, N1278, \r402/carry[9] ,
         \r402/carry[8] , \r402/carry[7] , \r402/carry[6] , \r402/carry[5] ,
         \r402/carry[4] , \r402/carry[3] , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1195, n1198, n1201, n1202, n1204, n1205, n1207, n1209,
         n1210, n1270, n1273, n1275, n1277, n1279, n1281, n1283, n1285, n1287,
         n1289, n1291, n1293, n1295, n1297, n1299, n1301, n1303, n1305, n1307,
         n1309, n1311, n1313, n1315, n1317, n1319, n1321, n1323, n1325, n1327,
         n1329, n1331, n1333, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1368, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1402, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1436, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1470, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1504, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1538, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1572, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1607, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1872, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2137, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2339, n2341, n2343, n2345, n2347, n2349, n2351,
         n2353, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2382, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973;
  wire   [19:0] M2;
  wire   [19:0] N2;
  wire   [1:0] state;
  wire   [12:0] pixel_i;
  wire   [18:0] block_i;
  wire   [3:0] param_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35;

  Control_And_Registers_DW_cmp_0 gt_124 ( .A({N1387, N1367, N1366, N1365, 
        N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, 
        N1354, N1353, N1352, N1351, N1350, N1349}), .B({N1407, N1406, N1405, 
        N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, 
        N1394, N1393, N1392, N1391, N1390, N1389, N1388}), .TC(1'b0), .GE_LT(
        1'b0), .GE_GT_EQ(1'b1), .GE_LT_GT_LE(N1408) );
  Control_And_Registers_DW01_add_15 add_0_root_add_99_3 ( .A({N1216, N1215, 
        N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207}), .B({N1206, 
        N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197}), .CI(
        1'b0), .SUM({N77, N76, N75, N74, N73, N72, N71, N70, N69, N68}) );
  Control_And_Registers_DW01_inc_0 r409 ( .A({1'b0, block_i}), .SUM({N1387, 
        N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, 
        N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349}) );
  Control_And_Registers_DW01_inc_1 r405 ( .A({pixel_i[12:6], n9, pixel_i[4:1], 
        N1197}), .SUM({N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, 
        N1239, N1238, N1237, N1236, N1235}) );
  Control_And_Registers_DW_mult_uns_2 mult_58 ( .a({data_in[15:8], n8377, 
        n8319, n8261, n8203, n8161, n8107, n8051, n8666}), .b({data_in[15:8], 
        n8377, n8319, n8261, n8203, n8161, n8105, n8049, n7994}), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, N147, N146, N145, 
        N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, 
        N132, N131, N130, SYNOPSYS_UNCONNECTED__12, N128}) );
  Control_And_Registers_DW_mult_uns_1 mult_56 ( .a({data_in[15:8], n8377, 
        n8319, n8261, n8203, n8161, n8106, n8050, n7994}), .b({data_in[15:8], 
        n8868, n8839, n8810, n8781, n8768, n8151, n8095, n8666}), .product({
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, N127, N126, N125, 
        N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, 
        N112, N111, N110, SYNOPSYS_UNCONNECTED__25, N108}) );
  Control_And_Registers_DW01_add_18 add_1_root_add_0_root_add_110_4 ( .A(
        N2[9:0]), .B({N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, 
        N1198, N1197}), .CI(1'b0), .SUM({N1287, N1286, N1285, N1284, N1283, 
        N1282, N1281, N1280, N1279, N1278}) );
  Control_And_Registers_DW01_add_17 add_0_root_add_0_root_add_110_4 ( .A({
        N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278}), 
        .B({N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, 
        N1207}), .CI(1'b0), .SUM({N87, N86, N85, N84, N83, N82, N81, N80, N79, 
        N78}) );
  Control_And_Registers_DW_mult_uns_0 r403 ( .a(block_i[9:0]), .b(M2[9:0]), 
        .product({SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, N1216, N1215, 
        N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207}) );
  Control_And_Registers_DW_div_uns_5 div_124 ( .a(N2), .b(M2), .quotient({
        N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, 
        N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388})
         );
  DFFHQX1 Image_Done_reg ( .D(n2425), .CK(clk), .Q(Image_Done) );
  EDFFX1 \param_i_reg[3]  ( .D(1'b0), .E(n1239), .CK(clk), .Q(param_i[3]) );
  EDFFX1 \registers_reg[1021][7]  ( .D(n8396), .E(n931), .CK(clk), .Q(
        \registers[1021][7] ) );
  EDFFX1 \registers_reg[1021][6]  ( .D(n8338), .E(n931), .CK(clk), .Q(
        \registers[1021][6] ) );
  EDFFX1 \registers_reg[1021][5]  ( .D(n8280), .E(n931), .CK(clk), .Q(
        \registers[1021][5] ) );
  EDFFX1 \registers_reg[1021][4]  ( .D(n8222), .E(n931), .CK(clk), .Q(
        \registers[1021][4] ) );
  EDFFX1 \registers_reg[1021][3]  ( .D(n8177), .E(n931), .CK(clk), .Q(
        \registers[1021][3] ) );
  EDFFX1 \registers_reg[1021][2]  ( .D(n8126), .E(n931), .CK(clk), .Q(
        \registers[1021][2] ) );
  EDFFX1 \registers_reg[1021][1]  ( .D(n8070), .E(n931), .CK(clk), .Q(
        \registers[1021][1] ) );
  EDFFX1 \registers_reg[1021][0]  ( .D(n8012), .E(n931), .CK(clk), .Q(
        \registers[1021][0] ) );
  EDFFX1 \registers_reg[1017][7]  ( .D(n8397), .E(n927), .CK(clk), .Q(
        \registers[1017][7] ) );
  EDFFX1 \registers_reg[1017][6]  ( .D(n8339), .E(n927), .CK(clk), .Q(
        \registers[1017][6] ) );
  EDFFX1 \registers_reg[1017][5]  ( .D(n8281), .E(n927), .CK(clk), .Q(
        \registers[1017][5] ) );
  EDFFX1 \registers_reg[1017][4]  ( .D(n8223), .E(n927), .CK(clk), .Q(
        \registers[1017][4] ) );
  EDFFX1 \registers_reg[1017][3]  ( .D(n8178), .E(n927), .CK(clk), .Q(
        \registers[1017][3] ) );
  EDFFX1 \registers_reg[1017][2]  ( .D(n8127), .E(n927), .CK(clk), .Q(
        \registers[1017][2] ) );
  EDFFX1 \registers_reg[1017][1]  ( .D(n8071), .E(n927), .CK(clk), .Q(
        \registers[1017][1] ) );
  EDFFX1 \registers_reg[1017][0]  ( .D(n8010), .E(n927), .CK(clk), .Q(
        \registers[1017][0] ) );
  EDFFX1 \registers_reg[1013][7]  ( .D(n8395), .E(n923), .CK(clk), .Q(
        \registers[1013][7] ) );
  EDFFX1 \registers_reg[1013][6]  ( .D(n8337), .E(n923), .CK(clk), .Q(
        \registers[1013][6] ) );
  EDFFX1 \registers_reg[1013][5]  ( .D(n8279), .E(n923), .CK(clk), .Q(
        \registers[1013][5] ) );
  EDFFX1 \registers_reg[1013][4]  ( .D(n8221), .E(n923), .CK(clk), .Q(
        \registers[1013][4] ) );
  EDFFX1 \registers_reg[1013][3]  ( .D(n8176), .E(n923), .CK(clk), .Q(
        \registers[1013][3] ) );
  EDFFX1 \registers_reg[1013][2]  ( .D(n8128), .E(n923), .CK(clk), .Q(
        \registers[1013][2] ) );
  EDFFX1 \registers_reg[1013][1]  ( .D(n8072), .E(n923), .CK(clk), .Q(
        \registers[1013][1] ) );
  EDFFX1 \registers_reg[1013][0]  ( .D(n8011), .E(n923), .CK(clk), .Q(
        \registers[1013][0] ) );
  EDFFX1 \registers_reg[1009][7]  ( .D(n8396), .E(n236), .CK(clk), .Q(
        \registers[1009][7] ) );
  EDFFX1 \registers_reg[1009][6]  ( .D(n8338), .E(n236), .CK(clk), .Q(
        \registers[1009][6] ) );
  EDFFX1 \registers_reg[1009][5]  ( .D(n8280), .E(n236), .CK(clk), .Q(
        \registers[1009][5] ) );
  EDFFX1 \registers_reg[1009][4]  ( .D(n8222), .E(n236), .CK(clk), .Q(
        \registers[1009][4] ) );
  EDFFX1 \registers_reg[1009][3]  ( .D(n8177), .E(n236), .CK(clk), .Q(
        \registers[1009][3] ) );
  EDFFX1 \registers_reg[1009][2]  ( .D(n8126), .E(n236), .CK(clk), .Q(
        \registers[1009][2] ) );
  EDFFX1 \registers_reg[1009][1]  ( .D(n8070), .E(n236), .CK(clk), .Q(
        \registers[1009][1] ) );
  EDFFX1 \registers_reg[1009][0]  ( .D(n8012), .E(n236), .CK(clk), .Q(
        \registers[1009][0] ) );
  EDFFX1 \registers_reg[1005][7]  ( .D(n8397), .E(n232), .CK(clk), .Q(
        \registers[1005][7] ) );
  EDFFX1 \registers_reg[1005][6]  ( .D(n8339), .E(n232), .CK(clk), .Q(
        \registers[1005][6] ) );
  EDFFX1 \registers_reg[1005][5]  ( .D(n8281), .E(n232), .CK(clk), .Q(
        \registers[1005][5] ) );
  EDFFX1 \registers_reg[1005][4]  ( .D(n8223), .E(n232), .CK(clk), .Q(
        \registers[1005][4] ) );
  EDFFX1 \registers_reg[1005][3]  ( .D(n8178), .E(n232), .CK(clk), .Q(
        \registers[1005][3] ) );
  EDFFX1 \registers_reg[1005][2]  ( .D(n8127), .E(n232), .CK(clk), .Q(
        \registers[1005][2] ) );
  EDFFX1 \registers_reg[1005][1]  ( .D(n8071), .E(n232), .CK(clk), .Q(
        \registers[1005][1] ) );
  EDFFX1 \registers_reg[1005][0]  ( .D(n8010), .E(n232), .CK(clk), .Q(
        \registers[1005][0] ) );
  EDFFX1 \registers_reg[1001][7]  ( .D(n8395), .E(n228), .CK(clk), .Q(
        \registers[1001][7] ) );
  EDFFX1 \registers_reg[1001][6]  ( .D(n8337), .E(n228), .CK(clk), .Q(
        \registers[1001][6] ) );
  EDFFX1 \registers_reg[1001][5]  ( .D(n8279), .E(n228), .CK(clk), .Q(
        \registers[1001][5] ) );
  EDFFX1 \registers_reg[1001][4]  ( .D(n8221), .E(n228), .CK(clk), .Q(
        \registers[1001][4] ) );
  EDFFX1 \registers_reg[1001][3]  ( .D(n8173), .E(n228), .CK(clk), .Q(
        \registers[1001][3] ) );
  EDFFX1 \registers_reg[1001][2]  ( .D(n8128), .E(n228), .CK(clk), .Q(
        \registers[1001][2] ) );
  EDFFX1 \registers_reg[1001][1]  ( .D(n8072), .E(n228), .CK(clk), .Q(
        \registers[1001][1] ) );
  EDFFX1 \registers_reg[1001][0]  ( .D(n8011), .E(n228), .CK(clk), .Q(
        \registers[1001][0] ) );
  EDFFX1 \registers_reg[997][7]  ( .D(n8396), .E(n384), .CK(clk), .Q(
        \registers[997][7] ) );
  EDFFX1 \registers_reg[997][6]  ( .D(n8338), .E(n384), .CK(clk), .Q(
        \registers[997][6] ) );
  EDFFX1 \registers_reg[997][5]  ( .D(n8280), .E(n384), .CK(clk), .Q(
        \registers[997][5] ) );
  EDFFX1 \registers_reg[997][4]  ( .D(n8222), .E(n384), .CK(clk), .Q(
        \registers[997][4] ) );
  EDFFX1 \registers_reg[997][3]  ( .D(n8174), .E(n384), .CK(clk), .Q(
        \registers[997][3] ) );
  EDFFX1 \registers_reg[997][2]  ( .D(n8126), .E(n384), .CK(clk), .Q(
        \registers[997][2] ) );
  EDFFX1 \registers_reg[997][1]  ( .D(n8070), .E(n384), .CK(clk), .Q(
        \registers[997][1] ) );
  EDFFX1 \registers_reg[997][0]  ( .D(n8012), .E(n384), .CK(clk), .Q(
        \registers[997][0] ) );
  EDFFX1 \registers_reg[993][7]  ( .D(n8397), .E(n380), .CK(clk), .Q(
        \registers[993][7] ) );
  EDFFX1 \registers_reg[993][6]  ( .D(n8339), .E(n380), .CK(clk), .Q(
        \registers[993][6] ) );
  EDFFX1 \registers_reg[993][5]  ( .D(n8281), .E(n380), .CK(clk), .Q(
        \registers[993][5] ) );
  EDFFX1 \registers_reg[993][4]  ( .D(n8223), .E(n380), .CK(clk), .Q(
        \registers[993][4] ) );
  EDFFX1 \registers_reg[993][3]  ( .D(n8175), .E(n380), .CK(clk), .Q(
        \registers[993][3] ) );
  EDFFX1 \registers_reg[993][2]  ( .D(n8127), .E(n380), .CK(clk), .Q(
        \registers[993][2] ) );
  EDFFX1 \registers_reg[993][1]  ( .D(n8071), .E(n380), .CK(clk), .Q(
        \registers[993][1] ) );
  EDFFX1 \registers_reg[993][0]  ( .D(n8010), .E(n380), .CK(clk), .Q(
        \registers[993][0] ) );
  EDFFX1 \registers_reg[989][7]  ( .D(n8395), .E(n919), .CK(clk), .Q(
        \registers[989][7] ) );
  EDFFX1 \registers_reg[989][6]  ( .D(n8337), .E(n919), .CK(clk), .Q(
        \registers[989][6] ) );
  EDFFX1 \registers_reg[989][5]  ( .D(n8279), .E(n919), .CK(clk), .Q(
        \registers[989][5] ) );
  EDFFX1 \registers_reg[989][4]  ( .D(n8221), .E(n919), .CK(clk), .Q(
        \registers[989][4] ) );
  EDFFX1 \registers_reg[989][3]  ( .D(n8173), .E(n919), .CK(clk), .Q(
        \registers[989][3] ) );
  EDFFX1 \registers_reg[989][2]  ( .D(n8128), .E(n919), .CK(clk), .Q(
        \registers[989][2] ) );
  EDFFX1 \registers_reg[989][1]  ( .D(n8072), .E(n919), .CK(clk), .Q(
        \registers[989][1] ) );
  EDFFX1 \registers_reg[989][0]  ( .D(n8011), .E(n919), .CK(clk), .Q(
        \registers[989][0] ) );
  EDFFX1 \registers_reg[985][7]  ( .D(n8396), .E(n915), .CK(clk), .Q(
        \registers[985][7] ) );
  EDFFX1 \registers_reg[985][6]  ( .D(n8338), .E(n915), .CK(clk), .Q(
        \registers[985][6] ) );
  EDFFX1 \registers_reg[985][5]  ( .D(n8280), .E(n915), .CK(clk), .Q(
        \registers[985][5] ) );
  EDFFX1 \registers_reg[985][4]  ( .D(n8222), .E(n915), .CK(clk), .Q(
        \registers[985][4] ) );
  EDFFX1 \registers_reg[985][3]  ( .D(n8174), .E(n915), .CK(clk), .Q(
        \registers[985][3] ) );
  EDFFX1 \registers_reg[985][2]  ( .D(n8123), .E(n915), .CK(clk), .Q(
        \registers[985][2] ) );
  EDFFX1 \registers_reg[985][1]  ( .D(n8067), .E(n915), .CK(clk), .Q(
        \registers[985][1] ) );
  EDFFX1 \registers_reg[985][0]  ( .D(n8012), .E(n915), .CK(clk), .Q(
        \registers[985][0] ) );
  EDFFX1 \registers_reg[981][7]  ( .D(n8397), .E(n911), .CK(clk), .Q(
        \registers[981][7] ) );
  EDFFX1 \registers_reg[981][6]  ( .D(n8339), .E(n911), .CK(clk), .Q(
        \registers[981][6] ) );
  EDFFX1 \registers_reg[981][5]  ( .D(n8281), .E(n911), .CK(clk), .Q(
        \registers[981][5] ) );
  EDFFX1 \registers_reg[981][4]  ( .D(n8223), .E(n911), .CK(clk), .Q(
        \registers[981][4] ) );
  EDFFX1 \registers_reg[981][3]  ( .D(n8175), .E(n911), .CK(clk), .Q(
        \registers[981][3] ) );
  EDFFX1 \registers_reg[981][2]  ( .D(n8124), .E(n911), .CK(clk), .Q(
        \registers[981][2] ) );
  EDFFX1 \registers_reg[981][1]  ( .D(n8068), .E(n911), .CK(clk), .Q(
        \registers[981][1] ) );
  EDFFX1 \registers_reg[981][0]  ( .D(n8007), .E(n911), .CK(clk), .Q(
        \registers[981][0] ) );
  EDFFX1 \registers_reg[977][7]  ( .D(n8393), .E(n224), .CK(clk), .Q(
        \registers[977][7] ) );
  EDFFX1 \registers_reg[977][6]  ( .D(n8335), .E(n224), .CK(clk), .Q(
        \registers[977][6] ) );
  EDFFX1 \registers_reg[977][5]  ( .D(n8277), .E(n224), .CK(clk), .Q(
        \registers[977][5] ) );
  EDFFX1 \registers_reg[977][4]  ( .D(n8219), .E(n224), .CK(clk), .Q(
        \registers[977][4] ) );
  EDFFX1 \registers_reg[977][3]  ( .D(n8173), .E(n224), .CK(clk), .Q(
        \registers[977][3] ) );
  EDFFX1 \registers_reg[977][2]  ( .D(n8125), .E(n224), .CK(clk), .Q(
        \registers[977][2] ) );
  EDFFX1 \registers_reg[977][1]  ( .D(n8069), .E(n224), .CK(clk), .Q(
        \registers[977][1] ) );
  EDFFX1 \registers_reg[977][0]  ( .D(n8008), .E(n224), .CK(clk), .Q(
        \registers[977][0] ) );
  EDFFX1 \registers_reg[973][7]  ( .D(n8394), .E(n220), .CK(clk), .Q(
        \registers[973][7] ) );
  EDFFX1 \registers_reg[973][6]  ( .D(n8336), .E(n220), .CK(clk), .Q(
        \registers[973][6] ) );
  EDFFX1 \registers_reg[973][5]  ( .D(n8278), .E(n220), .CK(clk), .Q(
        \registers[973][5] ) );
  EDFFX1 \registers_reg[973][4]  ( .D(n8220), .E(n220), .CK(clk), .Q(
        \registers[973][4] ) );
  EDFFX1 \registers_reg[973][3]  ( .D(n8174), .E(n220), .CK(clk), .Q(
        \registers[973][3] ) );
  EDFFX1 \registers_reg[973][2]  ( .D(n8123), .E(n220), .CK(clk), .Q(
        \registers[973][2] ) );
  EDFFX1 \registers_reg[973][1]  ( .D(n8067), .E(n220), .CK(clk), .Q(
        \registers[973][1] ) );
  EDFFX1 \registers_reg[973][0]  ( .D(n8009), .E(n220), .CK(clk), .Q(
        \registers[973][0] ) );
  EDFFX1 \registers_reg[969][7]  ( .D(n8392), .E(n216), .CK(clk), .Q(
        \registers[969][7] ) );
  EDFFX1 \registers_reg[969][6]  ( .D(n8334), .E(n216), .CK(clk), .Q(
        \registers[969][6] ) );
  EDFFX1 \registers_reg[969][5]  ( .D(n8276), .E(n216), .CK(clk), .Q(
        \registers[969][5] ) );
  EDFFX1 \registers_reg[969][4]  ( .D(n8218), .E(n216), .CK(clk), .Q(
        \registers[969][4] ) );
  EDFFX1 \registers_reg[969][3]  ( .D(n8175), .E(n216), .CK(clk), .Q(
        \registers[969][3] ) );
  EDFFX1 \registers_reg[969][2]  ( .D(n8124), .E(n216), .CK(clk), .Q(
        \registers[969][2] ) );
  EDFFX1 \registers_reg[969][1]  ( .D(n8068), .E(n216), .CK(clk), .Q(
        \registers[969][1] ) );
  EDFFX1 \registers_reg[969][0]  ( .D(n8007), .E(n216), .CK(clk), .Q(
        \registers[969][0] ) );
  EDFFX1 \registers_reg[965][7]  ( .D(n8393), .E(n377), .CK(clk), .Q(
        \registers[965][7] ) );
  EDFFX1 \registers_reg[965][6]  ( .D(n8335), .E(n377), .CK(clk), .Q(
        \registers[965][6] ) );
  EDFFX1 \registers_reg[965][5]  ( .D(n8277), .E(n377), .CK(clk), .Q(
        \registers[965][5] ) );
  EDFFX1 \registers_reg[965][4]  ( .D(n8219), .E(n377), .CK(clk), .Q(
        \registers[965][4] ) );
  EDFFX1 \registers_reg[965][3]  ( .D(n8173), .E(n377), .CK(clk), .Q(
        \registers[965][3] ) );
  EDFFX1 \registers_reg[965][2]  ( .D(n8125), .E(n377), .CK(clk), .Q(
        \registers[965][2] ) );
  EDFFX1 \registers_reg[965][1]  ( .D(n8069), .E(n377), .CK(clk), .Q(
        \registers[965][1] ) );
  EDFFX1 \registers_reg[965][0]  ( .D(n8008), .E(n377), .CK(clk), .Q(
        \registers[965][0] ) );
  EDFFX1 \registers_reg[961][7]  ( .D(n8394), .E(n373), .CK(clk), .Q(
        \registers[961][7] ) );
  EDFFX1 \registers_reg[961][6]  ( .D(n8336), .E(n373), .CK(clk), .Q(
        \registers[961][6] ) );
  EDFFX1 \registers_reg[961][5]  ( .D(n8278), .E(n373), .CK(clk), .Q(
        \registers[961][5] ) );
  EDFFX1 \registers_reg[961][4]  ( .D(n8220), .E(n373), .CK(clk), .Q(
        \registers[961][4] ) );
  EDFFX1 \registers_reg[961][3]  ( .D(n8174), .E(n373), .CK(clk), .Q(
        \registers[961][3] ) );
  EDFFX1 \registers_reg[961][2]  ( .D(n8123), .E(n373), .CK(clk), .Q(
        \registers[961][2] ) );
  EDFFX1 \registers_reg[961][1]  ( .D(n8067), .E(n373), .CK(clk), .Q(
        \registers[961][1] ) );
  EDFFX1 \registers_reg[961][0]  ( .D(n8009), .E(n373), .CK(clk), .Q(
        \registers[961][0] ) );
  EDFFX1 \registers_reg[957][7]  ( .D(n8393), .E(n907), .CK(clk), .Q(
        \registers[957][7] ) );
  EDFFX1 \registers_reg[957][6]  ( .D(n8335), .E(n907), .CK(clk), .Q(
        \registers[957][6] ) );
  EDFFX1 \registers_reg[957][5]  ( .D(n8277), .E(n907), .CK(clk), .Q(
        \registers[957][5] ) );
  EDFFX1 \registers_reg[957][4]  ( .D(n8219), .E(n907), .CK(clk), .Q(
        \registers[957][4] ) );
  EDFFX1 \registers_reg[957][3]  ( .D(n8173), .E(n907), .CK(clk), .Q(
        \registers[957][3] ) );
  EDFFX1 \registers_reg[957][2]  ( .D(n8125), .E(n907), .CK(clk), .Q(
        \registers[957][2] ) );
  EDFFX1 \registers_reg[957][1]  ( .D(n8069), .E(n907), .CK(clk), .Q(
        \registers[957][1] ) );
  EDFFX1 \registers_reg[957][0]  ( .D(n8008), .E(n907), .CK(clk), .Q(
        \registers[957][0] ) );
  EDFFX1 \registers_reg[953][7]  ( .D(n8394), .E(n903), .CK(clk), .Q(
        \registers[953][7] ) );
  EDFFX1 \registers_reg[953][6]  ( .D(n8336), .E(n903), .CK(clk), .Q(
        \registers[953][6] ) );
  EDFFX1 \registers_reg[953][5]  ( .D(n8278), .E(n903), .CK(clk), .Q(
        \registers[953][5] ) );
  EDFFX1 \registers_reg[953][4]  ( .D(n8220), .E(n903), .CK(clk), .Q(
        \registers[953][4] ) );
  EDFFX1 \registers_reg[953][3]  ( .D(n8174), .E(n903), .CK(clk), .Q(
        \registers[953][3] ) );
  EDFFX1 \registers_reg[953][2]  ( .D(n8123), .E(n903), .CK(clk), .Q(
        \registers[953][2] ) );
  EDFFX1 \registers_reg[953][1]  ( .D(n8067), .E(n903), .CK(clk), .Q(
        \registers[953][1] ) );
  EDFFX1 \registers_reg[953][0]  ( .D(n8009), .E(n903), .CK(clk), .Q(
        \registers[953][0] ) );
  EDFFX1 \registers_reg[949][7]  ( .D(n8392), .E(n899), .CK(clk), .Q(
        \registers[949][7] ) );
  EDFFX1 \registers_reg[949][6]  ( .D(n8334), .E(n899), .CK(clk), .Q(
        \registers[949][6] ) );
  EDFFX1 \registers_reg[949][5]  ( .D(n8276), .E(n899), .CK(clk), .Q(
        \registers[949][5] ) );
  EDFFX1 \registers_reg[949][4]  ( .D(n8218), .E(n899), .CK(clk), .Q(
        \registers[949][4] ) );
  EDFFX1 \registers_reg[949][3]  ( .D(n8175), .E(n899), .CK(clk), .Q(
        \registers[949][3] ) );
  EDFFX1 \registers_reg[949][2]  ( .D(n8124), .E(n899), .CK(clk), .Q(
        \registers[949][2] ) );
  EDFFX1 \registers_reg[949][1]  ( .D(n8068), .E(n899), .CK(clk), .Q(
        \registers[949][1] ) );
  EDFFX1 \registers_reg[949][0]  ( .D(n8007), .E(n899), .CK(clk), .Q(
        \registers[949][0] ) );
  EDFFX1 \registers_reg[945][7]  ( .D(n8393), .E(n212), .CK(clk), .Q(
        \registers[945][7] ) );
  EDFFX1 \registers_reg[945][6]  ( .D(n8335), .E(n212), .CK(clk), .Q(
        \registers[945][6] ) );
  EDFFX1 \registers_reg[945][5]  ( .D(n8277), .E(n212), .CK(clk), .Q(
        \registers[945][5] ) );
  EDFFX1 \registers_reg[945][4]  ( .D(n8219), .E(n212), .CK(clk), .Q(
        \registers[945][4] ) );
  EDFFX1 \registers_reg[945][3]  ( .D(n8173), .E(n212), .CK(clk), .Q(
        \registers[945][3] ) );
  EDFFX1 \registers_reg[945][2]  ( .D(n8125), .E(n212), .CK(clk), .Q(
        \registers[945][2] ) );
  EDFFX1 \registers_reg[945][1]  ( .D(n8069), .E(n212), .CK(clk), .Q(
        \registers[945][1] ) );
  EDFFX1 \registers_reg[945][0]  ( .D(n8008), .E(n212), .CK(clk), .Q(
        \registers[945][0] ) );
  EDFFX1 \registers_reg[941][7]  ( .D(n8394), .E(n208), .CK(clk), .Q(
        \registers[941][7] ) );
  EDFFX1 \registers_reg[941][6]  ( .D(n8336), .E(n208), .CK(clk), .Q(
        \registers[941][6] ) );
  EDFFX1 \registers_reg[941][5]  ( .D(n8278), .E(n208), .CK(clk), .Q(
        \registers[941][5] ) );
  EDFFX1 \registers_reg[941][4]  ( .D(n8220), .E(n208), .CK(clk), .Q(
        \registers[941][4] ) );
  EDFFX1 \registers_reg[941][3]  ( .D(n8171), .E(n208), .CK(clk), .Q(
        \registers[941][3] ) );
  EDFFX1 \registers_reg[941][2]  ( .D(n8123), .E(n208), .CK(clk), .Q(
        \registers[941][2] ) );
  EDFFX1 \registers_reg[941][1]  ( .D(n8067), .E(n208), .CK(clk), .Q(
        \registers[941][1] ) );
  EDFFX1 \registers_reg[941][0]  ( .D(n8009), .E(n208), .CK(clk), .Q(
        \registers[941][0] ) );
  EDFFX1 \registers_reg[937][7]  ( .D(n8392), .E(n204), .CK(clk), .Q(
        \registers[937][7] ) );
  EDFFX1 \registers_reg[937][6]  ( .D(n8334), .E(n204), .CK(clk), .Q(
        \registers[937][6] ) );
  EDFFX1 \registers_reg[937][5]  ( .D(n8276), .E(n204), .CK(clk), .Q(
        \registers[937][5] ) );
  EDFFX1 \registers_reg[937][4]  ( .D(n8218), .E(n204), .CK(clk), .Q(
        \registers[937][4] ) );
  EDFFX1 \registers_reg[937][3]  ( .D(n8172), .E(n204), .CK(clk), .Q(
        \registers[937][3] ) );
  EDFFX1 \registers_reg[937][2]  ( .D(n8124), .E(n204), .CK(clk), .Q(
        \registers[937][2] ) );
  EDFFX1 \registers_reg[937][1]  ( .D(n8068), .E(n204), .CK(clk), .Q(
        \registers[937][1] ) );
  EDFFX1 \registers_reg[937][0]  ( .D(n8007), .E(n204), .CK(clk), .Q(
        \registers[937][0] ) );
  EDFFX1 \registers_reg[933][7]  ( .D(n8393), .E(n370), .CK(clk), .Q(
        \registers[933][7] ) );
  EDFFX1 \registers_reg[933][6]  ( .D(n8335), .E(n370), .CK(clk), .Q(
        \registers[933][6] ) );
  EDFFX1 \registers_reg[933][5]  ( .D(n8277), .E(n370), .CK(clk), .Q(
        \registers[933][5] ) );
  EDFFX1 \registers_reg[933][4]  ( .D(n8219), .E(n370), .CK(clk), .Q(
        \registers[933][4] ) );
  EDFFX1 \registers_reg[933][3]  ( .D(n8170), .E(n370), .CK(clk), .Q(
        \registers[933][3] ) );
  EDFFX1 \registers_reg[933][2]  ( .D(n8122), .E(n370), .CK(clk), .Q(
        \registers[933][2] ) );
  EDFFX1 \registers_reg[933][1]  ( .D(n8066), .E(n370), .CK(clk), .Q(
        \registers[933][1] ) );
  EDFFX1 \registers_reg[933][0]  ( .D(n8005), .E(n370), .CK(clk), .Q(
        \registers[933][0] ) );
  EDFFX1 \registers_reg[929][7]  ( .D(n8389), .E(n366), .CK(clk), .Q(
        \registers[929][7] ) );
  EDFFX1 \registers_reg[929][6]  ( .D(n8331), .E(n366), .CK(clk), .Q(
        \registers[929][6] ) );
  EDFFX1 \registers_reg[929][5]  ( .D(n8273), .E(n366), .CK(clk), .Q(
        \registers[929][5] ) );
  EDFFX1 \registers_reg[929][4]  ( .D(n8215), .E(n366), .CK(clk), .Q(
        \registers[929][4] ) );
  EDFFX1 \registers_reg[929][3]  ( .D(n8171), .E(n366), .CK(clk), .Q(
        \registers[929][3] ) );
  EDFFX1 \registers_reg[929][2]  ( .D(n8120), .E(n366), .CK(clk), .Q(
        \registers[929][2] ) );
  EDFFX1 \registers_reg[929][1]  ( .D(n8064), .E(n366), .CK(clk), .Q(
        \registers[929][1] ) );
  EDFFX1 \registers_reg[929][0]  ( .D(n8006), .E(n366), .CK(clk), .Q(
        \registers[929][0] ) );
  EDFFX1 \registers_reg[925][7]  ( .D(n8390), .E(n895), .CK(clk), .Q(
        \registers[925][7] ) );
  EDFFX1 \registers_reg[925][6]  ( .D(n8332), .E(n895), .CK(clk), .Q(
        \registers[925][6] ) );
  EDFFX1 \registers_reg[925][5]  ( .D(n8274), .E(n895), .CK(clk), .Q(
        \registers[925][5] ) );
  EDFFX1 \registers_reg[925][4]  ( .D(n8216), .E(n895), .CK(clk), .Q(
        \registers[925][4] ) );
  EDFFX1 \registers_reg[925][3]  ( .D(n8172), .E(n895), .CK(clk), .Q(
        \registers[925][3] ) );
  EDFFX1 \registers_reg[925][2]  ( .D(n8121), .E(n895), .CK(clk), .Q(
        \registers[925][2] ) );
  EDFFX1 \registers_reg[925][1]  ( .D(n8065), .E(n895), .CK(clk), .Q(
        \registers[925][1] ) );
  EDFFX1 \registers_reg[925][0]  ( .D(n8004), .E(n895), .CK(clk), .Q(
        \registers[925][0] ) );
  EDFFX1 \registers_reg[921][7]  ( .D(n8391), .E(n891), .CK(clk), .Q(
        \registers[921][7] ) );
  EDFFX1 \registers_reg[921][6]  ( .D(n8333), .E(n891), .CK(clk), .Q(
        \registers[921][6] ) );
  EDFFX1 \registers_reg[921][5]  ( .D(n8275), .E(n891), .CK(clk), .Q(
        \registers[921][5] ) );
  EDFFX1 \registers_reg[921][4]  ( .D(n8217), .E(n891), .CK(clk), .Q(
        \registers[921][4] ) );
  EDFFX1 \registers_reg[921][3]  ( .D(n8170), .E(n891), .CK(clk), .Q(
        \registers[921][3] ) );
  EDFFX1 \registers_reg[921][2]  ( .D(n8122), .E(n891), .CK(clk), .Q(
        \registers[921][2] ) );
  EDFFX1 \registers_reg[921][1]  ( .D(n8066), .E(n891), .CK(clk), .Q(
        \registers[921][1] ) );
  EDFFX1 \registers_reg[921][0]  ( .D(n8005), .E(n891), .CK(clk), .Q(
        \registers[921][0] ) );
  EDFFX1 \registers_reg[917][7]  ( .D(n8389), .E(n887), .CK(clk), .Q(
        \registers[917][7] ) );
  EDFFX1 \registers_reg[917][6]  ( .D(n8331), .E(n887), .CK(clk), .Q(
        \registers[917][6] ) );
  EDFFX1 \registers_reg[917][5]  ( .D(n8273), .E(n887), .CK(clk), .Q(
        \registers[917][5] ) );
  EDFFX1 \registers_reg[917][4]  ( .D(n8215), .E(n887), .CK(clk), .Q(
        \registers[917][4] ) );
  EDFFX1 \registers_reg[917][3]  ( .D(n8171), .E(n887), .CK(clk), .Q(
        \registers[917][3] ) );
  EDFFX1 \registers_reg[917][2]  ( .D(n8120), .E(n887), .CK(clk), .Q(
        \registers[917][2] ) );
  EDFFX1 \registers_reg[917][1]  ( .D(n8064), .E(n887), .CK(clk), .Q(
        \registers[917][1] ) );
  EDFFX1 \registers_reg[917][0]  ( .D(n8006), .E(n887), .CK(clk), .Q(
        \registers[917][0] ) );
  EDFFX1 \registers_reg[913][7]  ( .D(n8390), .E(n200), .CK(clk), .Q(
        \registers[913][7] ) );
  EDFFX1 \registers_reg[913][6]  ( .D(n8332), .E(n200), .CK(clk), .Q(
        \registers[913][6] ) );
  EDFFX1 \registers_reg[913][5]  ( .D(n8274), .E(n200), .CK(clk), .Q(
        \registers[913][5] ) );
  EDFFX1 \registers_reg[913][4]  ( .D(n8216), .E(n200), .CK(clk), .Q(
        \registers[913][4] ) );
  EDFFX1 \registers_reg[913][3]  ( .D(n8172), .E(n200), .CK(clk), .Q(
        \registers[913][3] ) );
  EDFFX1 \registers_reg[913][2]  ( .D(n8121), .E(n200), .CK(clk), .Q(
        \registers[913][2] ) );
  EDFFX1 \registers_reg[913][1]  ( .D(n8065), .E(n200), .CK(clk), .Q(
        \registers[913][1] ) );
  EDFFX1 \registers_reg[913][0]  ( .D(n8004), .E(n200), .CK(clk), .Q(
        \registers[913][0] ) );
  EDFFX1 \registers_reg[909][7]  ( .D(n8391), .E(n196), .CK(clk), .Q(
        \registers[909][7] ) );
  EDFFX1 \registers_reg[909][6]  ( .D(n8333), .E(n196), .CK(clk), .Q(
        \registers[909][6] ) );
  EDFFX1 \registers_reg[909][5]  ( .D(n8275), .E(n196), .CK(clk), .Q(
        \registers[909][5] ) );
  EDFFX1 \registers_reg[909][4]  ( .D(n8217), .E(n196), .CK(clk), .Q(
        \registers[909][4] ) );
  EDFFX1 \registers_reg[909][3]  ( .D(n8170), .E(n196), .CK(clk), .Q(
        \registers[909][3] ) );
  EDFFX1 \registers_reg[909][2]  ( .D(n8122), .E(n196), .CK(clk), .Q(
        \registers[909][2] ) );
  EDFFX1 \registers_reg[909][1]  ( .D(n8066), .E(n196), .CK(clk), .Q(
        \registers[909][1] ) );
  EDFFX1 \registers_reg[909][0]  ( .D(n8005), .E(n196), .CK(clk), .Q(
        \registers[909][0] ) );
  EDFFX1 \registers_reg[905][7]  ( .D(n8389), .E(n192), .CK(clk), .Q(
        \registers[905][7] ) );
  EDFFX1 \registers_reg[905][6]  ( .D(n8331), .E(n192), .CK(clk), .Q(
        \registers[905][6] ) );
  EDFFX1 \registers_reg[905][5]  ( .D(n8273), .E(n192), .CK(clk), .Q(
        \registers[905][5] ) );
  EDFFX1 \registers_reg[905][4]  ( .D(n8215), .E(n192), .CK(clk), .Q(
        \registers[905][4] ) );
  EDFFX1 \registers_reg[905][3]  ( .D(n8171), .E(n192), .CK(clk), .Q(
        \registers[905][3] ) );
  EDFFX1 \registers_reg[905][2]  ( .D(n8120), .E(n192), .CK(clk), .Q(
        \registers[905][2] ) );
  EDFFX1 \registers_reg[905][1]  ( .D(n8064), .E(n192), .CK(clk), .Q(
        \registers[905][1] ) );
  EDFFX1 \registers_reg[905][0]  ( .D(n8006), .E(n192), .CK(clk), .Q(
        \registers[905][0] ) );
  EDFFX1 \registers_reg[901][7]  ( .D(n8390), .E(n363), .CK(clk), .Q(
        \registers[901][7] ) );
  EDFFX1 \registers_reg[901][6]  ( .D(n8332), .E(n363), .CK(clk), .Q(
        \registers[901][6] ) );
  EDFFX1 \registers_reg[901][5]  ( .D(n8274), .E(n363), .CK(clk), .Q(
        \registers[901][5] ) );
  EDFFX1 \registers_reg[901][4]  ( .D(n8216), .E(n363), .CK(clk), .Q(
        \registers[901][4] ) );
  EDFFX1 \registers_reg[901][3]  ( .D(n8172), .E(n363), .CK(clk), .Q(
        \registers[901][3] ) );
  EDFFX1 \registers_reg[901][2]  ( .D(n8121), .E(n363), .CK(clk), .Q(
        \registers[901][2] ) );
  EDFFX1 \registers_reg[901][1]  ( .D(n8065), .E(n363), .CK(clk), .Q(
        \registers[901][1] ) );
  EDFFX1 \registers_reg[901][0]  ( .D(n8004), .E(n363), .CK(clk), .Q(
        \registers[901][0] ) );
  EDFFX1 \registers_reg[897][7]  ( .D(n8391), .E(n359), .CK(clk), .Q(
        \registers[897][7] ) );
  EDFFX1 \registers_reg[897][6]  ( .D(n8333), .E(n359), .CK(clk), .Q(
        \registers[897][6] ) );
  EDFFX1 \registers_reg[897][5]  ( .D(n8275), .E(n359), .CK(clk), .Q(
        \registers[897][5] ) );
  EDFFX1 \registers_reg[897][4]  ( .D(n8217), .E(n359), .CK(clk), .Q(
        \registers[897][4] ) );
  EDFFX1 \registers_reg[897][3]  ( .D(n8170), .E(n359), .CK(clk), .Q(
        \registers[897][3] ) );
  EDFFX1 \registers_reg[897][2]  ( .D(n8122), .E(n359), .CK(clk), .Q(
        \registers[897][2] ) );
  EDFFX1 \registers_reg[897][1]  ( .D(n8066), .E(n359), .CK(clk), .Q(
        \registers[897][1] ) );
  EDFFX1 \registers_reg[897][0]  ( .D(n8005), .E(n359), .CK(clk), .Q(
        \registers[897][0] ) );
  EDFFX1 \registers_reg[893][7]  ( .D(n8404), .E(n883), .CK(clk), .Q(
        \registers[893][7] ) );
  EDFFX1 \registers_reg[893][6]  ( .D(n8346), .E(n883), .CK(clk), .Q(
        \registers[893][6] ) );
  EDFFX1 \registers_reg[893][5]  ( .D(n8288), .E(n883), .CK(clk), .Q(
        \registers[893][5] ) );
  EDFFX1 \registers_reg[893][4]  ( .D(n8230), .E(n883), .CK(clk), .Q(
        \registers[893][4] ) );
  EDFFX1 \registers_reg[893][3]  ( .D(n8182), .E(n883), .CK(clk), .Q(
        \registers[893][3] ) );
  EDFFX1 \registers_reg[893][2]  ( .D(n8137), .E(n883), .CK(clk), .Q(
        \registers[893][2] ) );
  EDFFX1 \registers_reg[893][1]  ( .D(n8081), .E(n883), .CK(clk), .Q(
        \registers[893][1] ) );
  EDFFX1 \registers_reg[893][0]  ( .D(n8020), .E(n883), .CK(clk), .Q(
        \registers[893][0] ) );
  EDFFX1 \registers_reg[889][7]  ( .D(n8405), .E(n879), .CK(clk), .Q(
        \registers[889][7] ) );
  EDFFX1 \registers_reg[889][6]  ( .D(n8347), .E(n879), .CK(clk), .Q(
        \registers[889][6] ) );
  EDFFX1 \registers_reg[889][5]  ( .D(n8289), .E(n879), .CK(clk), .Q(
        \registers[889][5] ) );
  EDFFX1 \registers_reg[889][4]  ( .D(n8231), .E(n879), .CK(clk), .Q(
        \registers[889][4] ) );
  EDFFX1 \registers_reg[889][3]  ( .D(n8183), .E(n879), .CK(clk), .Q(
        \registers[889][3] ) );
  EDFFX1 \registers_reg[889][2]  ( .D(n8135), .E(n879), .CK(clk), .Q(
        \registers[889][2] ) );
  EDFFX1 \registers_reg[889][1]  ( .D(n8079), .E(n879), .CK(clk), .Q(
        \registers[889][1] ) );
  EDFFX1 \registers_reg[889][0]  ( .D(n8021), .E(n879), .CK(clk), .Q(
        \registers[889][0] ) );
  EDFFX1 \registers_reg[885][7]  ( .D(n8406), .E(n875), .CK(clk), .Q(
        \registers[885][7] ) );
  EDFFX1 \registers_reg[885][6]  ( .D(n8348), .E(n875), .CK(clk), .Q(
        \registers[885][6] ) );
  EDFFX1 \registers_reg[885][5]  ( .D(n8290), .E(n875), .CK(clk), .Q(
        \registers[885][5] ) );
  EDFFX1 \registers_reg[885][4]  ( .D(n8232), .E(n875), .CK(clk), .Q(
        \registers[885][4] ) );
  EDFFX1 \registers_reg[885][3]  ( .D(n8184), .E(n875), .CK(clk), .Q(
        \registers[885][3] ) );
  EDFFX1 \registers_reg[885][2]  ( .D(n8136), .E(n875), .CK(clk), .Q(
        \registers[885][2] ) );
  EDFFX1 \registers_reg[885][1]  ( .D(n8080), .E(n875), .CK(clk), .Q(
        \registers[885][1] ) );
  EDFFX1 \registers_reg[885][0]  ( .D(n8019), .E(n875), .CK(clk), .Q(
        \registers[885][0] ) );
  EDFFX1 \registers_reg[881][7]  ( .D(n8404), .E(n188), .CK(clk), .Q(
        \registers[881][7] ) );
  EDFFX1 \registers_reg[881][6]  ( .D(n8346), .E(n188), .CK(clk), .Q(
        \registers[881][6] ) );
  EDFFX1 \registers_reg[881][5]  ( .D(n8288), .E(n188), .CK(clk), .Q(
        \registers[881][5] ) );
  EDFFX1 \registers_reg[881][4]  ( .D(n8230), .E(n188), .CK(clk), .Q(
        \registers[881][4] ) );
  EDFFX1 \registers_reg[881][3]  ( .D(n8182), .E(n188), .CK(clk), .Q(
        \registers[881][3] ) );
  EDFFX1 \registers_reg[881][2]  ( .D(n8134), .E(n188), .CK(clk), .Q(
        \registers[881][2] ) );
  EDFFX1 \registers_reg[881][1]  ( .D(n8078), .E(n188), .CK(clk), .Q(
        \registers[881][1] ) );
  EDFFX1 \registers_reg[881][0]  ( .D(n8017), .E(n188), .CK(clk), .Q(
        \registers[881][0] ) );
  EDFFX1 \registers_reg[877][7]  ( .D(n8405), .E(n184), .CK(clk), .Q(
        \registers[877][7] ) );
  EDFFX1 \registers_reg[877][6]  ( .D(n8347), .E(n184), .CK(clk), .Q(
        \registers[877][6] ) );
  EDFFX1 \registers_reg[877][5]  ( .D(n8289), .E(n184), .CK(clk), .Q(
        \registers[877][5] ) );
  EDFFX1 \registers_reg[877][4]  ( .D(n8231), .E(n184), .CK(clk), .Q(
        \registers[877][4] ) );
  EDFFX1 \registers_reg[877][3]  ( .D(n8183), .E(n184), .CK(clk), .Q(
        \registers[877][3] ) );
  EDFFX1 \registers_reg[877][2]  ( .D(n8132), .E(n184), .CK(clk), .Q(
        \registers[877][2] ) );
  EDFFX1 \registers_reg[877][1]  ( .D(n8076), .E(n184), .CK(clk), .Q(
        \registers[877][1] ) );
  EDFFX1 \registers_reg[877][0]  ( .D(n8018), .E(n184), .CK(clk), .Q(
        \registers[877][0] ) );
  EDFFX1 \registers_reg[873][7]  ( .D(n8401), .E(n180), .CK(clk), .Q(
        \registers[873][7] ) );
  EDFFX1 \registers_reg[873][6]  ( .D(n8343), .E(n180), .CK(clk), .Q(
        \registers[873][6] ) );
  EDFFX1 \registers_reg[873][5]  ( .D(n8285), .E(n180), .CK(clk), .Q(
        \registers[873][5] ) );
  EDFFX1 \registers_reg[873][4]  ( .D(n8227), .E(n180), .CK(clk), .Q(
        \registers[873][4] ) );
  EDFFX1 \registers_reg[873][3]  ( .D(n8181), .E(n180), .CK(clk), .Q(
        \registers[873][3] ) );
  EDFFX1 \registers_reg[873][2]  ( .D(n8133), .E(n180), .CK(clk), .Q(
        \registers[873][2] ) );
  EDFFX1 \registers_reg[873][1]  ( .D(n8077), .E(n180), .CK(clk), .Q(
        \registers[873][1] ) );
  EDFFX1 \registers_reg[873][0]  ( .D(n8016), .E(n180), .CK(clk), .Q(
        \registers[873][0] ) );
  EDFFX1 \registers_reg[869][7]  ( .D(n8402), .E(n356), .CK(clk), .Q(
        \registers[869][7] ) );
  EDFFX1 \registers_reg[869][6]  ( .D(n8344), .E(n356), .CK(clk), .Q(
        \registers[869][6] ) );
  EDFFX1 \registers_reg[869][5]  ( .D(n8286), .E(n356), .CK(clk), .Q(
        \registers[869][5] ) );
  EDFFX1 \registers_reg[869][4]  ( .D(n8228), .E(n356), .CK(clk), .Q(
        \registers[869][4] ) );
  EDFFX1 \registers_reg[869][3]  ( .D(n8179), .E(n356), .CK(clk), .Q(
        \registers[869][3] ) );
  EDFFX1 \registers_reg[869][2]  ( .D(n8134), .E(n356), .CK(clk), .Q(
        \registers[869][2] ) );
  EDFFX1 \registers_reg[869][1]  ( .D(n8078), .E(n356), .CK(clk), .Q(
        \registers[869][1] ) );
  EDFFX1 \registers_reg[869][0]  ( .D(n8017), .E(n356), .CK(clk), .Q(
        \registers[869][0] ) );
  EDFFX1 \registers_reg[865][7]  ( .D(n8403), .E(n352), .CK(clk), .Q(
        \registers[865][7] ) );
  EDFFX1 \registers_reg[865][6]  ( .D(n8345), .E(n352), .CK(clk), .Q(
        \registers[865][6] ) );
  EDFFX1 \registers_reg[865][5]  ( .D(n8287), .E(n352), .CK(clk), .Q(
        \registers[865][5] ) );
  EDFFX1 \registers_reg[865][4]  ( .D(n8229), .E(n352), .CK(clk), .Q(
        \registers[865][4] ) );
  EDFFX1 \registers_reg[865][3]  ( .D(n8180), .E(n352), .CK(clk), .Q(
        \registers[865][3] ) );
  EDFFX1 \registers_reg[865][2]  ( .D(n8132), .E(n352), .CK(clk), .Q(
        \registers[865][2] ) );
  EDFFX1 \registers_reg[865][1]  ( .D(n8076), .E(n352), .CK(clk), .Q(
        \registers[865][1] ) );
  EDFFX1 \registers_reg[865][0]  ( .D(n8018), .E(n352), .CK(clk), .Q(
        \registers[865][0] ) );
  EDFFX1 \registers_reg[861][7]  ( .D(n8401), .E(n871), .CK(clk), .Q(
        \registers[861][7] ) );
  EDFFX1 \registers_reg[861][6]  ( .D(n8343), .E(n871), .CK(clk), .Q(
        \registers[861][6] ) );
  EDFFX1 \registers_reg[861][5]  ( .D(n8285), .E(n871), .CK(clk), .Q(
        \registers[861][5] ) );
  EDFFX1 \registers_reg[861][4]  ( .D(n8227), .E(n871), .CK(clk), .Q(
        \registers[861][4] ) );
  EDFFX1 \registers_reg[861][3]  ( .D(n8181), .E(n871), .CK(clk), .Q(
        \registers[861][3] ) );
  EDFFX1 \registers_reg[861][2]  ( .D(n8133), .E(n871), .CK(clk), .Q(
        \registers[861][2] ) );
  EDFFX1 \registers_reg[861][1]  ( .D(n8077), .E(n871), .CK(clk), .Q(
        \registers[861][1] ) );
  EDFFX1 \registers_reg[861][0]  ( .D(n8016), .E(n871), .CK(clk), .Q(
        \registers[861][0] ) );
  EDFFX1 \registers_reg[857][7]  ( .D(n8402), .E(n867), .CK(clk), .Q(
        \registers[857][7] ) );
  EDFFX1 \registers_reg[857][6]  ( .D(n8344), .E(n867), .CK(clk), .Q(
        \registers[857][6] ) );
  EDFFX1 \registers_reg[857][5]  ( .D(n8286), .E(n867), .CK(clk), .Q(
        \registers[857][5] ) );
  EDFFX1 \registers_reg[857][4]  ( .D(n8228), .E(n867), .CK(clk), .Q(
        \registers[857][4] ) );
  EDFFX1 \registers_reg[857][3]  ( .D(n8179), .E(n867), .CK(clk), .Q(
        \registers[857][3] ) );
  EDFFX1 \registers_reg[857][2]  ( .D(n8134), .E(n867), .CK(clk), .Q(
        \registers[857][2] ) );
  EDFFX1 \registers_reg[857][1]  ( .D(n8078), .E(n867), .CK(clk), .Q(
        \registers[857][1] ) );
  EDFFX1 \registers_reg[857][0]  ( .D(n8017), .E(n867), .CK(clk), .Q(
        \registers[857][0] ) );
  EDFFX1 \registers_reg[853][7]  ( .D(n8403), .E(n863), .CK(clk), .Q(
        \registers[853][7] ) );
  EDFFX1 \registers_reg[853][6]  ( .D(n8345), .E(n863), .CK(clk), .Q(
        \registers[853][6] ) );
  EDFFX1 \registers_reg[853][5]  ( .D(n8287), .E(n863), .CK(clk), .Q(
        \registers[853][5] ) );
  EDFFX1 \registers_reg[853][4]  ( .D(n8229), .E(n863), .CK(clk), .Q(
        \registers[853][4] ) );
  EDFFX1 \registers_reg[853][3]  ( .D(n8180), .E(n863), .CK(clk), .Q(
        \registers[853][3] ) );
  EDFFX1 \registers_reg[853][2]  ( .D(n8132), .E(n863), .CK(clk), .Q(
        \registers[853][2] ) );
  EDFFX1 \registers_reg[853][1]  ( .D(n8076), .E(n863), .CK(clk), .Q(
        \registers[853][1] ) );
  EDFFX1 \registers_reg[853][0]  ( .D(n8018), .E(n863), .CK(clk), .Q(
        \registers[853][0] ) );
  EDFFX1 \registers_reg[849][7]  ( .D(n8401), .E(n176), .CK(clk), .Q(
        \registers[849][7] ) );
  EDFFX1 \registers_reg[849][6]  ( .D(n8343), .E(n176), .CK(clk), .Q(
        \registers[849][6] ) );
  EDFFX1 \registers_reg[849][5]  ( .D(n8285), .E(n176), .CK(clk), .Q(
        \registers[849][5] ) );
  EDFFX1 \registers_reg[849][4]  ( .D(n8227), .E(n176), .CK(clk), .Q(
        \registers[849][4] ) );
  EDFFX1 \registers_reg[849][3]  ( .D(n8181), .E(n176), .CK(clk), .Q(
        \registers[849][3] ) );
  EDFFX1 \registers_reg[849][2]  ( .D(n8133), .E(n176), .CK(clk), .Q(
        \registers[849][2] ) );
  EDFFX1 \registers_reg[849][1]  ( .D(n8077), .E(n176), .CK(clk), .Q(
        \registers[849][1] ) );
  EDFFX1 \registers_reg[849][0]  ( .D(n8016), .E(n176), .CK(clk), .Q(
        \registers[849][0] ) );
  EDFFX1 \registers_reg[845][7]  ( .D(n8402), .E(n172), .CK(clk), .Q(
        \registers[845][7] ) );
  EDFFX1 \registers_reg[845][6]  ( .D(n8344), .E(n172), .CK(clk), .Q(
        \registers[845][6] ) );
  EDFFX1 \registers_reg[845][5]  ( .D(n8286), .E(n172), .CK(clk), .Q(
        \registers[845][5] ) );
  EDFFX1 \registers_reg[845][4]  ( .D(n8228), .E(n172), .CK(clk), .Q(
        \registers[845][4] ) );
  EDFFX1 \registers_reg[845][3]  ( .D(n8179), .E(n172), .CK(clk), .Q(
        \registers[845][3] ) );
  EDFFX1 \registers_reg[845][2]  ( .D(n8134), .E(n172), .CK(clk), .Q(
        \registers[845][2] ) );
  EDFFX1 \registers_reg[845][1]  ( .D(n8078), .E(n172), .CK(clk), .Q(
        \registers[845][1] ) );
  EDFFX1 \registers_reg[845][0]  ( .D(n8017), .E(n172), .CK(clk), .Q(
        \registers[845][0] ) );
  EDFFX1 \registers_reg[841][7]  ( .D(n8403), .E(n168), .CK(clk), .Q(
        \registers[841][7] ) );
  EDFFX1 \registers_reg[841][6]  ( .D(n8345), .E(n168), .CK(clk), .Q(
        \registers[841][6] ) );
  EDFFX1 \registers_reg[841][5]  ( .D(n8287), .E(n168), .CK(clk), .Q(
        \registers[841][5] ) );
  EDFFX1 \registers_reg[841][4]  ( .D(n8229), .E(n168), .CK(clk), .Q(
        \registers[841][4] ) );
  EDFFX1 \registers_reg[841][3]  ( .D(n8180), .E(n168), .CK(clk), .Q(
        \registers[841][3] ) );
  EDFFX1 \registers_reg[841][2]  ( .D(n8132), .E(n168), .CK(clk), .Q(
        \registers[841][2] ) );
  EDFFX1 \registers_reg[841][1]  ( .D(n8076), .E(n168), .CK(clk), .Q(
        \registers[841][1] ) );
  EDFFX1 \registers_reg[841][0]  ( .D(n8018), .E(n168), .CK(clk), .Q(
        \registers[841][0] ) );
  EDFFX1 \registers_reg[837][7]  ( .D(n8401), .E(n349), .CK(clk), .Q(
        \registers[837][7] ) );
  EDFFX1 \registers_reg[837][6]  ( .D(n8343), .E(n349), .CK(clk), .Q(
        \registers[837][6] ) );
  EDFFX1 \registers_reg[837][5]  ( .D(n8285), .E(n349), .CK(clk), .Q(
        \registers[837][5] ) );
  EDFFX1 \registers_reg[837][4]  ( .D(n8227), .E(n349), .CK(clk), .Q(
        \registers[837][4] ) );
  EDFFX1 \registers_reg[837][3]  ( .D(n8181), .E(n349), .CK(clk), .Q(
        \registers[837][3] ) );
  EDFFX1 \registers_reg[837][2]  ( .D(n8133), .E(n349), .CK(clk), .Q(
        \registers[837][2] ) );
  EDFFX1 \registers_reg[837][1]  ( .D(n8077), .E(n349), .CK(clk), .Q(
        \registers[837][1] ) );
  EDFFX1 \registers_reg[837][0]  ( .D(n8016), .E(n349), .CK(clk), .Q(
        \registers[837][0] ) );
  EDFFX1 \registers_reg[833][7]  ( .D(n8402), .E(n345), .CK(clk), .Q(
        \registers[833][7] ) );
  EDFFX1 \registers_reg[833][6]  ( .D(n8344), .E(n345), .CK(clk), .Q(
        \registers[833][6] ) );
  EDFFX1 \registers_reg[833][5]  ( .D(n8286), .E(n345), .CK(clk), .Q(
        \registers[833][5] ) );
  EDFFX1 \registers_reg[833][4]  ( .D(n8228), .E(n345), .CK(clk), .Q(
        \registers[833][4] ) );
  EDFFX1 \registers_reg[833][3]  ( .D(n8179), .E(n345), .CK(clk), .Q(
        \registers[833][3] ) );
  EDFFX1 \registers_reg[833][2]  ( .D(n8134), .E(n345), .CK(clk), .Q(
        \registers[833][2] ) );
  EDFFX1 \registers_reg[833][1]  ( .D(n8078), .E(n345), .CK(clk), .Q(
        \registers[833][1] ) );
  EDFFX1 \registers_reg[833][0]  ( .D(n8017), .E(n345), .CK(clk), .Q(
        \registers[833][0] ) );
  EDFFX1 \registers_reg[829][7]  ( .D(n8401), .E(n859), .CK(clk), .Q(
        \registers[829][7] ) );
  EDFFX1 \registers_reg[829][6]  ( .D(n8343), .E(n859), .CK(clk), .Q(
        \registers[829][6] ) );
  EDFFX1 \registers_reg[829][5]  ( .D(n8285), .E(n859), .CK(clk), .Q(
        \registers[829][5] ) );
  EDFFX1 \registers_reg[829][4]  ( .D(n8227), .E(n859), .CK(clk), .Q(
        \registers[829][4] ) );
  EDFFX1 \registers_reg[829][3]  ( .D(n8181), .E(n859), .CK(clk), .Q(
        \registers[829][3] ) );
  EDFFX1 \registers_reg[829][2]  ( .D(n8130), .E(n859), .CK(clk), .Q(
        \registers[829][2] ) );
  EDFFX1 \registers_reg[829][1]  ( .D(n8074), .E(n859), .CK(clk), .Q(
        \registers[829][1] ) );
  EDFFX1 \registers_reg[829][0]  ( .D(n8013), .E(n859), .CK(clk), .Q(
        \registers[829][0] ) );
  EDFFX1 \registers_reg[825][7]  ( .D(n8402), .E(n855), .CK(clk), .Q(
        \registers[825][7] ) );
  EDFFX1 \registers_reg[825][6]  ( .D(n8344), .E(n855), .CK(clk), .Q(
        \registers[825][6] ) );
  EDFFX1 \registers_reg[825][5]  ( .D(n8286), .E(n855), .CK(clk), .Q(
        \registers[825][5] ) );
  EDFFX1 \registers_reg[825][4]  ( .D(n8228), .E(n855), .CK(clk), .Q(
        \registers[825][4] ) );
  EDFFX1 \registers_reg[825][3]  ( .D(n8179), .E(n855), .CK(clk), .Q(
        \registers[825][3] ) );
  EDFFX1 \registers_reg[825][2]  ( .D(n8131), .E(n855), .CK(clk), .Q(
        \registers[825][2] ) );
  EDFFX1 \registers_reg[825][1]  ( .D(n8075), .E(n855), .CK(clk), .Q(
        \registers[825][1] ) );
  EDFFX1 \registers_reg[825][0]  ( .D(n8014), .E(n855), .CK(clk), .Q(
        \registers[825][0] ) );
  EDFFX1 \registers_reg[821][7]  ( .D(n8398), .E(n851), .CK(clk), .Q(
        \registers[821][7] ) );
  EDFFX1 \registers_reg[821][6]  ( .D(n8340), .E(n851), .CK(clk), .Q(
        \registers[821][6] ) );
  EDFFX1 \registers_reg[821][5]  ( .D(n8282), .E(n851), .CK(clk), .Q(
        \registers[821][5] ) );
  EDFFX1 \registers_reg[821][4]  ( .D(n8224), .E(n851), .CK(clk), .Q(
        \registers[821][4] ) );
  EDFFX1 \registers_reg[821][3]  ( .D(n8180), .E(n851), .CK(clk), .Q(
        \registers[821][3] ) );
  EDFFX1 \registers_reg[821][2]  ( .D(n8129), .E(n851), .CK(clk), .Q(
        \registers[821][2] ) );
  EDFFX1 \registers_reg[821][1]  ( .D(n8073), .E(n851), .CK(clk), .Q(
        \registers[821][1] ) );
  EDFFX1 \registers_reg[821][0]  ( .D(n8015), .E(n851), .CK(clk), .Q(
        \registers[821][0] ) );
  EDFFX1 \registers_reg[817][7]  ( .D(n8399), .E(n164), .CK(clk), .Q(
        \registers[817][7] ) );
  EDFFX1 \registers_reg[817][6]  ( .D(n8341), .E(n164), .CK(clk), .Q(
        \registers[817][6] ) );
  EDFFX1 \registers_reg[817][5]  ( .D(n8283), .E(n164), .CK(clk), .Q(
        \registers[817][5] ) );
  EDFFX1 \registers_reg[817][4]  ( .D(n8225), .E(n164), .CK(clk), .Q(
        \registers[817][4] ) );
  EDFFX1 \registers_reg[817][3]  ( .D(n8181), .E(n164), .CK(clk), .Q(
        \registers[817][3] ) );
  EDFFX1 \registers_reg[817][2]  ( .D(n8130), .E(n164), .CK(clk), .Q(
        \registers[817][2] ) );
  EDFFX1 \registers_reg[817][1]  ( .D(n8074), .E(n164), .CK(clk), .Q(
        \registers[817][1] ) );
  EDFFX1 \registers_reg[817][0]  ( .D(n8013), .E(n164), .CK(clk), .Q(
        \registers[817][0] ) );
  EDFFX1 \registers_reg[813][7]  ( .D(n8400), .E(n160), .CK(clk), .Q(
        \registers[813][7] ) );
  EDFFX1 \registers_reg[813][6]  ( .D(n8342), .E(n160), .CK(clk), .Q(
        \registers[813][6] ) );
  EDFFX1 \registers_reg[813][5]  ( .D(n8284), .E(n160), .CK(clk), .Q(
        \registers[813][5] ) );
  EDFFX1 \registers_reg[813][4]  ( .D(n8226), .E(n160), .CK(clk), .Q(
        \registers[813][4] ) );
  EDFFX1 \registers_reg[813][3]  ( .D(n8176), .E(n160), .CK(clk), .Q(
        \registers[813][3] ) );
  EDFFX1 \registers_reg[813][2]  ( .D(n8131), .E(n160), .CK(clk), .Q(
        \registers[813][2] ) );
  EDFFX1 \registers_reg[813][1]  ( .D(n8075), .E(n160), .CK(clk), .Q(
        \registers[813][1] ) );
  EDFFX1 \registers_reg[813][0]  ( .D(n8014), .E(n160), .CK(clk), .Q(
        \registers[813][0] ) );
  EDFFX1 \registers_reg[809][7]  ( .D(n8398), .E(n156), .CK(clk), .Q(
        \registers[809][7] ) );
  EDFFX1 \registers_reg[809][6]  ( .D(n8340), .E(n156), .CK(clk), .Q(
        \registers[809][6] ) );
  EDFFX1 \registers_reg[809][5]  ( .D(n8282), .E(n156), .CK(clk), .Q(
        \registers[809][5] ) );
  EDFFX1 \registers_reg[809][4]  ( .D(n8224), .E(n156), .CK(clk), .Q(
        \registers[809][4] ) );
  EDFFX1 \registers_reg[809][3]  ( .D(n8177), .E(n156), .CK(clk), .Q(
        \registers[809][3] ) );
  EDFFX1 \registers_reg[809][2]  ( .D(n8129), .E(n156), .CK(clk), .Q(
        \registers[809][2] ) );
  EDFFX1 \registers_reg[809][1]  ( .D(n8073), .E(n156), .CK(clk), .Q(
        \registers[809][1] ) );
  EDFFX1 \registers_reg[809][0]  ( .D(n8015), .E(n156), .CK(clk), .Q(
        \registers[809][0] ) );
  EDFFX1 \registers_reg[805][7]  ( .D(n8399), .E(n327), .CK(clk), .Q(
        \registers[805][7] ) );
  EDFFX1 \registers_reg[805][6]  ( .D(n8341), .E(n327), .CK(clk), .Q(
        \registers[805][6] ) );
  EDFFX1 \registers_reg[805][5]  ( .D(n8283), .E(n327), .CK(clk), .Q(
        \registers[805][5] ) );
  EDFFX1 \registers_reg[805][4]  ( .D(n8225), .E(n327), .CK(clk), .Q(
        \registers[805][4] ) );
  EDFFX1 \registers_reg[805][3]  ( .D(n8178), .E(n327), .CK(clk), .Q(
        \registers[805][3] ) );
  EDFFX1 \registers_reg[805][2]  ( .D(n8130), .E(n327), .CK(clk), .Q(
        \registers[805][2] ) );
  EDFFX1 \registers_reg[805][1]  ( .D(n8074), .E(n327), .CK(clk), .Q(
        \registers[805][1] ) );
  EDFFX1 \registers_reg[805][0]  ( .D(n8013), .E(n327), .CK(clk), .Q(
        \registers[805][0] ) );
  EDFFX1 \registers_reg[801][7]  ( .D(n8400), .E(n323), .CK(clk), .Q(
        \registers[801][7] ) );
  EDFFX1 \registers_reg[801][6]  ( .D(n8342), .E(n323), .CK(clk), .Q(
        \registers[801][6] ) );
  EDFFX1 \registers_reg[801][5]  ( .D(n8284), .E(n323), .CK(clk), .Q(
        \registers[801][5] ) );
  EDFFX1 \registers_reg[801][4]  ( .D(n8226), .E(n323), .CK(clk), .Q(
        \registers[801][4] ) );
  EDFFX1 \registers_reg[801][3]  ( .D(n8176), .E(n323), .CK(clk), .Q(
        \registers[801][3] ) );
  EDFFX1 \registers_reg[801][2]  ( .D(n8131), .E(n323), .CK(clk), .Q(
        \registers[801][2] ) );
  EDFFX1 \registers_reg[801][1]  ( .D(n8075), .E(n323), .CK(clk), .Q(
        \registers[801][1] ) );
  EDFFX1 \registers_reg[801][0]  ( .D(n8014), .E(n323), .CK(clk), .Q(
        \registers[801][0] ) );
  EDFFX1 \registers_reg[797][7]  ( .D(n8398), .E(n847), .CK(clk), .Q(
        \registers[797][7] ) );
  EDFFX1 \registers_reg[797][6]  ( .D(n8340), .E(n847), .CK(clk), .Q(
        \registers[797][6] ) );
  EDFFX1 \registers_reg[797][5]  ( .D(n8282), .E(n847), .CK(clk), .Q(
        \registers[797][5] ) );
  EDFFX1 \registers_reg[797][4]  ( .D(n8224), .E(n847), .CK(clk), .Q(
        \registers[797][4] ) );
  EDFFX1 \registers_reg[797][3]  ( .D(n8177), .E(n847), .CK(clk), .Q(
        \registers[797][3] ) );
  EDFFX1 \registers_reg[797][2]  ( .D(n8129), .E(n847), .CK(clk), .Q(
        \registers[797][2] ) );
  EDFFX1 \registers_reg[797][1]  ( .D(n8073), .E(n847), .CK(clk), .Q(
        \registers[797][1] ) );
  EDFFX1 \registers_reg[797][0]  ( .D(n8015), .E(n847), .CK(clk), .Q(
        \registers[797][0] ) );
  EDFFX1 \registers_reg[793][7]  ( .D(n8399), .E(n843), .CK(clk), .Q(
        \registers[793][7] ) );
  EDFFX1 \registers_reg[793][6]  ( .D(n8341), .E(n843), .CK(clk), .Q(
        \registers[793][6] ) );
  EDFFX1 \registers_reg[793][5]  ( .D(n8283), .E(n843), .CK(clk), .Q(
        \registers[793][5] ) );
  EDFFX1 \registers_reg[793][4]  ( .D(n8225), .E(n843), .CK(clk), .Q(
        \registers[793][4] ) );
  EDFFX1 \registers_reg[793][3]  ( .D(n8178), .E(n843), .CK(clk), .Q(
        \registers[793][3] ) );
  EDFFX1 \registers_reg[793][2]  ( .D(n8130), .E(n843), .CK(clk), .Q(
        \registers[793][2] ) );
  EDFFX1 \registers_reg[793][1]  ( .D(n8074), .E(n843), .CK(clk), .Q(
        \registers[793][1] ) );
  EDFFX1 \registers_reg[793][0]  ( .D(n8013), .E(n843), .CK(clk), .Q(
        \registers[793][0] ) );
  EDFFX1 \registers_reg[789][7]  ( .D(n8400), .E(n839), .CK(clk), .Q(
        \registers[789][7] ) );
  EDFFX1 \registers_reg[789][6]  ( .D(n8342), .E(n839), .CK(clk), .Q(
        \registers[789][6] ) );
  EDFFX1 \registers_reg[789][5]  ( .D(n8284), .E(n839), .CK(clk), .Q(
        \registers[789][5] ) );
  EDFFX1 \registers_reg[789][4]  ( .D(n8226), .E(n839), .CK(clk), .Q(
        \registers[789][4] ) );
  EDFFX1 \registers_reg[789][3]  ( .D(n8176), .E(n839), .CK(clk), .Q(
        \registers[789][3] ) );
  EDFFX1 \registers_reg[789][2]  ( .D(n8131), .E(n839), .CK(clk), .Q(
        \registers[789][2] ) );
  EDFFX1 \registers_reg[789][1]  ( .D(n8075), .E(n839), .CK(clk), .Q(
        \registers[789][1] ) );
  EDFFX1 \registers_reg[789][0]  ( .D(n8014), .E(n839), .CK(clk), .Q(
        \registers[789][0] ) );
  EDFFX1 \registers_reg[785][7]  ( .D(n8398), .E(n152), .CK(clk), .Q(
        \registers[785][7] ) );
  EDFFX1 \registers_reg[785][6]  ( .D(n8340), .E(n152), .CK(clk), .Q(
        \registers[785][6] ) );
  EDFFX1 \registers_reg[785][5]  ( .D(n8282), .E(n152), .CK(clk), .Q(
        \registers[785][5] ) );
  EDFFX1 \registers_reg[785][4]  ( .D(n8224), .E(n152), .CK(clk), .Q(
        \registers[785][4] ) );
  EDFFX1 \registers_reg[785][3]  ( .D(n8177), .E(n152), .CK(clk), .Q(
        \registers[785][3] ) );
  EDFFX1 \registers_reg[785][2]  ( .D(n8129), .E(n152), .CK(clk), .Q(
        \registers[785][2] ) );
  EDFFX1 \registers_reg[785][1]  ( .D(n8073), .E(n152), .CK(clk), .Q(
        \registers[785][1] ) );
  EDFFX1 \registers_reg[785][0]  ( .D(n8015), .E(n152), .CK(clk), .Q(
        \registers[785][0] ) );
  EDFFX1 \registers_reg[781][7]  ( .D(n8399), .E(n148), .CK(clk), .Q(
        \registers[781][7] ) );
  EDFFX1 \registers_reg[781][6]  ( .D(n8341), .E(n148), .CK(clk), .Q(
        \registers[781][6] ) );
  EDFFX1 \registers_reg[781][5]  ( .D(n8283), .E(n148), .CK(clk), .Q(
        \registers[781][5] ) );
  EDFFX1 \registers_reg[781][4]  ( .D(n8225), .E(n148), .CK(clk), .Q(
        \registers[781][4] ) );
  EDFFX1 \registers_reg[781][3]  ( .D(n8178), .E(n148), .CK(clk), .Q(
        \registers[781][3] ) );
  EDFFX1 \registers_reg[781][2]  ( .D(n8127), .E(n148), .CK(clk), .Q(
        \registers[781][2] ) );
  EDFFX1 \registers_reg[781][1]  ( .D(n8071), .E(n148), .CK(clk), .Q(
        \registers[781][1] ) );
  EDFFX1 \registers_reg[781][0]  ( .D(n8010), .E(n148), .CK(clk), .Q(
        \registers[781][0] ) );
  EDFFX1 \registers_reg[777][7]  ( .D(n8400), .E(n144), .CK(clk), .Q(
        \registers[777][7] ) );
  EDFFX1 \registers_reg[777][6]  ( .D(n8342), .E(n144), .CK(clk), .Q(
        \registers[777][6] ) );
  EDFFX1 \registers_reg[777][5]  ( .D(n8284), .E(n144), .CK(clk), .Q(
        \registers[777][5] ) );
  EDFFX1 \registers_reg[777][4]  ( .D(n8226), .E(n144), .CK(clk), .Q(
        \registers[777][4] ) );
  EDFFX1 \registers_reg[777][3]  ( .D(n8176), .E(n144), .CK(clk), .Q(
        \registers[777][3] ) );
  EDFFX1 \registers_reg[777][2]  ( .D(n8128), .E(n144), .CK(clk), .Q(
        \registers[777][2] ) );
  EDFFX1 \registers_reg[777][1]  ( .D(n8072), .E(n144), .CK(clk), .Q(
        \registers[777][1] ) );
  EDFFX1 \registers_reg[777][0]  ( .D(n8011), .E(n144), .CK(clk), .Q(
        \registers[777][0] ) );
  EDFFX1 \registers_reg[773][7]  ( .D(n8396), .E(n320), .CK(clk), .Q(
        \registers[773][7] ) );
  EDFFX1 \registers_reg[773][6]  ( .D(n8338), .E(n320), .CK(clk), .Q(
        \registers[773][6] ) );
  EDFFX1 \registers_reg[773][5]  ( .D(n8280), .E(n320), .CK(clk), .Q(
        \registers[773][5] ) );
  EDFFX1 \registers_reg[773][4]  ( .D(n8222), .E(n320), .CK(clk), .Q(
        \registers[773][4] ) );
  EDFFX1 \registers_reg[773][3]  ( .D(n8177), .E(n320), .CK(clk), .Q(
        \registers[773][3] ) );
  EDFFX1 \registers_reg[773][2]  ( .D(n8126), .E(n320), .CK(clk), .Q(
        \registers[773][2] ) );
  EDFFX1 \registers_reg[773][1]  ( .D(n8070), .E(n320), .CK(clk), .Q(
        \registers[773][1] ) );
  EDFFX1 \registers_reg[773][0]  ( .D(n8012), .E(n320), .CK(clk), .Q(
        \registers[773][0] ) );
  EDFFX1 \registers_reg[769][7]  ( .D(n8397), .E(n316), .CK(clk), .Q(
        \registers[769][7] ) );
  EDFFX1 \registers_reg[769][6]  ( .D(n8339), .E(n316), .CK(clk), .Q(
        \registers[769][6] ) );
  EDFFX1 \registers_reg[769][5]  ( .D(n8281), .E(n316), .CK(clk), .Q(
        \registers[769][5] ) );
  EDFFX1 \registers_reg[769][4]  ( .D(n8223), .E(n316), .CK(clk), .Q(
        \registers[769][4] ) );
  EDFFX1 \registers_reg[769][3]  ( .D(n8178), .E(n316), .CK(clk), .Q(
        \registers[769][3] ) );
  EDFFX1 \registers_reg[769][2]  ( .D(n8127), .E(n316), .CK(clk), .Q(
        \registers[769][2] ) );
  EDFFX1 \registers_reg[769][1]  ( .D(n8071), .E(n316), .CK(clk), .Q(
        \registers[769][1] ) );
  EDFFX1 \registers_reg[769][0]  ( .D(n8010), .E(n316), .CK(clk), .Q(
        \registers[769][0] ) );
  EDFFX1 \registers_reg[765][7]  ( .D(n8383), .E(n835), .CK(clk), .Q(
        \registers[765][7] ) );
  EDFFX1 \registers_reg[765][6]  ( .D(n8325), .E(n835), .CK(clk), .Q(
        \registers[765][6] ) );
  EDFFX1 \registers_reg[765][5]  ( .D(n8267), .E(n835), .CK(clk), .Q(
        \registers[765][5] ) );
  EDFFX1 \registers_reg[765][4]  ( .D(n8209), .E(n835), .CK(clk), .Q(
        \registers[765][4] ) );
  EDFFX1 \registers_reg[765][3]  ( .D(n8164), .E(n835), .CK(clk), .Q(
        \registers[765][3] ) );
  EDFFX1 \registers_reg[765][2]  ( .D(n8113), .E(n835), .CK(clk), .Q(
        \registers[765][2] ) );
  EDFFX1 \registers_reg[765][1]  ( .D(n8057), .E(n835), .CK(clk), .Q(
        \registers[765][1] ) );
  EDFFX1 \registers_reg[765][0]  ( .D(n7997), .E(n835), .CK(clk), .Q(
        \registers[765][0] ) );
  EDFFX1 \registers_reg[761][7]  ( .D(n8381), .E(n831), .CK(clk), .Q(
        \registers[761][7] ) );
  EDFFX1 \registers_reg[761][6]  ( .D(n8323), .E(n831), .CK(clk), .Q(
        \registers[761][6] ) );
  EDFFX1 \registers_reg[761][5]  ( .D(n8265), .E(n831), .CK(clk), .Q(
        \registers[761][5] ) );
  EDFFX1 \registers_reg[761][4]  ( .D(n8207), .E(n831), .CK(clk), .Q(
        \registers[761][4] ) );
  EDFFX1 \registers_reg[761][3]  ( .D(n8165), .E(n831), .CK(clk), .Q(
        \registers[761][3] ) );
  EDFFX1 \registers_reg[761][2]  ( .D(n8111), .E(n831), .CK(clk), .Q(
        \registers[761][2] ) );
  EDFFX1 \registers_reg[761][1]  ( .D(n8055), .E(n831), .CK(clk), .Q(
        \registers[761][1] ) );
  EDFFX1 \registers_reg[761][0]  ( .D(n7994), .E(n831), .CK(clk), .Q(
        \registers[761][0] ) );
  EDFFX1 \registers_reg[757][7]  ( .D(n8382), .E(n827), .CK(clk), .Q(
        \registers[757][7] ) );
  EDFFX1 \registers_reg[757][6]  ( .D(n8324), .E(n827), .CK(clk), .Q(
        \registers[757][6] ) );
  EDFFX1 \registers_reg[757][5]  ( .D(n8266), .E(n827), .CK(clk), .Q(
        \registers[757][5] ) );
  EDFFX1 \registers_reg[757][4]  ( .D(n8208), .E(n827), .CK(clk), .Q(
        \registers[757][4] ) );
  EDFFX1 \registers_reg[757][3]  ( .D(n8166), .E(n827), .CK(clk), .Q(
        \registers[757][3] ) );
  EDFFX1 \registers_reg[757][2]  ( .D(n8112), .E(n827), .CK(clk), .Q(
        \registers[757][2] ) );
  EDFFX1 \registers_reg[757][1]  ( .D(n8056), .E(n827), .CK(clk), .Q(
        \registers[757][1] ) );
  EDFFX1 \registers_reg[757][0]  ( .D(n7996), .E(n827), .CK(clk), .Q(
        \registers[757][0] ) );
  EDFFX1 \registers_reg[753][7]  ( .D(n8383), .E(n140), .CK(clk), .Q(
        \registers[753][7] ) );
  EDFFX1 \registers_reg[753][6]  ( .D(n8325), .E(n140), .CK(clk), .Q(
        \registers[753][6] ) );
  EDFFX1 \registers_reg[753][5]  ( .D(n8267), .E(n140), .CK(clk), .Q(
        \registers[753][5] ) );
  EDFFX1 \registers_reg[753][4]  ( .D(n8209), .E(n140), .CK(clk), .Q(
        \registers[753][4] ) );
  EDFFX1 \registers_reg[753][3]  ( .D(n8758), .E(n140), .CK(clk), .Q(
        \registers[753][3] ) );
  EDFFX1 \registers_reg[753][2]  ( .D(n8113), .E(n140), .CK(clk), .Q(
        \registers[753][2] ) );
  EDFFX1 \registers_reg[753][1]  ( .D(n8057), .E(n140), .CK(clk), .Q(
        \registers[753][1] ) );
  EDFFX1 \registers_reg[753][0]  ( .D(n7997), .E(n140), .CK(clk), .Q(
        \registers[753][0] ) );
  EDFFX1 \registers_reg[749][7]  ( .D(n8381), .E(n136), .CK(clk), .Q(
        \registers[749][7] ) );
  EDFFX1 \registers_reg[749][6]  ( .D(n8323), .E(n136), .CK(clk), .Q(
        \registers[749][6] ) );
  EDFFX1 \registers_reg[749][5]  ( .D(n8265), .E(n136), .CK(clk), .Q(
        \registers[749][5] ) );
  EDFFX1 \registers_reg[749][4]  ( .D(n8207), .E(n136), .CK(clk), .Q(
        \registers[749][4] ) );
  EDFFX1 \registers_reg[749][3]  ( .D(n8162), .E(n136), .CK(clk), .Q(
        \registers[749][3] ) );
  EDFFX1 \registers_reg[749][2]  ( .D(n8111), .E(n136), .CK(clk), .Q(
        \registers[749][2] ) );
  EDFFX1 \registers_reg[749][1]  ( .D(n8055), .E(n136), .CK(clk), .Q(
        \registers[749][1] ) );
  EDFFX1 \registers_reg[749][0]  ( .D(n8680), .E(n136), .CK(clk), .Q(
        \registers[749][0] ) );
  EDFFX1 \registers_reg[745][7]  ( .D(n8382), .E(n132), .CK(clk), .Q(
        \registers[745][7] ) );
  EDFFX1 \registers_reg[745][6]  ( .D(n8324), .E(n132), .CK(clk), .Q(
        \registers[745][6] ) );
  EDFFX1 \registers_reg[745][5]  ( .D(n8266), .E(n132), .CK(clk), .Q(
        \registers[745][5] ) );
  EDFFX1 \registers_reg[745][4]  ( .D(n8208), .E(n132), .CK(clk), .Q(
        \registers[745][4] ) );
  EDFFX1 \registers_reg[745][3]  ( .D(n8163), .E(n132), .CK(clk), .Q(
        \registers[745][3] ) );
  EDFFX1 \registers_reg[745][2]  ( .D(n8112), .E(n132), .CK(clk), .Q(
        \registers[745][2] ) );
  EDFFX1 \registers_reg[745][1]  ( .D(n8056), .E(n132), .CK(clk), .Q(
        \registers[745][1] ) );
  EDFFX1 \registers_reg[745][0]  ( .D(n7996), .E(n132), .CK(clk), .Q(
        \registers[745][0] ) );
  EDFFX1 \registers_reg[741][7]  ( .D(n8383), .E(n313), .CK(clk), .Q(
        \registers[741][7] ) );
  EDFFX1 \registers_reg[741][6]  ( .D(n8325), .E(n313), .CK(clk), .Q(
        \registers[741][6] ) );
  EDFFX1 \registers_reg[741][5]  ( .D(n8267), .E(n313), .CK(clk), .Q(
        \registers[741][5] ) );
  EDFFX1 \registers_reg[741][4]  ( .D(n8209), .E(n313), .CK(clk), .Q(
        \registers[741][4] ) );
  EDFFX1 \registers_reg[741][3]  ( .D(n8754), .E(n313), .CK(clk), .Q(
        \registers[741][3] ) );
  EDFFX1 \registers_reg[741][2]  ( .D(n8113), .E(n313), .CK(clk), .Q(
        \registers[741][2] ) );
  EDFFX1 \registers_reg[741][1]  ( .D(n8057), .E(n313), .CK(clk), .Q(
        \registers[741][1] ) );
  EDFFX1 \registers_reg[741][0]  ( .D(n7997), .E(n313), .CK(clk), .Q(
        \registers[741][0] ) );
  EDFFX1 \registers_reg[737][7]  ( .D(n8381), .E(n309), .CK(clk), .Q(
        \registers[737][7] ) );
  EDFFX1 \registers_reg[737][6]  ( .D(n8323), .E(n309), .CK(clk), .Q(
        \registers[737][6] ) );
  EDFFX1 \registers_reg[737][5]  ( .D(n8265), .E(n309), .CK(clk), .Q(
        \registers[737][5] ) );
  EDFFX1 \registers_reg[737][4]  ( .D(n8207), .E(n309), .CK(clk), .Q(
        \registers[737][4] ) );
  EDFFX1 \registers_reg[737][3]  ( .D(n8162), .E(n309), .CK(clk), .Q(
        \registers[737][3] ) );
  EDFFX1 \registers_reg[737][2]  ( .D(n8111), .E(n309), .CK(clk), .Q(
        \registers[737][2] ) );
  EDFFX1 \registers_reg[737][1]  ( .D(n8055), .E(n309), .CK(clk), .Q(
        \registers[737][1] ) );
  EDFFX1 \registers_reg[737][0]  ( .D(n8677), .E(n309), .CK(clk), .Q(
        \registers[737][0] ) );
  EDFFX1 \registers_reg[733][7]  ( .D(n8382), .E(n823), .CK(clk), .Q(
        \registers[733][7] ) );
  EDFFX1 \registers_reg[733][6]  ( .D(n8324), .E(n823), .CK(clk), .Q(
        \registers[733][6] ) );
  EDFFX1 \registers_reg[733][5]  ( .D(n8266), .E(n823), .CK(clk), .Q(
        \registers[733][5] ) );
  EDFFX1 \registers_reg[733][4]  ( .D(n8208), .E(n823), .CK(clk), .Q(
        \registers[733][4] ) );
  EDFFX1 \registers_reg[733][3]  ( .D(n8163), .E(n823), .CK(clk), .Q(
        \registers[733][3] ) );
  EDFFX1 \registers_reg[733][2]  ( .D(n8112), .E(n823), .CK(clk), .Q(
        \registers[733][2] ) );
  EDFFX1 \registers_reg[733][1]  ( .D(n8056), .E(n823), .CK(clk), .Q(
        \registers[733][1] ) );
  EDFFX1 \registers_reg[733][0]  ( .D(n7996), .E(n823), .CK(clk), .Q(
        \registers[733][0] ) );
  EDFFX1 \registers_reg[729][7]  ( .D(n8378), .E(n819), .CK(clk), .Q(
        \registers[729][7] ) );
  EDFFX1 \registers_reg[729][6]  ( .D(n8320), .E(n819), .CK(clk), .Q(
        \registers[729][6] ) );
  EDFFX1 \registers_reg[729][5]  ( .D(n8262), .E(n819), .CK(clk), .Q(
        \registers[729][5] ) );
  EDFFX1 \registers_reg[729][4]  ( .D(n8204), .E(n819), .CK(clk), .Q(
        \registers[729][4] ) );
  EDFFX1 \registers_reg[729][3]  ( .D(n8756), .E(n819), .CK(clk), .Q(
        \registers[729][3] ) );
  EDFFX1 \registers_reg[729][2]  ( .D(n8110), .E(n819), .CK(clk), .Q(
        \registers[729][2] ) );
  EDFFX1 \registers_reg[729][1]  ( .D(n8054), .E(n819), .CK(clk), .Q(
        \registers[729][1] ) );
  EDFFX1 \registers_reg[729][0]  ( .D(n8675), .E(n819), .CK(clk), .Q(
        \registers[729][0] ) );
  EDFFX1 \registers_reg[725][7]  ( .D(n8379), .E(n815), .CK(clk), .Q(
        \registers[725][7] ) );
  EDFFX1 \registers_reg[725][6]  ( .D(n8321), .E(n815), .CK(clk), .Q(
        \registers[725][6] ) );
  EDFFX1 \registers_reg[725][5]  ( .D(n8263), .E(n815), .CK(clk), .Q(
        \registers[725][5] ) );
  EDFFX1 \registers_reg[725][4]  ( .D(n8205), .E(n815), .CK(clk), .Q(
        \registers[725][4] ) );
  EDFFX1 \registers_reg[725][3]  ( .D(n8162), .E(n815), .CK(clk), .Q(
        \registers[725][3] ) );
  EDFFX1 \registers_reg[725][2]  ( .D(n8108), .E(n815), .CK(clk), .Q(
        \registers[725][2] ) );
  EDFFX1 \registers_reg[725][1]  ( .D(n8052), .E(n815), .CK(clk), .Q(
        \registers[725][1] ) );
  EDFFX1 \registers_reg[725][0]  ( .D(n8028), .E(n815), .CK(clk), .Q(
        \registers[725][0] ) );
  EDFFX1 \registers_reg[721][7]  ( .D(n8380), .E(n128), .CK(clk), .Q(
        \registers[721][7] ) );
  EDFFX1 \registers_reg[721][6]  ( .D(n8322), .E(n128), .CK(clk), .Q(
        \registers[721][6] ) );
  EDFFX1 \registers_reg[721][5]  ( .D(n8264), .E(n128), .CK(clk), .Q(
        \registers[721][5] ) );
  EDFFX1 \registers_reg[721][4]  ( .D(n8206), .E(n128), .CK(clk), .Q(
        \registers[721][4] ) );
  EDFFX1 \registers_reg[721][3]  ( .D(n8163), .E(n128), .CK(clk), .Q(
        \registers[721][3] ) );
  EDFFX1 \registers_reg[721][2]  ( .D(n8109), .E(n128), .CK(clk), .Q(
        \registers[721][2] ) );
  EDFFX1 \registers_reg[721][1]  ( .D(n8053), .E(n128), .CK(clk), .Q(
        \registers[721][1] ) );
  EDFFX1 \registers_reg[721][0]  ( .D(n7995), .E(n128), .CK(clk), .Q(
        \registers[721][0] ) );
  EDFFX1 \registers_reg[717][7]  ( .D(n8378), .E(n124), .CK(clk), .Q(
        \registers[717][7] ) );
  EDFFX1 \registers_reg[717][6]  ( .D(n8320), .E(n124), .CK(clk), .Q(
        \registers[717][6] ) );
  EDFFX1 \registers_reg[717][5]  ( .D(n8262), .E(n124), .CK(clk), .Q(
        \registers[717][5] ) );
  EDFFX1 \registers_reg[717][4]  ( .D(n8204), .E(n124), .CK(clk), .Q(
        \registers[717][4] ) );
  EDFFX1 \registers_reg[717][3]  ( .D(n8755), .E(n124), .CK(clk), .Q(
        \registers[717][3] ) );
  EDFFX1 \registers_reg[717][2]  ( .D(n8110), .E(n124), .CK(clk), .Q(
        \registers[717][2] ) );
  EDFFX1 \registers_reg[717][1]  ( .D(n8054), .E(n124), .CK(clk), .Q(
        \registers[717][1] ) );
  EDFFX1 \registers_reg[717][0]  ( .D(n8671), .E(n124), .CK(clk), .Q(
        \registers[717][0] ) );
  EDFFX1 \registers_reg[713][7]  ( .D(n8379), .E(n120), .CK(clk), .Q(
        \registers[713][7] ) );
  EDFFX1 \registers_reg[713][6]  ( .D(n8321), .E(n120), .CK(clk), .Q(
        \registers[713][6] ) );
  EDFFX1 \registers_reg[713][5]  ( .D(n8263), .E(n120), .CK(clk), .Q(
        \registers[713][5] ) );
  EDFFX1 \registers_reg[713][4]  ( .D(n8205), .E(n120), .CK(clk), .Q(
        \registers[713][4] ) );
  EDFFX1 \registers_reg[713][3]  ( .D(n8162), .E(n120), .CK(clk), .Q(
        \registers[713][3] ) );
  EDFFX1 \registers_reg[713][2]  ( .D(n8108), .E(n120), .CK(clk), .Q(
        \registers[713][2] ) );
  EDFFX1 \registers_reg[713][1]  ( .D(n8052), .E(n120), .CK(clk), .Q(
        \registers[713][1] ) );
  EDFFX1 \registers_reg[713][0]  ( .D(n8030), .E(n120), .CK(clk), .Q(
        \registers[713][0] ) );
  EDFFX1 \registers_reg[709][7]  ( .D(n8380), .E(n306), .CK(clk), .Q(
        \registers[709][7] ) );
  EDFFX1 \registers_reg[709][6]  ( .D(n8322), .E(n306), .CK(clk), .Q(
        \registers[709][6] ) );
  EDFFX1 \registers_reg[709][5]  ( .D(n8264), .E(n306), .CK(clk), .Q(
        \registers[709][5] ) );
  EDFFX1 \registers_reg[709][4]  ( .D(n8206), .E(n306), .CK(clk), .Q(
        \registers[709][4] ) );
  EDFFX1 \registers_reg[709][3]  ( .D(n8163), .E(n306), .CK(clk), .Q(
        \registers[709][3] ) );
  EDFFX1 \registers_reg[709][2]  ( .D(n8109), .E(n306), .CK(clk), .Q(
        \registers[709][2] ) );
  EDFFX1 \registers_reg[709][1]  ( .D(n8053), .E(n306), .CK(clk), .Q(
        \registers[709][1] ) );
  EDFFX1 \registers_reg[709][0]  ( .D(n7995), .E(n306), .CK(clk), .Q(
        \registers[709][0] ) );
  EDFFX1 \registers_reg[705][7]  ( .D(n8378), .E(n302), .CK(clk), .Q(
        \registers[705][7] ) );
  EDFFX1 \registers_reg[705][6]  ( .D(n8320), .E(n302), .CK(clk), .Q(
        \registers[705][6] ) );
  EDFFX1 \registers_reg[705][5]  ( .D(n8262), .E(n302), .CK(clk), .Q(
        \registers[705][5] ) );
  EDFFX1 \registers_reg[705][4]  ( .D(n8204), .E(n302), .CK(clk), .Q(
        \registers[705][4] ) );
  EDFFX1 \registers_reg[705][3]  ( .D(n8761), .E(n302), .CK(clk), .Q(
        \registers[705][3] ) );
  EDFFX1 \registers_reg[705][2]  ( .D(n8110), .E(n302), .CK(clk), .Q(
        \registers[705][2] ) );
  EDFFX1 \registers_reg[705][1]  ( .D(n8054), .E(n302), .CK(clk), .Q(
        \registers[705][1] ) );
  EDFFX1 \registers_reg[705][0]  ( .D(n8670), .E(n302), .CK(clk), .Q(
        \registers[705][0] ) );
  EDFFX1 \registers_reg[701][7]  ( .D(n8380), .E(n811), .CK(clk), .Q(
        \registers[701][7] ) );
  EDFFX1 \registers_reg[701][6]  ( .D(n8322), .E(n811), .CK(clk), .Q(
        \registers[701][6] ) );
  EDFFX1 \registers_reg[701][5]  ( .D(n8264), .E(n811), .CK(clk), .Q(
        \registers[701][5] ) );
  EDFFX1 \registers_reg[701][4]  ( .D(n8206), .E(n811), .CK(clk), .Q(
        \registers[701][4] ) );
  EDFFX1 \registers_reg[701][3]  ( .D(n8163), .E(n811), .CK(clk), .Q(
        \registers[701][3] ) );
  EDFFX1 \registers_reg[701][2]  ( .D(n8109), .E(n811), .CK(clk), .Q(
        \registers[701][2] ) );
  EDFFX1 \registers_reg[701][1]  ( .D(n8053), .E(n811), .CK(clk), .Q(
        \registers[701][1] ) );
  EDFFX1 \registers_reg[701][0]  ( .D(n7995), .E(n811), .CK(clk), .Q(
        \registers[701][0] ) );
  EDFFX1 \registers_reg[697][7]  ( .D(n8378), .E(n807), .CK(clk), .Q(
        \registers[697][7] ) );
  EDFFX1 \registers_reg[697][6]  ( .D(n8320), .E(n807), .CK(clk), .Q(
        \registers[697][6] ) );
  EDFFX1 \registers_reg[697][5]  ( .D(n8262), .E(n807), .CK(clk), .Q(
        \registers[697][5] ) );
  EDFFX1 \registers_reg[697][4]  ( .D(n8204), .E(n807), .CK(clk), .Q(
        \registers[697][4] ) );
  EDFFX1 \registers_reg[697][3]  ( .D(n8760), .E(n807), .CK(clk), .Q(
        \registers[697][3] ) );
  EDFFX1 \registers_reg[697][2]  ( .D(n8110), .E(n807), .CK(clk), .Q(
        \registers[697][2] ) );
  EDFFX1 \registers_reg[697][1]  ( .D(n8054), .E(n807), .CK(clk), .Q(
        \registers[697][1] ) );
  EDFFX1 \registers_reg[697][0]  ( .D(n8673), .E(n807), .CK(clk), .Q(
        \registers[697][0] ) );
  EDFFX1 \registers_reg[693][7]  ( .D(n8379), .E(n803), .CK(clk), .Q(
        \registers[693][7] ) );
  EDFFX1 \registers_reg[693][6]  ( .D(n8321), .E(n803), .CK(clk), .Q(
        \registers[693][6] ) );
  EDFFX1 \registers_reg[693][5]  ( .D(n8263), .E(n803), .CK(clk), .Q(
        \registers[693][5] ) );
  EDFFX1 \registers_reg[693][4]  ( .D(n8205), .E(n803), .CK(clk), .Q(
        \registers[693][4] ) );
  EDFFX1 \registers_reg[693][3]  ( .D(n8162), .E(n803), .CK(clk), .Q(
        \registers[693][3] ) );
  EDFFX1 \registers_reg[693][2]  ( .D(n8108), .E(n803), .CK(clk), .Q(
        \registers[693][2] ) );
  EDFFX1 \registers_reg[693][1]  ( .D(n8052), .E(n803), .CK(clk), .Q(
        \registers[693][1] ) );
  EDFFX1 \registers_reg[693][0]  ( .D(n8029), .E(n803), .CK(clk), .Q(
        \registers[693][0] ) );
  EDFFX1 \registers_reg[689][7]  ( .D(n8380), .E(n116), .CK(clk), .Q(
        \registers[689][7] ) );
  EDFFX1 \registers_reg[689][6]  ( .D(n8322), .E(n116), .CK(clk), .Q(
        \registers[689][6] ) );
  EDFFX1 \registers_reg[689][5]  ( .D(n8264), .E(n116), .CK(clk), .Q(
        \registers[689][5] ) );
  EDFFX1 \registers_reg[689][4]  ( .D(n8206), .E(n116), .CK(clk), .Q(
        \registers[689][4] ) );
  EDFFX1 \registers_reg[689][3]  ( .D(n8161), .E(n116), .CK(clk), .Q(
        \registers[689][3] ) );
  EDFFX1 \registers_reg[689][2]  ( .D(n8109), .E(n116), .CK(clk), .Q(
        \registers[689][2] ) );
  EDFFX1 \registers_reg[689][1]  ( .D(n8053), .E(n116), .CK(clk), .Q(
        \registers[689][1] ) );
  EDFFX1 \registers_reg[689][0]  ( .D(n7995), .E(n116), .CK(clk), .Q(
        \registers[689][0] ) );
  EDFFX1 \registers_reg[685][7]  ( .D(n8378), .E(n112), .CK(clk), .Q(
        \registers[685][7] ) );
  EDFFX1 \registers_reg[685][6]  ( .D(n8320), .E(n112), .CK(clk), .Q(
        \registers[685][6] ) );
  EDFFX1 \registers_reg[685][5]  ( .D(n8262), .E(n112), .CK(clk), .Q(
        \registers[685][5] ) );
  EDFFX1 \registers_reg[685][4]  ( .D(n8204), .E(n112), .CK(clk), .Q(
        \registers[685][4] ) );
  EDFFX1 \registers_reg[685][3]  ( .D(n8161), .E(n112), .CK(clk), .Q(
        \registers[685][3] ) );
  EDFFX1 \registers_reg[685][2]  ( .D(n8110), .E(n112), .CK(clk), .Q(
        \registers[685][2] ) );
  EDFFX1 \registers_reg[685][1]  ( .D(n8054), .E(n112), .CK(clk), .Q(
        \registers[685][1] ) );
  EDFFX1 \registers_reg[685][0]  ( .D(n8672), .E(n112), .CK(clk), .Q(
        \registers[685][0] ) );
  EDFFX1 \registers_reg[681][7]  ( .D(n8379), .E(n108), .CK(clk), .Q(
        \registers[681][7] ) );
  EDFFX1 \registers_reg[681][6]  ( .D(n8321), .E(n108), .CK(clk), .Q(
        \registers[681][6] ) );
  EDFFX1 \registers_reg[681][5]  ( .D(n8263), .E(n108), .CK(clk), .Q(
        \registers[681][5] ) );
  EDFFX1 \registers_reg[681][4]  ( .D(n8205), .E(n108), .CK(clk), .Q(
        \registers[681][4] ) );
  EDFFX1 \registers_reg[681][3]  ( .D(n8161), .E(n108), .CK(clk), .Q(
        \registers[681][3] ) );
  EDFFX1 \registers_reg[681][2]  ( .D(n8105), .E(n108), .CK(clk), .Q(
        \registers[681][2] ) );
  EDFFX1 \registers_reg[681][1]  ( .D(n8049), .E(n108), .CK(clk), .Q(
        \registers[681][1] ) );
  EDFFX1 \registers_reg[681][0]  ( .D(n8687), .E(n108), .CK(clk), .Q(
        \registers[681][0] ) );
  EDFFX1 \registers_reg[677][7]  ( .D(n8377), .E(n299), .CK(clk), .Q(
        \registers[677][7] ) );
  EDFFX1 \registers_reg[677][6]  ( .D(n8319), .E(n299), .CK(clk), .Q(
        \registers[677][6] ) );
  EDFFX1 \registers_reg[677][5]  ( .D(n8261), .E(n299), .CK(clk), .Q(
        \registers[677][5] ) );
  EDFFX1 \registers_reg[677][4]  ( .D(n8203), .E(n299), .CK(clk), .Q(
        \registers[677][4] ) );
  EDFFX1 \registers_reg[677][3]  ( .D(n8161), .E(n299), .CK(clk), .Q(
        \registers[677][3] ) );
  EDFFX1 \registers_reg[677][2]  ( .D(n8106), .E(n299), .CK(clk), .Q(
        \registers[677][2] ) );
  EDFFX1 \registers_reg[677][1]  ( .D(n8050), .E(n299), .CK(clk), .Q(
        \registers[677][1] ) );
  EDFFX1 \registers_reg[677][0]  ( .D(n7994), .E(n299), .CK(clk), .Q(
        \registers[677][0] ) );
  EDFFX1 \registers_reg[673][7]  ( .D(n8377), .E(n295), .CK(clk), .Q(
        \registers[673][7] ) );
  EDFFX1 \registers_reg[673][6]  ( .D(n8319), .E(n295), .CK(clk), .Q(
        \registers[673][6] ) );
  EDFFX1 \registers_reg[673][5]  ( .D(n8261), .E(n295), .CK(clk), .Q(
        \registers[673][5] ) );
  EDFFX1 \registers_reg[673][4]  ( .D(n8203), .E(n295), .CK(clk), .Q(
        \registers[673][4] ) );
  EDFFX1 \registers_reg[673][3]  ( .D(n8175), .E(n295), .CK(clk), .Q(
        \registers[673][3] ) );
  EDFFX1 \registers_reg[673][2]  ( .D(n8107), .E(n295), .CK(clk), .Q(
        \registers[673][2] ) );
  EDFFX1 \registers_reg[673][1]  ( .D(n8051), .E(n295), .CK(clk), .Q(
        \registers[673][1] ) );
  EDFFX1 \registers_reg[673][0]  ( .D(n7994), .E(n295), .CK(clk), .Q(
        \registers[673][0] ) );
  EDFFX1 \registers_reg[669][7]  ( .D(n8394), .E(n799), .CK(clk), .Q(
        \registers[669][7] ) );
  EDFFX1 \registers_reg[669][6]  ( .D(n8336), .E(n799), .CK(clk), .Q(
        \registers[669][6] ) );
  EDFFX1 \registers_reg[669][5]  ( .D(n8278), .E(n799), .CK(clk), .Q(
        \registers[669][5] ) );
  EDFFX1 \registers_reg[669][4]  ( .D(n8220), .E(n799), .CK(clk), .Q(
        \registers[669][4] ) );
  EDFFX1 \registers_reg[669][3]  ( .D(n8179), .E(n799), .CK(clk), .Q(
        \registers[669][3] ) );
  EDFFX1 \registers_reg[669][2]  ( .D(n8105), .E(n799), .CK(clk), .Q(
        \registers[669][2] ) );
  EDFFX1 \registers_reg[669][1]  ( .D(n8049), .E(n799), .CK(clk), .Q(
        \registers[669][1] ) );
  EDFFX1 \registers_reg[669][0]  ( .D(n7994), .E(n799), .CK(clk), .Q(
        \registers[669][0] ) );
  EDFFX1 \registers_reg[665][7]  ( .D(n8391), .E(n795), .CK(clk), .Q(
        \registers[665][7] ) );
  EDFFX1 \registers_reg[665][6]  ( .D(n8333), .E(n795), .CK(clk), .Q(
        \registers[665][6] ) );
  EDFFX1 \registers_reg[665][5]  ( .D(n8275), .E(n795), .CK(clk), .Q(
        \registers[665][5] ) );
  EDFFX1 \registers_reg[665][4]  ( .D(n8217), .E(n795), .CK(clk), .Q(
        \registers[665][4] ) );
  EDFFX1 \registers_reg[665][3]  ( .D(n8180), .E(n795), .CK(clk), .Q(
        \registers[665][3] ) );
  EDFFX1 \registers_reg[665][2]  ( .D(n8106), .E(n795), .CK(clk), .Q(
        \registers[665][2] ) );
  EDFFX1 \registers_reg[665][1]  ( .D(n8050), .E(n795), .CK(clk), .Q(
        \registers[665][1] ) );
  EDFFX1 \registers_reg[665][0]  ( .D(n8668), .E(n795), .CK(clk), .Q(
        \registers[665][0] ) );
  EDFFX1 \registers_reg[661][7]  ( .D(n8388), .E(n791), .CK(clk), .Q(
        \registers[661][7] ) );
  EDFFX1 \registers_reg[661][6]  ( .D(n8330), .E(n791), .CK(clk), .Q(
        \registers[661][6] ) );
  EDFFX1 \registers_reg[661][5]  ( .D(n8272), .E(n791), .CK(clk), .Q(
        \registers[661][5] ) );
  EDFFX1 \registers_reg[661][4]  ( .D(n8214), .E(n791), .CK(clk), .Q(
        \registers[661][4] ) );
  EDFFX1 \registers_reg[661][3]  ( .D(n8181), .E(n791), .CK(clk), .Q(
        \registers[661][3] ) );
  EDFFX1 \registers_reg[661][2]  ( .D(n8107), .E(n791), .CK(clk), .Q(
        \registers[661][2] ) );
  EDFFX1 \registers_reg[661][1]  ( .D(n8051), .E(n791), .CK(clk), .Q(
        \registers[661][1] ) );
  EDFFX1 \registers_reg[661][0]  ( .D(n8669), .E(n791), .CK(clk), .Q(
        \registers[661][0] ) );
  EDFFX1 \registers_reg[657][7]  ( .D(n8385), .E(n104), .CK(clk), .Q(
        \registers[657][7] ) );
  EDFFX1 \registers_reg[657][6]  ( .D(n8327), .E(n104), .CK(clk), .Q(
        \registers[657][6] ) );
  EDFFX1 \registers_reg[657][5]  ( .D(n8269), .E(n104), .CK(clk), .Q(
        \registers[657][5] ) );
  EDFFX1 \registers_reg[657][4]  ( .D(n8211), .E(n104), .CK(clk), .Q(
        \registers[657][4] ) );
  EDFFX1 \registers_reg[657][3]  ( .D(n8177), .E(n104), .CK(clk), .Q(
        \registers[657][3] ) );
  EDFFX1 \registers_reg[657][2]  ( .D(n8105), .E(n104), .CK(clk), .Q(
        \registers[657][2] ) );
  EDFFX1 \registers_reg[657][1]  ( .D(n8049), .E(n104), .CK(clk), .Q(
        \registers[657][1] ) );
  EDFFX1 \registers_reg[657][0]  ( .D(n8667), .E(n104), .CK(clk), .Q(
        \registers[657][0] ) );
  EDFFX1 \registers_reg[653][7]  ( .D(n8383), .E(n100), .CK(clk), .Q(
        \registers[653][7] ) );
  EDFFX1 \registers_reg[653][6]  ( .D(n8325), .E(n100), .CK(clk), .Q(
        \registers[653][6] ) );
  EDFFX1 \registers_reg[653][5]  ( .D(n8267), .E(n100), .CK(clk), .Q(
        \registers[653][5] ) );
  EDFFX1 \registers_reg[653][4]  ( .D(n8209), .E(n100), .CK(clk), .Q(
        \registers[653][4] ) );
  EDFFX1 \registers_reg[653][3]  ( .D(n8178), .E(n100), .CK(clk), .Q(
        \registers[653][3] ) );
  EDFFX1 \registers_reg[653][2]  ( .D(n8106), .E(n100), .CK(clk), .Q(
        \registers[653][2] ) );
  EDFFX1 \registers_reg[653][1]  ( .D(n8050), .E(n100), .CK(clk), .Q(
        \registers[653][1] ) );
  EDFFX1 \registers_reg[653][0]  ( .D(n8666), .E(n100), .CK(clk), .Q(
        \registers[653][0] ) );
  EDFFX1 \registers_reg[649][7]  ( .D(n8380), .E(n96), .CK(clk), .Q(
        \registers[649][7] ) );
  EDFFX1 \registers_reg[649][6]  ( .D(n8322), .E(n96), .CK(clk), .Q(
        \registers[649][6] ) );
  EDFFX1 \registers_reg[649][5]  ( .D(n8264), .E(n96), .CK(clk), .Q(
        \registers[649][5] ) );
  EDFFX1 \registers_reg[649][4]  ( .D(n8206), .E(n96), .CK(clk), .Q(
        \registers[649][4] ) );
  EDFFX1 \registers_reg[649][3]  ( .D(n8176), .E(n96), .CK(clk), .Q(
        \registers[649][3] ) );
  EDFFX1 \registers_reg[649][2]  ( .D(n8107), .E(n96), .CK(clk), .Q(
        \registers[649][2] ) );
  EDFFX1 \registers_reg[649][1]  ( .D(n8051), .E(n96), .CK(clk), .Q(
        \registers[649][1] ) );
  EDFFX1 \registers_reg[649][0]  ( .D(n8048), .E(n96), .CK(clk), .Q(
        \registers[649][0] ) );
  EDFFX1 \registers_reg[645][7]  ( .D(n8397), .E(n292), .CK(clk), .Q(
        \registers[645][7] ) );
  EDFFX1 \registers_reg[645][6]  ( .D(n8339), .E(n292), .CK(clk), .Q(
        \registers[645][6] ) );
  EDFFX1 \registers_reg[645][5]  ( .D(n8281), .E(n292), .CK(clk), .Q(
        \registers[645][5] ) );
  EDFFX1 \registers_reg[645][4]  ( .D(n8223), .E(n292), .CK(clk), .Q(
        \registers[645][4] ) );
  EDFFX1 \registers_reg[645][3]  ( .D(n8763), .E(n292), .CK(clk), .Q(
        \registers[645][3] ) );
  EDFFX1 \registers_reg[645][2]  ( .D(n8105), .E(n292), .CK(clk), .Q(
        \registers[645][2] ) );
  EDFFX1 \registers_reg[645][1]  ( .D(n8049), .E(n292), .CK(clk), .Q(
        \registers[645][1] ) );
  EDFFX1 \registers_reg[645][0]  ( .D(n8032), .E(n292), .CK(clk), .Q(
        \registers[645][0] ) );
  EDFFX1 \registers_reg[641][7]  ( .D(n8400), .E(n288), .CK(clk), .Q(
        \registers[641][7] ) );
  EDFFX1 \registers_reg[641][6]  ( .D(n8342), .E(n288), .CK(clk), .Q(
        \registers[641][6] ) );
  EDFFX1 \registers_reg[641][5]  ( .D(n8284), .E(n288), .CK(clk), .Q(
        \registers[641][5] ) );
  EDFFX1 \registers_reg[641][4]  ( .D(n8226), .E(n288), .CK(clk), .Q(
        \registers[641][4] ) );
  EDFFX1 \registers_reg[641][3]  ( .D(n8762), .E(n288), .CK(clk), .Q(
        \registers[641][3] ) );
  EDFFX1 \registers_reg[641][2]  ( .D(n8106), .E(n288), .CK(clk), .Q(
        \registers[641][2] ) );
  EDFFX1 \registers_reg[641][1]  ( .D(n8050), .E(n288), .CK(clk), .Q(
        \registers[641][1] ) );
  EDFFX1 \registers_reg[641][0]  ( .D(n8012), .E(n288), .CK(clk), .Q(
        \registers[641][0] ) );
  EDFFX1 \registers_reg[637][7]  ( .D(n8391), .E(n787), .CK(clk), .Q(
        \registers[637][7] ) );
  EDFFX1 \registers_reg[637][6]  ( .D(n8333), .E(n787), .CK(clk), .Q(
        \registers[637][6] ) );
  EDFFX1 \registers_reg[637][5]  ( .D(n8275), .E(n787), .CK(clk), .Q(
        \registers[637][5] ) );
  EDFFX1 \registers_reg[637][4]  ( .D(n8217), .E(n787), .CK(clk), .Q(
        \registers[637][4] ) );
  EDFFX1 \registers_reg[637][3]  ( .D(n8170), .E(n787), .CK(clk), .Q(
        \registers[637][3] ) );
  EDFFX1 \registers_reg[637][2]  ( .D(n8122), .E(n787), .CK(clk), .Q(
        \registers[637][2] ) );
  EDFFX1 \registers_reg[637][1]  ( .D(n8066), .E(n787), .CK(clk), .Q(
        \registers[637][1] ) );
  EDFFX1 \registers_reg[637][0]  ( .D(n8004), .E(n787), .CK(clk), .Q(
        \registers[637][0] ) );
  EDFFX1 \registers_reg[633][7]  ( .D(n8389), .E(n783), .CK(clk), .Q(
        \registers[633][7] ) );
  EDFFX1 \registers_reg[633][6]  ( .D(n8331), .E(n783), .CK(clk), .Q(
        \registers[633][6] ) );
  EDFFX1 \registers_reg[633][5]  ( .D(n8273), .E(n783), .CK(clk), .Q(
        \registers[633][5] ) );
  EDFFX1 \registers_reg[633][4]  ( .D(n8215), .E(n783), .CK(clk), .Q(
        \registers[633][4] ) );
  EDFFX1 \registers_reg[633][3]  ( .D(n8171), .E(n783), .CK(clk), .Q(
        \registers[633][3] ) );
  EDFFX1 \registers_reg[633][2]  ( .D(n8120), .E(n783), .CK(clk), .Q(
        \registers[633][2] ) );
  EDFFX1 \registers_reg[633][1]  ( .D(n8064), .E(n783), .CK(clk), .Q(
        \registers[633][1] ) );
  EDFFX1 \registers_reg[633][0]  ( .D(n8005), .E(n783), .CK(clk), .Q(
        \registers[633][0] ) );
  EDFFX1 \registers_reg[629][7]  ( .D(n8390), .E(n779), .CK(clk), .Q(
        \registers[629][7] ) );
  EDFFX1 \registers_reg[629][6]  ( .D(n8332), .E(n779), .CK(clk), .Q(
        \registers[629][6] ) );
  EDFFX1 \registers_reg[629][5]  ( .D(n8274), .E(n779), .CK(clk), .Q(
        \registers[629][5] ) );
  EDFFX1 \registers_reg[629][4]  ( .D(n8216), .E(n779), .CK(clk), .Q(
        \registers[629][4] ) );
  EDFFX1 \registers_reg[629][3]  ( .D(n8172), .E(n779), .CK(clk), .Q(
        \registers[629][3] ) );
  EDFFX1 \registers_reg[629][2]  ( .D(n8118), .E(n779), .CK(clk), .Q(
        \registers[629][2] ) );
  EDFFX1 \registers_reg[629][1]  ( .D(n8062), .E(n779), .CK(clk), .Q(
        \registers[629][1] ) );
  EDFFX1 \registers_reg[629][0]  ( .D(n8006), .E(n779), .CK(clk), .Q(
        \registers[629][0] ) );
  EDFFX1 \registers_reg[625][7]  ( .D(n8386), .E(n92), .CK(clk), .Q(
        \registers[625][7] ) );
  EDFFX1 \registers_reg[625][6]  ( .D(n8328), .E(n92), .CK(clk), .Q(
        \registers[625][6] ) );
  EDFFX1 \registers_reg[625][5]  ( .D(n8270), .E(n92), .CK(clk), .Q(
        \registers[625][5] ) );
  EDFFX1 \registers_reg[625][4]  ( .D(n8212), .E(n92), .CK(clk), .Q(
        \registers[625][4] ) );
  EDFFX1 \registers_reg[625][3]  ( .D(n8167), .E(n92), .CK(clk), .Q(
        \registers[625][3] ) );
  EDFFX1 \registers_reg[625][2]  ( .D(n8119), .E(n92), .CK(clk), .Q(
        \registers[625][2] ) );
  EDFFX1 \registers_reg[625][1]  ( .D(n8063), .E(n92), .CK(clk), .Q(
        \registers[625][1] ) );
  EDFFX1 \registers_reg[625][0]  ( .D(n8001), .E(n92), .CK(clk), .Q(
        \registers[625][0] ) );
  EDFFX1 \registers_reg[621][7]  ( .D(n8387), .E(n88), .CK(clk), .Q(
        \registers[621][7] ) );
  EDFFX1 \registers_reg[621][6]  ( .D(n8329), .E(n88), .CK(clk), .Q(
        \registers[621][6] ) );
  EDFFX1 \registers_reg[621][5]  ( .D(n8271), .E(n88), .CK(clk), .Q(
        \registers[621][5] ) );
  EDFFX1 \registers_reg[621][4]  ( .D(n8213), .E(n88), .CK(clk), .Q(
        \registers[621][4] ) );
  EDFFX1 \registers_reg[621][3]  ( .D(n8168), .E(n88), .CK(clk), .Q(
        \registers[621][3] ) );
  EDFFX1 \registers_reg[621][2]  ( .D(n8117), .E(n88), .CK(clk), .Q(
        \registers[621][2] ) );
  EDFFX1 \registers_reg[621][1]  ( .D(n8061), .E(n88), .CK(clk), .Q(
        \registers[621][1] ) );
  EDFFX1 \registers_reg[621][0]  ( .D(n8002), .E(n88), .CK(clk), .Q(
        \registers[621][0] ) );
  EDFFX1 \registers_reg[617][7]  ( .D(n8388), .E(n84), .CK(clk), .Q(
        \registers[617][7] ) );
  EDFFX1 \registers_reg[617][6]  ( .D(n8330), .E(n84), .CK(clk), .Q(
        \registers[617][6] ) );
  EDFFX1 \registers_reg[617][5]  ( .D(n8272), .E(n84), .CK(clk), .Q(
        \registers[617][5] ) );
  EDFFX1 \registers_reg[617][4]  ( .D(n8214), .E(n84), .CK(clk), .Q(
        \registers[617][4] ) );
  EDFFX1 \registers_reg[617][3]  ( .D(n8169), .E(n84), .CK(clk), .Q(
        \registers[617][3] ) );
  EDFFX1 \registers_reg[617][2]  ( .D(n8118), .E(n84), .CK(clk), .Q(
        \registers[617][2] ) );
  EDFFX1 \registers_reg[617][1]  ( .D(n8062), .E(n84), .CK(clk), .Q(
        \registers[617][1] ) );
  EDFFX1 \registers_reg[617][0]  ( .D(n8003), .E(n84), .CK(clk), .Q(
        \registers[617][0] ) );
  EDFFX1 \registers_reg[613][7]  ( .D(n8386), .E(n285), .CK(clk), .Q(
        \registers[613][7] ) );
  EDFFX1 \registers_reg[613][6]  ( .D(n8328), .E(n285), .CK(clk), .Q(
        \registers[613][6] ) );
  EDFFX1 \registers_reg[613][5]  ( .D(n8270), .E(n285), .CK(clk), .Q(
        \registers[613][5] ) );
  EDFFX1 \registers_reg[613][4]  ( .D(n8212), .E(n285), .CK(clk), .Q(
        \registers[613][4] ) );
  EDFFX1 \registers_reg[613][3]  ( .D(n8167), .E(n285), .CK(clk), .Q(
        \registers[613][3] ) );
  EDFFX1 \registers_reg[613][2]  ( .D(n8119), .E(n285), .CK(clk), .Q(
        \registers[613][2] ) );
  EDFFX1 \registers_reg[613][1]  ( .D(n8063), .E(n285), .CK(clk), .Q(
        \registers[613][1] ) );
  EDFFX1 \registers_reg[613][0]  ( .D(n8001), .E(n285), .CK(clk), .Q(
        \registers[613][0] ) );
  EDFFX1 \registers_reg[609][7]  ( .D(n8387), .E(n281), .CK(clk), .Q(
        \registers[609][7] ) );
  EDFFX1 \registers_reg[609][6]  ( .D(n8329), .E(n281), .CK(clk), .Q(
        \registers[609][6] ) );
  EDFFX1 \registers_reg[609][5]  ( .D(n8271), .E(n281), .CK(clk), .Q(
        \registers[609][5] ) );
  EDFFX1 \registers_reg[609][4]  ( .D(n8213), .E(n281), .CK(clk), .Q(
        \registers[609][4] ) );
  EDFFX1 \registers_reg[609][3]  ( .D(n8168), .E(n281), .CK(clk), .Q(
        \registers[609][3] ) );
  EDFFX1 \registers_reg[609][2]  ( .D(n8117), .E(n281), .CK(clk), .Q(
        \registers[609][2] ) );
  EDFFX1 \registers_reg[609][1]  ( .D(n8061), .E(n281), .CK(clk), .Q(
        \registers[609][1] ) );
  EDFFX1 \registers_reg[609][0]  ( .D(n8002), .E(n281), .CK(clk), .Q(
        \registers[609][0] ) );
  EDFFX1 \registers_reg[605][7]  ( .D(n8388), .E(n775), .CK(clk), .Q(
        \registers[605][7] ) );
  EDFFX1 \registers_reg[605][6]  ( .D(n8330), .E(n775), .CK(clk), .Q(
        \registers[605][6] ) );
  EDFFX1 \registers_reg[605][5]  ( .D(n8272), .E(n775), .CK(clk), .Q(
        \registers[605][5] ) );
  EDFFX1 \registers_reg[605][4]  ( .D(n8214), .E(n775), .CK(clk), .Q(
        \registers[605][4] ) );
  EDFFX1 \registers_reg[605][3]  ( .D(n8169), .E(n775), .CK(clk), .Q(
        \registers[605][3] ) );
  EDFFX1 \registers_reg[605][2]  ( .D(n8118), .E(n775), .CK(clk), .Q(
        \registers[605][2] ) );
  EDFFX1 \registers_reg[605][1]  ( .D(n8062), .E(n775), .CK(clk), .Q(
        \registers[605][1] ) );
  EDFFX1 \registers_reg[605][0]  ( .D(n8003), .E(n775), .CK(clk), .Q(
        \registers[605][0] ) );
  EDFFX1 \registers_reg[601][7]  ( .D(n8386), .E(n771), .CK(clk), .Q(
        \registers[601][7] ) );
  EDFFX1 \registers_reg[601][6]  ( .D(n8328), .E(n771), .CK(clk), .Q(
        \registers[601][6] ) );
  EDFFX1 \registers_reg[601][5]  ( .D(n8270), .E(n771), .CK(clk), .Q(
        \registers[601][5] ) );
  EDFFX1 \registers_reg[601][4]  ( .D(n8212), .E(n771), .CK(clk), .Q(
        \registers[601][4] ) );
  EDFFX1 \registers_reg[601][3]  ( .D(n8167), .E(n771), .CK(clk), .Q(
        \registers[601][3] ) );
  EDFFX1 \registers_reg[601][2]  ( .D(n8119), .E(n771), .CK(clk), .Q(
        \registers[601][2] ) );
  EDFFX1 \registers_reg[601][1]  ( .D(n8063), .E(n771), .CK(clk), .Q(
        \registers[601][1] ) );
  EDFFX1 \registers_reg[601][0]  ( .D(n8001), .E(n771), .CK(clk), .Q(
        \registers[601][0] ) );
  EDFFX1 \registers_reg[597][7]  ( .D(n8387), .E(n767), .CK(clk), .Q(
        \registers[597][7] ) );
  EDFFX1 \registers_reg[597][6]  ( .D(n8329), .E(n767), .CK(clk), .Q(
        \registers[597][6] ) );
  EDFFX1 \registers_reg[597][5]  ( .D(n8271), .E(n767), .CK(clk), .Q(
        \registers[597][5] ) );
  EDFFX1 \registers_reg[597][4]  ( .D(n8213), .E(n767), .CK(clk), .Q(
        \registers[597][4] ) );
  EDFFX1 \registers_reg[597][3]  ( .D(n8168), .E(n767), .CK(clk), .Q(
        \registers[597][3] ) );
  EDFFX1 \registers_reg[597][2]  ( .D(n8117), .E(n767), .CK(clk), .Q(
        \registers[597][2] ) );
  EDFFX1 \registers_reg[597][1]  ( .D(n8061), .E(n767), .CK(clk), .Q(
        \registers[597][1] ) );
  EDFFX1 \registers_reg[597][0]  ( .D(n8002), .E(n767), .CK(clk), .Q(
        \registers[597][0] ) );
  EDFFX1 \registers_reg[593][7]  ( .D(n8388), .E(n80), .CK(clk), .Q(
        \registers[593][7] ) );
  EDFFX1 \registers_reg[593][6]  ( .D(n8330), .E(n80), .CK(clk), .Q(
        \registers[593][6] ) );
  EDFFX1 \registers_reg[593][5]  ( .D(n8272), .E(n80), .CK(clk), .Q(
        \registers[593][5] ) );
  EDFFX1 \registers_reg[593][4]  ( .D(n8214), .E(n80), .CK(clk), .Q(
        \registers[593][4] ) );
  EDFFX1 \registers_reg[593][3]  ( .D(n8169), .E(n80), .CK(clk), .Q(
        \registers[593][3] ) );
  EDFFX1 \registers_reg[593][2]  ( .D(n8118), .E(n80), .CK(clk), .Q(
        \registers[593][2] ) );
  EDFFX1 \registers_reg[593][1]  ( .D(n8062), .E(n80), .CK(clk), .Q(
        \registers[593][1] ) );
  EDFFX1 \registers_reg[593][0]  ( .D(n8003), .E(n80), .CK(clk), .Q(
        \registers[593][0] ) );
  EDFFX1 \registers_reg[589][7]  ( .D(n8386), .E(n76), .CK(clk), .Q(
        \registers[589][7] ) );
  EDFFX1 \registers_reg[589][6]  ( .D(n8328), .E(n76), .CK(clk), .Q(
        \registers[589][6] ) );
  EDFFX1 \registers_reg[589][5]  ( .D(n8270), .E(n76), .CK(clk), .Q(
        \registers[589][5] ) );
  EDFFX1 \registers_reg[589][4]  ( .D(n8212), .E(n76), .CK(clk), .Q(
        \registers[589][4] ) );
  EDFFX1 \registers_reg[589][3]  ( .D(n8167), .E(n76), .CK(clk), .Q(
        \registers[589][3] ) );
  EDFFX1 \registers_reg[589][2]  ( .D(n8119), .E(n76), .CK(clk), .Q(
        \registers[589][2] ) );
  EDFFX1 \registers_reg[589][1]  ( .D(n8063), .E(n76), .CK(clk), .Q(
        \registers[589][1] ) );
  EDFFX1 \registers_reg[589][0]  ( .D(n8001), .E(n76), .CK(clk), .Q(
        \registers[589][0] ) );
  EDFFX1 \registers_reg[585][7]  ( .D(n8387), .E(n72), .CK(clk), .Q(
        \registers[585][7] ) );
  EDFFX1 \registers_reg[585][6]  ( .D(n8329), .E(n72), .CK(clk), .Q(
        \registers[585][6] ) );
  EDFFX1 \registers_reg[585][5]  ( .D(n8271), .E(n72), .CK(clk), .Q(
        \registers[585][5] ) );
  EDFFX1 \registers_reg[585][4]  ( .D(n8213), .E(n72), .CK(clk), .Q(
        \registers[585][4] ) );
  EDFFX1 \registers_reg[585][3]  ( .D(n8168), .E(n72), .CK(clk), .Q(
        \registers[585][3] ) );
  EDFFX1 \registers_reg[585][2]  ( .D(n8117), .E(n72), .CK(clk), .Q(
        \registers[585][2] ) );
  EDFFX1 \registers_reg[585][1]  ( .D(n8061), .E(n72), .CK(clk), .Q(
        \registers[585][1] ) );
  EDFFX1 \registers_reg[585][0]  ( .D(n8002), .E(n72), .CK(clk), .Q(
        \registers[585][0] ) );
  EDFFX1 \registers_reg[581][7]  ( .D(n8388), .E(n278), .CK(clk), .Q(
        \registers[581][7] ) );
  EDFFX1 \registers_reg[581][6]  ( .D(n8330), .E(n278), .CK(clk), .Q(
        \registers[581][6] ) );
  EDFFX1 \registers_reg[581][5]  ( .D(n8272), .E(n278), .CK(clk), .Q(
        \registers[581][5] ) );
  EDFFX1 \registers_reg[581][4]  ( .D(n8214), .E(n278), .CK(clk), .Q(
        \registers[581][4] ) );
  EDFFX1 \registers_reg[581][3]  ( .D(n8169), .E(n278), .CK(clk), .Q(
        \registers[581][3] ) );
  EDFFX1 \registers_reg[581][2]  ( .D(n8118), .E(n278), .CK(clk), .Q(
        \registers[581][2] ) );
  EDFFX1 \registers_reg[581][1]  ( .D(n8062), .E(n278), .CK(clk), .Q(
        \registers[581][1] ) );
  EDFFX1 \registers_reg[581][0]  ( .D(n8003), .E(n278), .CK(clk), .Q(
        \registers[581][0] ) );
  EDFFX1 \registers_reg[577][7]  ( .D(n8386), .E(n274), .CK(clk), .Q(
        \registers[577][7] ) );
  EDFFX1 \registers_reg[577][6]  ( .D(n8328), .E(n274), .CK(clk), .Q(
        \registers[577][6] ) );
  EDFFX1 \registers_reg[577][5]  ( .D(n8270), .E(n274), .CK(clk), .Q(
        \registers[577][5] ) );
  EDFFX1 \registers_reg[577][4]  ( .D(n8212), .E(n274), .CK(clk), .Q(
        \registers[577][4] ) );
  EDFFX1 \registers_reg[577][3]  ( .D(n8167), .E(n274), .CK(clk), .Q(
        \registers[577][3] ) );
  EDFFX1 \registers_reg[577][2]  ( .D(n8116), .E(n274), .CK(clk), .Q(
        \registers[577][2] ) );
  EDFFX1 \registers_reg[577][1]  ( .D(n8060), .E(n274), .CK(clk), .Q(
        \registers[577][1] ) );
  EDFFX1 \registers_reg[577][0]  ( .D(n7998), .E(n274), .CK(clk), .Q(
        \registers[577][0] ) );
  EDFFX1 \registers_reg[573][7]  ( .D(n8384), .E(n763), .CK(clk), .Q(
        \registers[573][7] ) );
  EDFFX1 \registers_reg[573][6]  ( .D(n8326), .E(n763), .CK(clk), .Q(
        \registers[573][6] ) );
  EDFFX1 \registers_reg[573][5]  ( .D(n8268), .E(n763), .CK(clk), .Q(
        \registers[573][5] ) );
  EDFFX1 \registers_reg[573][4]  ( .D(n8210), .E(n763), .CK(clk), .Q(
        \registers[573][4] ) );
  EDFFX1 \registers_reg[573][3]  ( .D(n8169), .E(n763), .CK(clk), .Q(
        \registers[573][3] ) );
  EDFFX1 \registers_reg[573][2]  ( .D(n8115), .E(n763), .CK(clk), .Q(
        \registers[573][2] ) );
  EDFFX1 \registers_reg[573][1]  ( .D(n8059), .E(n763), .CK(clk), .Q(
        \registers[573][1] ) );
  EDFFX1 \registers_reg[573][0]  ( .D(n8000), .E(n763), .CK(clk), .Q(
        \registers[573][0] ) );
  EDFFX1 \registers_reg[569][7]  ( .D(n8883), .E(n759), .CK(clk), .Q(
        \registers[569][7] ) );
  EDFFX1 \registers_reg[569][6]  ( .D(n8854), .E(n759), .CK(clk), .Q(
        \registers[569][6] ) );
  EDFFX1 \registers_reg[569][5]  ( .D(n8825), .E(n759), .CK(clk), .Q(
        \registers[569][5] ) );
  EDFFX1 \registers_reg[569][4]  ( .D(n8796), .E(n759), .CK(clk), .Q(
        \registers[569][4] ) );
  EDFFX1 \registers_reg[569][3]  ( .D(n8167), .E(n759), .CK(clk), .Q(
        \registers[569][3] ) );
  EDFFX1 \registers_reg[569][2]  ( .D(n8116), .E(n759), .CK(clk), .Q(
        \registers[569][2] ) );
  EDFFX1 \registers_reg[569][1]  ( .D(n8060), .E(n759), .CK(clk), .Q(
        \registers[569][1] ) );
  EDFFX1 \registers_reg[569][0]  ( .D(n7998), .E(n759), .CK(clk), .Q(
        \registers[569][0] ) );
  EDFFX1 \registers_reg[565][7]  ( .D(n8385), .E(n755), .CK(clk), .Q(
        \registers[565][7] ) );
  EDFFX1 \registers_reg[565][6]  ( .D(n8327), .E(n755), .CK(clk), .Q(
        \registers[565][6] ) );
  EDFFX1 \registers_reg[565][5]  ( .D(n8269), .E(n755), .CK(clk), .Q(
        \registers[565][5] ) );
  EDFFX1 \registers_reg[565][4]  ( .D(n8211), .E(n755), .CK(clk), .Q(
        \registers[565][4] ) );
  EDFFX1 \registers_reg[565][3]  ( .D(n8168), .E(n755), .CK(clk), .Q(
        \registers[565][3] ) );
  EDFFX1 \registers_reg[565][2]  ( .D(n8114), .E(n755), .CK(clk), .Q(
        \registers[565][2] ) );
  EDFFX1 \registers_reg[565][1]  ( .D(n8058), .E(n755), .CK(clk), .Q(
        \registers[565][1] ) );
  EDFFX1 \registers_reg[565][0]  ( .D(n7999), .E(n755), .CK(clk), .Q(
        \registers[565][0] ) );
  EDFFX1 \registers_reg[561][7]  ( .D(n8384), .E(n68), .CK(clk), .Q(
        \registers[561][7] ) );
  EDFFX1 \registers_reg[561][6]  ( .D(n8326), .E(n68), .CK(clk), .Q(
        \registers[561][6] ) );
  EDFFX1 \registers_reg[561][5]  ( .D(n8268), .E(n68), .CK(clk), .Q(
        \registers[561][5] ) );
  EDFFX1 \registers_reg[561][4]  ( .D(n8210), .E(n68), .CK(clk), .Q(
        \registers[561][4] ) );
  EDFFX1 \registers_reg[561][3]  ( .D(n8166), .E(n68), .CK(clk), .Q(
        \registers[561][3] ) );
  EDFFX1 \registers_reg[561][2]  ( .D(n8115), .E(n68), .CK(clk), .Q(
        \registers[561][2] ) );
  EDFFX1 \registers_reg[561][1]  ( .D(n8059), .E(n68), .CK(clk), .Q(
        \registers[561][1] ) );
  EDFFX1 \registers_reg[561][0]  ( .D(n8000), .E(n68), .CK(clk), .Q(
        \registers[561][0] ) );
  EDFFX1 \registers_reg[557][7]  ( .D(n8433), .E(n64), .CK(clk), .Q(
        \registers[557][7] ) );
  EDFFX1 \registers_reg[557][6]  ( .D(n8375), .E(n64), .CK(clk), .Q(
        \registers[557][6] ) );
  EDFFX1 \registers_reg[557][5]  ( .D(n8317), .E(n64), .CK(clk), .Q(
        \registers[557][5] ) );
  EDFFX1 \registers_reg[557][4]  ( .D(n8259), .E(n64), .CK(clk), .Q(
        \registers[557][4] ) );
  EDFFX1 \registers_reg[557][3]  ( .D(n8164), .E(n64), .CK(clk), .Q(
        \registers[557][3] ) );
  EDFFX1 \registers_reg[557][2]  ( .D(n8116), .E(n64), .CK(clk), .Q(
        \registers[557][2] ) );
  EDFFX1 \registers_reg[557][1]  ( .D(n8060), .E(n64), .CK(clk), .Q(
        \registers[557][1] ) );
  EDFFX1 \registers_reg[557][0]  ( .D(n7998), .E(n64), .CK(clk), .Q(
        \registers[557][0] ) );
  EDFFX1 \registers_reg[553][7]  ( .D(n8385), .E(n60), .CK(clk), .Q(
        \registers[553][7] ) );
  EDFFX1 \registers_reg[553][6]  ( .D(n8327), .E(n60), .CK(clk), .Q(
        \registers[553][6] ) );
  EDFFX1 \registers_reg[553][5]  ( .D(n8269), .E(n60), .CK(clk), .Q(
        \registers[553][5] ) );
  EDFFX1 \registers_reg[553][4]  ( .D(n8211), .E(n60), .CK(clk), .Q(
        \registers[553][4] ) );
  EDFFX1 \registers_reg[553][3]  ( .D(n8165), .E(n60), .CK(clk), .Q(
        \registers[553][3] ) );
  EDFFX1 \registers_reg[553][2]  ( .D(n8114), .E(n60), .CK(clk), .Q(
        \registers[553][2] ) );
  EDFFX1 \registers_reg[553][1]  ( .D(n8058), .E(n60), .CK(clk), .Q(
        \registers[553][1] ) );
  EDFFX1 \registers_reg[553][0]  ( .D(n7999), .E(n60), .CK(clk), .Q(
        \registers[553][0] ) );
  EDFFX1 \registers_reg[549][7]  ( .D(n8384), .E(n271), .CK(clk), .Q(
        \registers[549][7] ) );
  EDFFX1 \registers_reg[549][6]  ( .D(n8326), .E(n271), .CK(clk), .Q(
        \registers[549][6] ) );
  EDFFX1 \registers_reg[549][5]  ( .D(n8268), .E(n271), .CK(clk), .Q(
        \registers[549][5] ) );
  EDFFX1 \registers_reg[549][4]  ( .D(n8210), .E(n271), .CK(clk), .Q(
        \registers[549][4] ) );
  EDFFX1 \registers_reg[549][3]  ( .D(n8166), .E(n271), .CK(clk), .Q(
        \registers[549][3] ) );
  EDFFX1 \registers_reg[549][2]  ( .D(n8115), .E(n271), .CK(clk), .Q(
        \registers[549][2] ) );
  EDFFX1 \registers_reg[549][1]  ( .D(n8059), .E(n271), .CK(clk), .Q(
        \registers[549][1] ) );
  EDFFX1 \registers_reg[549][0]  ( .D(n8000), .E(n271), .CK(clk), .Q(
        \registers[549][0] ) );
  EDFFX1 \registers_reg[545][7]  ( .D(n8434), .E(n267), .CK(clk), .Q(
        \registers[545][7] ) );
  EDFFX1 \registers_reg[545][6]  ( .D(n8376), .E(n267), .CK(clk), .Q(
        \registers[545][6] ) );
  EDFFX1 \registers_reg[545][5]  ( .D(n8318), .E(n267), .CK(clk), .Q(
        \registers[545][5] ) );
  EDFFX1 \registers_reg[545][4]  ( .D(n8260), .E(n267), .CK(clk), .Q(
        \registers[545][4] ) );
  EDFFX1 \registers_reg[545][3]  ( .D(n8164), .E(n267), .CK(clk), .Q(
        \registers[545][3] ) );
  EDFFX1 \registers_reg[545][2]  ( .D(n8116), .E(n267), .CK(clk), .Q(
        \registers[545][2] ) );
  EDFFX1 \registers_reg[545][1]  ( .D(n8060), .E(n267), .CK(clk), .Q(
        \registers[545][1] ) );
  EDFFX1 \registers_reg[545][0]  ( .D(n7998), .E(n267), .CK(clk), .Q(
        \registers[545][0] ) );
  EDFFX1 \registers_reg[541][7]  ( .D(n8385), .E(n751), .CK(clk), .Q(
        \registers[541][7] ) );
  EDFFX1 \registers_reg[541][6]  ( .D(n8327), .E(n751), .CK(clk), .Q(
        \registers[541][6] ) );
  EDFFX1 \registers_reg[541][5]  ( .D(n8269), .E(n751), .CK(clk), .Q(
        \registers[541][5] ) );
  EDFFX1 \registers_reg[541][4]  ( .D(n8211), .E(n751), .CK(clk), .Q(
        \registers[541][4] ) );
  EDFFX1 \registers_reg[541][3]  ( .D(n8165), .E(n751), .CK(clk), .Q(
        \registers[541][3] ) );
  EDFFX1 \registers_reg[541][2]  ( .D(n8114), .E(n751), .CK(clk), .Q(
        \registers[541][2] ) );
  EDFFX1 \registers_reg[541][1]  ( .D(n8058), .E(n751), .CK(clk), .Q(
        \registers[541][1] ) );
  EDFFX1 \registers_reg[541][0]  ( .D(n7999), .E(n751), .CK(clk), .Q(
        \registers[541][0] ) );
  EDFFX1 \registers_reg[537][7]  ( .D(n8384), .E(n747), .CK(clk), .Q(
        \registers[537][7] ) );
  EDFFX1 \registers_reg[537][6]  ( .D(n8326), .E(n747), .CK(clk), .Q(
        \registers[537][6] ) );
  EDFFX1 \registers_reg[537][5]  ( .D(n8268), .E(n747), .CK(clk), .Q(
        \registers[537][5] ) );
  EDFFX1 \registers_reg[537][4]  ( .D(n8210), .E(n747), .CK(clk), .Q(
        \registers[537][4] ) );
  EDFFX1 \registers_reg[537][3]  ( .D(n8166), .E(n747), .CK(clk), .Q(
        \registers[537][3] ) );
  EDFFX1 \registers_reg[537][2]  ( .D(n8115), .E(n747), .CK(clk), .Q(
        \registers[537][2] ) );
  EDFFX1 \registers_reg[537][1]  ( .D(n8059), .E(n747), .CK(clk), .Q(
        \registers[537][1] ) );
  EDFFX1 \registers_reg[537][0]  ( .D(n8000), .E(n747), .CK(clk), .Q(
        \registers[537][0] ) );
  EDFFX1 \registers_reg[533][7]  ( .D(n8875), .E(n743), .CK(clk), .Q(
        \registers[533][7] ) );
  EDFFX1 \registers_reg[533][6]  ( .D(n8846), .E(n743), .CK(clk), .Q(
        \registers[533][6] ) );
  EDFFX1 \registers_reg[533][5]  ( .D(n8817), .E(n743), .CK(clk), .Q(
        \registers[533][5] ) );
  EDFFX1 \registers_reg[533][4]  ( .D(n8788), .E(n743), .CK(clk), .Q(
        \registers[533][4] ) );
  EDFFX1 \registers_reg[533][3]  ( .D(n8164), .E(n743), .CK(clk), .Q(
        \registers[533][3] ) );
  EDFFX1 \registers_reg[533][2]  ( .D(n8116), .E(n743), .CK(clk), .Q(
        \registers[533][2] ) );
  EDFFX1 \registers_reg[533][1]  ( .D(n8060), .E(n743), .CK(clk), .Q(
        \registers[533][1] ) );
  EDFFX1 \registers_reg[533][0]  ( .D(n7998), .E(n743), .CK(clk), .Q(
        \registers[533][0] ) );
  EDFFX1 \registers_reg[529][7]  ( .D(n8385), .E(n56), .CK(clk), .Q(
        \registers[529][7] ) );
  EDFFX1 \registers_reg[529][6]  ( .D(n8327), .E(n56), .CK(clk), .Q(
        \registers[529][6] ) );
  EDFFX1 \registers_reg[529][5]  ( .D(n8269), .E(n56), .CK(clk), .Q(
        \registers[529][5] ) );
  EDFFX1 \registers_reg[529][4]  ( .D(n8211), .E(n56), .CK(clk), .Q(
        \registers[529][4] ) );
  EDFFX1 \registers_reg[529][3]  ( .D(n8165), .E(n56), .CK(clk), .Q(
        \registers[529][3] ) );
  EDFFX1 \registers_reg[529][2]  ( .D(n8111), .E(n56), .CK(clk), .Q(
        \registers[529][2] ) );
  EDFFX1 \registers_reg[529][1]  ( .D(n8055), .E(n56), .CK(clk), .Q(
        \registers[529][1] ) );
  EDFFX1 \registers_reg[529][0]  ( .D(n7999), .E(n56), .CK(clk), .Q(
        \registers[529][0] ) );
  EDFFX1 \registers_reg[525][7]  ( .D(n8382), .E(n51), .CK(clk), .Q(
        \registers[525][7] ) );
  EDFFX1 \registers_reg[525][6]  ( .D(n8324), .E(n51), .CK(clk), .Q(
        \registers[525][6] ) );
  EDFFX1 \registers_reg[525][5]  ( .D(n8266), .E(n51), .CK(clk), .Q(
        \registers[525][5] ) );
  EDFFX1 \registers_reg[525][4]  ( .D(n8208), .E(n51), .CK(clk), .Q(
        \registers[525][4] ) );
  EDFFX1 \registers_reg[525][3]  ( .D(n8166), .E(n51), .CK(clk), .Q(
        \registers[525][3] ) );
  EDFFX1 \registers_reg[525][2]  ( .D(n8112), .E(n51), .CK(clk), .Q(
        \registers[525][2] ) );
  EDFFX1 \registers_reg[525][1]  ( .D(n8056), .E(n51), .CK(clk), .Q(
        \registers[525][1] ) );
  EDFFX1 \registers_reg[525][0]  ( .D(n8676), .E(n51), .CK(clk), .Q(
        \registers[525][0] ) );
  EDFFX1 \registers_reg[521][7]  ( .D(n8383), .E(n47), .CK(clk), .Q(
        \registers[521][7] ) );
  EDFFX1 \registers_reg[521][6]  ( .D(n8325), .E(n47), .CK(clk), .Q(
        \registers[521][6] ) );
  EDFFX1 \registers_reg[521][5]  ( .D(n8267), .E(n47), .CK(clk), .Q(
        \registers[521][5] ) );
  EDFFX1 \registers_reg[521][4]  ( .D(n8209), .E(n47), .CK(clk), .Q(
        \registers[521][4] ) );
  EDFFX1 \registers_reg[521][3]  ( .D(n8164), .E(n47), .CK(clk), .Q(
        \registers[521][3] ) );
  EDFFX1 \registers_reg[521][2]  ( .D(n8113), .E(n47), .CK(clk), .Q(
        \registers[521][2] ) );
  EDFFX1 \registers_reg[521][1]  ( .D(n8057), .E(n47), .CK(clk), .Q(
        \registers[521][1] ) );
  EDFFX1 \registers_reg[521][0]  ( .D(n7996), .E(n47), .CK(clk), .Q(
        \registers[521][0] ) );
  EDFFX1 \registers_reg[517][7]  ( .D(n8381), .E(n264), .CK(clk), .Q(
        \registers[517][7] ) );
  EDFFX1 \registers_reg[517][6]  ( .D(n8323), .E(n264), .CK(clk), .Q(
        \registers[517][6] ) );
  EDFFX1 \registers_reg[517][5]  ( .D(n8265), .E(n264), .CK(clk), .Q(
        \registers[517][5] ) );
  EDFFX1 \registers_reg[517][4]  ( .D(n8207), .E(n264), .CK(clk), .Q(
        \registers[517][4] ) );
  EDFFX1 \registers_reg[517][3]  ( .D(n8165), .E(n264), .CK(clk), .Q(
        \registers[517][3] ) );
  EDFFX1 \registers_reg[517][2]  ( .D(n8111), .E(n264), .CK(clk), .Q(
        \registers[517][2] ) );
  EDFFX1 \registers_reg[517][1]  ( .D(n8055), .E(n264), .CK(clk), .Q(
        \registers[517][1] ) );
  EDFFX1 \registers_reg[517][0]  ( .D(n7997), .E(n264), .CK(clk), .Q(
        \registers[517][0] ) );
  EDFFX1 \registers_reg[513][7]  ( .D(n8387), .E(n260), .CK(clk), .Q(
        \registers[513][7] ) );
  EDFFX1 \registers_reg[513][6]  ( .D(n8329), .E(n260), .CK(clk), .Q(
        \registers[513][6] ) );
  EDFFX1 \registers_reg[513][5]  ( .D(n8271), .E(n260), .CK(clk), .Q(
        \registers[513][5] ) );
  EDFFX1 \registers_reg[513][4]  ( .D(n8213), .E(n260), .CK(clk), .Q(
        \registers[513][4] ) );
  EDFFX1 \registers_reg[513][3]  ( .D(n8168), .E(n260), .CK(clk), .Q(
        \registers[513][3] ) );
  EDFFX1 \registers_reg[513][2]  ( .D(n8114), .E(n260), .CK(clk), .Q(
        \registers[513][2] ) );
  EDFFX1 \registers_reg[513][1]  ( .D(n8058), .E(n260), .CK(clk), .Q(
        \registers[513][1] ) );
  EDFFX1 \registers_reg[513][0]  ( .D(n8687), .E(n260), .CK(clk), .Q(
        \registers[513][0] ) );
  EDFFX1 \registers_reg[509][7]  ( .D(n8405), .E(n739), .CK(clk), .Q(
        \registers[509][7] ) );
  EDFFX1 \registers_reg[509][6]  ( .D(n8347), .E(n739), .CK(clk), .Q(
        \registers[509][6] ) );
  EDFFX1 \registers_reg[509][5]  ( .D(n8289), .E(n739), .CK(clk), .Q(
        \registers[509][5] ) );
  EDFFX1 \registers_reg[509][4]  ( .D(n8231), .E(n739), .CK(clk), .Q(
        \registers[509][4] ) );
  EDFFX1 \registers_reg[509][3]  ( .D(n8201), .E(n739), .CK(clk), .Q(
        \registers[509][3] ) );
  EDFFX1 \registers_reg[509][2]  ( .D(n8155), .E(n739), .CK(clk), .Q(
        \registers[509][2] ) );
  EDFFX1 \registers_reg[509][1]  ( .D(n8099), .E(n739), .CK(clk), .Q(
        \registers[509][1] ) );
  EDFFX1 \registers_reg[509][0]  ( .D(n8042), .E(n739), .CK(clk), .Q(
        \registers[509][0] ) );
  EDFFX1 \registers_reg[505][7]  ( .D(n8426), .E(n735), .CK(clk), .Q(
        \registers[505][7] ) );
  EDFFX1 \registers_reg[505][6]  ( .D(n8368), .E(n735), .CK(clk), .Q(
        \registers[505][6] ) );
  EDFFX1 \registers_reg[505][5]  ( .D(n8310), .E(n735), .CK(clk), .Q(
        \registers[505][5] ) );
  EDFFX1 \registers_reg[505][4]  ( .D(n8252), .E(n735), .CK(clk), .Q(
        \registers[505][4] ) );
  EDFFX1 \registers_reg[505][3]  ( .D(n8202), .E(n735), .CK(clk), .Q(
        \registers[505][3] ) );
  EDFFX1 \registers_reg[505][2]  ( .D(n8156), .E(n735), .CK(clk), .Q(
        \registers[505][2] ) );
  EDFFX1 \registers_reg[505][1]  ( .D(n8100), .E(n735), .CK(clk), .Q(
        \registers[505][1] ) );
  EDFFX1 \registers_reg[505][0]  ( .D(n8040), .E(n735), .CK(clk), .Q(
        \registers[505][0] ) );
  EDFFX1 \registers_reg[501][7]  ( .D(n8427), .E(n731), .CK(clk), .Q(
        \registers[501][7] ) );
  EDFFX1 \registers_reg[501][6]  ( .D(n8369), .E(n731), .CK(clk), .Q(
        \registers[501][6] ) );
  EDFFX1 \registers_reg[501][5]  ( .D(n8311), .E(n731), .CK(clk), .Q(
        \registers[501][5] ) );
  EDFFX1 \registers_reg[501][4]  ( .D(n8253), .E(n731), .CK(clk), .Q(
        \registers[501][4] ) );
  EDFFX1 \registers_reg[501][3]  ( .D(n8200), .E(n731), .CK(clk), .Q(
        \registers[501][3] ) );
  EDFFX1 \registers_reg[501][2]  ( .D(n8157), .E(n731), .CK(clk), .Q(
        \registers[501][2] ) );
  EDFFX1 \registers_reg[501][1]  ( .D(n8101), .E(n731), .CK(clk), .Q(
        \registers[501][1] ) );
  EDFFX1 \registers_reg[501][0]  ( .D(n8041), .E(n731), .CK(clk), .Q(
        \registers[501][0] ) );
  EDFFX1 \registers_reg[497][7]  ( .D(n8425), .E(n43), .CK(clk), .Q(
        \registers[497][7] ) );
  EDFFX1 \registers_reg[497][6]  ( .D(n8367), .E(n43), .CK(clk), .Q(
        \registers[497][6] ) );
  EDFFX1 \registers_reg[497][5]  ( .D(n8309), .E(n43), .CK(clk), .Q(
        \registers[497][5] ) );
  EDFFX1 \registers_reg[497][4]  ( .D(n8251), .E(n43), .CK(clk), .Q(
        \registers[497][4] ) );
  EDFFX1 \registers_reg[497][3]  ( .D(n8201), .E(n43), .CK(clk), .Q(
        \registers[497][3] ) );
  EDFFX1 \registers_reg[497][2]  ( .D(n8155), .E(n43), .CK(clk), .Q(
        \registers[497][2] ) );
  EDFFX1 \registers_reg[497][1]  ( .D(n8099), .E(n43), .CK(clk), .Q(
        \registers[497][1] ) );
  EDFFX1 \registers_reg[497][0]  ( .D(n8042), .E(n43), .CK(clk), .Q(
        \registers[497][0] ) );
  EDFFX1 \registers_reg[493][7]  ( .D(n8426), .E(n39), .CK(clk), .Q(
        \registers[493][7] ) );
  EDFFX1 \registers_reg[493][6]  ( .D(n8368), .E(n39), .CK(clk), .Q(
        \registers[493][6] ) );
  EDFFX1 \registers_reg[493][5]  ( .D(n8310), .E(n39), .CK(clk), .Q(
        \registers[493][5] ) );
  EDFFX1 \registers_reg[493][4]  ( .D(n8252), .E(n39), .CK(clk), .Q(
        \registers[493][4] ) );
  EDFFX1 \registers_reg[493][3]  ( .D(n8202), .E(n39), .CK(clk), .Q(
        \registers[493][3] ) );
  EDFFX1 \registers_reg[493][2]  ( .D(n8156), .E(n39), .CK(clk), .Q(
        \registers[493][2] ) );
  EDFFX1 \registers_reg[493][1]  ( .D(n8100), .E(n39), .CK(clk), .Q(
        \registers[493][1] ) );
  EDFFX1 \registers_reg[493][0]  ( .D(n8040), .E(n39), .CK(clk), .Q(
        \registers[493][0] ) );
  EDFFX1 \registers_reg[489][7]  ( .D(n8427), .E(n35), .CK(clk), .Q(
        \registers[489][7] ) );
  EDFFX1 \registers_reg[489][6]  ( .D(n8369), .E(n35), .CK(clk), .Q(
        \registers[489][6] ) );
  EDFFX1 \registers_reg[489][5]  ( .D(n8311), .E(n35), .CK(clk), .Q(
        \registers[489][5] ) );
  EDFFX1 \registers_reg[489][4]  ( .D(n8253), .E(n35), .CK(clk), .Q(
        \registers[489][4] ) );
  EDFFX1 \registers_reg[489][3]  ( .D(n8200), .E(n35), .CK(clk), .Q(
        \registers[489][3] ) );
  EDFFX1 \registers_reg[489][2]  ( .D(n8157), .E(n35), .CK(clk), .Q(
        \registers[489][2] ) );
  EDFFX1 \registers_reg[489][1]  ( .D(n8101), .E(n35), .CK(clk), .Q(
        \registers[489][1] ) );
  EDFFX1 \registers_reg[489][0]  ( .D(n8041), .E(n35), .CK(clk), .Q(
        \registers[489][0] ) );
  EDFFX1 \registers_reg[485][7]  ( .D(n8425), .E(n257), .CK(clk), .Q(
        \registers[485][7] ) );
  EDFFX1 \registers_reg[485][6]  ( .D(n8367), .E(n257), .CK(clk), .Q(
        \registers[485][6] ) );
  EDFFX1 \registers_reg[485][5]  ( .D(n8309), .E(n257), .CK(clk), .Q(
        \registers[485][5] ) );
  EDFFX1 \registers_reg[485][4]  ( .D(n8251), .E(n257), .CK(clk), .Q(
        \registers[485][4] ) );
  EDFFX1 \registers_reg[485][3]  ( .D(n8198), .E(n257), .CK(clk), .Q(
        \registers[485][3] ) );
  EDFFX1 \registers_reg[485][2]  ( .D(n8155), .E(n257), .CK(clk), .Q(
        \registers[485][2] ) );
  EDFFX1 \registers_reg[485][1]  ( .D(n8099), .E(n257), .CK(clk), .Q(
        \registers[485][1] ) );
  EDFFX1 \registers_reg[485][0]  ( .D(n8042), .E(n257), .CK(clk), .Q(
        \registers[485][0] ) );
  EDFFX1 \registers_reg[481][7]  ( .D(n8426), .E(n253), .CK(clk), .Q(
        \registers[481][7] ) );
  EDFFX1 \registers_reg[481][6]  ( .D(n8368), .E(n253), .CK(clk), .Q(
        \registers[481][6] ) );
  EDFFX1 \registers_reg[481][5]  ( .D(n8310), .E(n253), .CK(clk), .Q(
        \registers[481][5] ) );
  EDFFX1 \registers_reg[481][4]  ( .D(n8252), .E(n253), .CK(clk), .Q(
        \registers[481][4] ) );
  EDFFX1 \registers_reg[481][3]  ( .D(n8199), .E(n253), .CK(clk), .Q(
        \registers[481][3] ) );
  EDFFX1 \registers_reg[481][2]  ( .D(n8156), .E(n253), .CK(clk), .Q(
        \registers[481][2] ) );
  EDFFX1 \registers_reg[481][1]  ( .D(n8100), .E(n253), .CK(clk), .Q(
        \registers[481][1] ) );
  EDFFX1 \registers_reg[481][0]  ( .D(n8040), .E(n253), .CK(clk), .Q(
        \registers[481][0] ) );
  EDFFX1 \registers_reg[477][7]  ( .D(n8427), .E(n727), .CK(clk), .Q(
        \registers[477][7] ) );
  EDFFX1 \registers_reg[477][6]  ( .D(n8369), .E(n727), .CK(clk), .Q(
        \registers[477][6] ) );
  EDFFX1 \registers_reg[477][5]  ( .D(n8311), .E(n727), .CK(clk), .Q(
        \registers[477][5] ) );
  EDFFX1 \registers_reg[477][4]  ( .D(n8253), .E(n727), .CK(clk), .Q(
        \registers[477][4] ) );
  EDFFX1 \registers_reg[477][3]  ( .D(n8197), .E(n727), .CK(clk), .Q(
        \registers[477][3] ) );
  EDFFX1 \registers_reg[477][2]  ( .D(n8157), .E(n727), .CK(clk), .Q(
        \registers[477][2] ) );
  EDFFX1 \registers_reg[477][1]  ( .D(n8101), .E(n727), .CK(clk), .Q(
        \registers[477][1] ) );
  EDFFX1 \registers_reg[477][0]  ( .D(n8041), .E(n727), .CK(clk), .Q(
        \registers[477][0] ) );
  EDFFX1 \registers_reg[473][7]  ( .D(n8425), .E(n723), .CK(clk), .Q(
        \registers[473][7] ) );
  EDFFX1 \registers_reg[473][6]  ( .D(n8367), .E(n723), .CK(clk), .Q(
        \registers[473][6] ) );
  EDFFX1 \registers_reg[473][5]  ( .D(n8309), .E(n723), .CK(clk), .Q(
        \registers[473][5] ) );
  EDFFX1 \registers_reg[473][4]  ( .D(n8251), .E(n723), .CK(clk), .Q(
        \registers[473][4] ) );
  EDFFX1 \registers_reg[473][3]  ( .D(n8198), .E(n723), .CK(clk), .Q(
        \registers[473][3] ) );
  EDFFX1 \registers_reg[473][2]  ( .D(n8152), .E(n723), .CK(clk), .Q(
        \registers[473][2] ) );
  EDFFX1 \registers_reg[473][1]  ( .D(n8096), .E(n723), .CK(clk), .Q(
        \registers[473][1] ) );
  EDFFX1 \registers_reg[473][0]  ( .D(n8042), .E(n723), .CK(clk), .Q(
        \registers[473][0] ) );
  EDFFX1 \registers_reg[469][7]  ( .D(n8426), .E(n719), .CK(clk), .Q(
        \registers[469][7] ) );
  EDFFX1 \registers_reg[469][6]  ( .D(n8368), .E(n719), .CK(clk), .Q(
        \registers[469][6] ) );
  EDFFX1 \registers_reg[469][5]  ( .D(n8310), .E(n719), .CK(clk), .Q(
        \registers[469][5] ) );
  EDFFX1 \registers_reg[469][4]  ( .D(n8252), .E(n719), .CK(clk), .Q(
        \registers[469][4] ) );
  EDFFX1 \registers_reg[469][3]  ( .D(n8199), .E(n719), .CK(clk), .Q(
        \registers[469][3] ) );
  EDFFX1 \registers_reg[469][2]  ( .D(n8153), .E(n719), .CK(clk), .Q(
        \registers[469][2] ) );
  EDFFX1 \registers_reg[469][1]  ( .D(n8097), .E(n719), .CK(clk), .Q(
        \registers[469][1] ) );
  EDFFX1 \registers_reg[469][0]  ( .D(n8037), .E(n719), .CK(clk), .Q(
        \registers[469][0] ) );
  EDFFX1 \registers_reg[465][7]  ( .D(n8427), .E(n31), .CK(clk), .Q(
        \registers[465][7] ) );
  EDFFX1 \registers_reg[465][6]  ( .D(n8369), .E(n31), .CK(clk), .Q(
        \registers[465][6] ) );
  EDFFX1 \registers_reg[465][5]  ( .D(n8311), .E(n31), .CK(clk), .Q(
        \registers[465][5] ) );
  EDFFX1 \registers_reg[465][4]  ( .D(n8253), .E(n31), .CK(clk), .Q(
        \registers[465][4] ) );
  EDFFX1 \registers_reg[465][3]  ( .D(n8197), .E(n31), .CK(clk), .Q(
        \registers[465][3] ) );
  EDFFX1 \registers_reg[465][2]  ( .D(n8154), .E(n31), .CK(clk), .Q(
        \registers[465][2] ) );
  EDFFX1 \registers_reg[465][1]  ( .D(n8098), .E(n31), .CK(clk), .Q(
        \registers[465][1] ) );
  EDFFX1 \registers_reg[465][0]  ( .D(n8038), .E(n31), .CK(clk), .Q(
        \registers[465][0] ) );
  EDFFX1 \registers_reg[461][7]  ( .D(n8425), .E(n27), .CK(clk), .Q(
        \registers[461][7] ) );
  EDFFX1 \registers_reg[461][6]  ( .D(n8367), .E(n27), .CK(clk), .Q(
        \registers[461][6] ) );
  EDFFX1 \registers_reg[461][5]  ( .D(n8309), .E(n27), .CK(clk), .Q(
        \registers[461][5] ) );
  EDFFX1 \registers_reg[461][4]  ( .D(n8251), .E(n27), .CK(clk), .Q(
        \registers[461][4] ) );
  EDFFX1 \registers_reg[461][3]  ( .D(n8198), .E(n27), .CK(clk), .Q(
        \registers[461][3] ) );
  EDFFX1 \registers_reg[461][2]  ( .D(n8152), .E(n27), .CK(clk), .Q(
        \registers[461][2] ) );
  EDFFX1 \registers_reg[461][1]  ( .D(n8096), .E(n27), .CK(clk), .Q(
        \registers[461][1] ) );
  EDFFX1 \registers_reg[461][0]  ( .D(n8039), .E(n27), .CK(clk), .Q(
        \registers[461][0] ) );
  EDFFX1 \registers_reg[457][7]  ( .D(n8426), .E(n23), .CK(clk), .Q(
        \registers[457][7] ) );
  EDFFX1 \registers_reg[457][6]  ( .D(n8368), .E(n23), .CK(clk), .Q(
        \registers[457][6] ) );
  EDFFX1 \registers_reg[457][5]  ( .D(n8310), .E(n23), .CK(clk), .Q(
        \registers[457][5] ) );
  EDFFX1 \registers_reg[457][4]  ( .D(n8252), .E(n23), .CK(clk), .Q(
        \registers[457][4] ) );
  EDFFX1 \registers_reg[457][3]  ( .D(n8199), .E(n23), .CK(clk), .Q(
        \registers[457][3] ) );
  EDFFX1 \registers_reg[457][2]  ( .D(n8153), .E(n23), .CK(clk), .Q(
        \registers[457][2] ) );
  EDFFX1 \registers_reg[457][1]  ( .D(n8097), .E(n23), .CK(clk), .Q(
        \registers[457][1] ) );
  EDFFX1 \registers_reg[457][0]  ( .D(n8037), .E(n23), .CK(clk), .Q(
        \registers[457][0] ) );
  EDFFX1 \registers_reg[453][7]  ( .D(n8422), .E(n250), .CK(clk), .Q(
        \registers[453][7] ) );
  EDFFX1 \registers_reg[453][6]  ( .D(n8364), .E(n250), .CK(clk), .Q(
        \registers[453][6] ) );
  EDFFX1 \registers_reg[453][5]  ( .D(n8306), .E(n250), .CK(clk), .Q(
        \registers[453][5] ) );
  EDFFX1 \registers_reg[453][4]  ( .D(n8248), .E(n250), .CK(clk), .Q(
        \registers[453][4] ) );
  EDFFX1 \registers_reg[453][3]  ( .D(n8197), .E(n250), .CK(clk), .Q(
        \registers[453][3] ) );
  EDFFX1 \registers_reg[453][2]  ( .D(n8154), .E(n250), .CK(clk), .Q(
        \registers[453][2] ) );
  EDFFX1 \registers_reg[453][1]  ( .D(n8098), .E(n250), .CK(clk), .Q(
        \registers[453][1] ) );
  EDFFX1 \registers_reg[453][0]  ( .D(n8038), .E(n250), .CK(clk), .Q(
        \registers[453][0] ) );
  EDFFX1 \registers_reg[449][7]  ( .D(n8423), .E(n246), .CK(clk), .Q(
        \registers[449][7] ) );
  EDFFX1 \registers_reg[449][6]  ( .D(n8365), .E(n246), .CK(clk), .Q(
        \registers[449][6] ) );
  EDFFX1 \registers_reg[449][5]  ( .D(n8307), .E(n246), .CK(clk), .Q(
        \registers[449][5] ) );
  EDFFX1 \registers_reg[449][4]  ( .D(n8249), .E(n246), .CK(clk), .Q(
        \registers[449][4] ) );
  EDFFX1 \registers_reg[449][3]  ( .D(n8198), .E(n246), .CK(clk), .Q(
        \registers[449][3] ) );
  EDFFX1 \registers_reg[449][2]  ( .D(n8152), .E(n246), .CK(clk), .Q(
        \registers[449][2] ) );
  EDFFX1 \registers_reg[449][1]  ( .D(n8096), .E(n246), .CK(clk), .Q(
        \registers[449][1] ) );
  EDFFX1 \registers_reg[449][0]  ( .D(n8039), .E(n246), .CK(clk), .Q(
        \registers[449][0] ) );
  EDFFX1 \registers_reg[445][7]  ( .D(n8422), .E(n715), .CK(clk), .Q(
        \registers[445][7] ) );
  EDFFX1 \registers_reg[445][6]  ( .D(n8364), .E(n715), .CK(clk), .Q(
        \registers[445][6] ) );
  EDFFX1 \registers_reg[445][5]  ( .D(n8306), .E(n715), .CK(clk), .Q(
        \registers[445][5] ) );
  EDFFX1 \registers_reg[445][4]  ( .D(n8248), .E(n715), .CK(clk), .Q(
        \registers[445][4] ) );
  EDFFX1 \registers_reg[445][3]  ( .D(n8197), .E(n715), .CK(clk), .Q(
        \registers[445][3] ) );
  EDFFX1 \registers_reg[445][2]  ( .D(n8154), .E(n715), .CK(clk), .Q(
        \registers[445][2] ) );
  EDFFX1 \registers_reg[445][1]  ( .D(n8098), .E(n715), .CK(clk), .Q(
        \registers[445][1] ) );
  EDFFX1 \registers_reg[445][0]  ( .D(n8038), .E(n715), .CK(clk), .Q(
        \registers[445][0] ) );
  EDFFX1 \registers_reg[441][7]  ( .D(n8423), .E(n711), .CK(clk), .Q(
        \registers[441][7] ) );
  EDFFX1 \registers_reg[441][6]  ( .D(n8365), .E(n711), .CK(clk), .Q(
        \registers[441][6] ) );
  EDFFX1 \registers_reg[441][5]  ( .D(n8307), .E(n711), .CK(clk), .Q(
        \registers[441][5] ) );
  EDFFX1 \registers_reg[441][4]  ( .D(n8249), .E(n711), .CK(clk), .Q(
        \registers[441][4] ) );
  EDFFX1 \registers_reg[441][3]  ( .D(n8198), .E(n711), .CK(clk), .Q(
        \registers[441][3] ) );
  EDFFX1 \registers_reg[441][2]  ( .D(n8152), .E(n711), .CK(clk), .Q(
        \registers[441][2] ) );
  EDFFX1 \registers_reg[441][1]  ( .D(n8096), .E(n711), .CK(clk), .Q(
        \registers[441][1] ) );
  EDFFX1 \registers_reg[441][0]  ( .D(n8039), .E(n711), .CK(clk), .Q(
        \registers[441][0] ) );
  EDFFX1 \registers_reg[437][7]  ( .D(n8424), .E(n707), .CK(clk), .Q(
        \registers[437][7] ) );
  EDFFX1 \registers_reg[437][6]  ( .D(n8366), .E(n707), .CK(clk), .Q(
        \registers[437][6] ) );
  EDFFX1 \registers_reg[437][5]  ( .D(n8308), .E(n707), .CK(clk), .Q(
        \registers[437][5] ) );
  EDFFX1 \registers_reg[437][4]  ( .D(n8250), .E(n707), .CK(clk), .Q(
        \registers[437][4] ) );
  EDFFX1 \registers_reg[437][3]  ( .D(n8199), .E(n707), .CK(clk), .Q(
        \registers[437][3] ) );
  EDFFX1 \registers_reg[437][2]  ( .D(n8153), .E(n707), .CK(clk), .Q(
        \registers[437][2] ) );
  EDFFX1 \registers_reg[437][1]  ( .D(n8097), .E(n707), .CK(clk), .Q(
        \registers[437][1] ) );
  EDFFX1 \registers_reg[437][0]  ( .D(n8037), .E(n707), .CK(clk), .Q(
        \registers[437][0] ) );
  EDFFX1 \registers_reg[433][7]  ( .D(n8422), .E(n19), .CK(clk), .Q(
        \registers[433][7] ) );
  EDFFX1 \registers_reg[433][6]  ( .D(n8364), .E(n19), .CK(clk), .Q(
        \registers[433][6] ) );
  EDFFX1 \registers_reg[433][5]  ( .D(n8306), .E(n19), .CK(clk), .Q(
        \registers[433][5] ) );
  EDFFX1 \registers_reg[433][4]  ( .D(n8248), .E(n19), .CK(clk), .Q(
        \registers[433][4] ) );
  EDFFX1 \registers_reg[433][3]  ( .D(n8197), .E(n19), .CK(clk), .Q(
        \registers[433][3] ) );
  EDFFX1 \registers_reg[433][2]  ( .D(n8154), .E(n19), .CK(clk), .Q(
        \registers[433][2] ) );
  EDFFX1 \registers_reg[433][1]  ( .D(n8098), .E(n19), .CK(clk), .Q(
        \registers[433][1] ) );
  EDFFX1 \registers_reg[433][0]  ( .D(n8038), .E(n19), .CK(clk), .Q(
        \registers[433][0] ) );
  EDFFX1 \registers_reg[429][7]  ( .D(n8423), .E(n15), .CK(clk), .Q(
        \registers[429][7] ) );
  EDFFX1 \registers_reg[429][6]  ( .D(n8365), .E(n15), .CK(clk), .Q(
        \registers[429][6] ) );
  EDFFX1 \registers_reg[429][5]  ( .D(n8307), .E(n15), .CK(clk), .Q(
        \registers[429][5] ) );
  EDFFX1 \registers_reg[429][4]  ( .D(n8249), .E(n15), .CK(clk), .Q(
        \registers[429][4] ) );
  EDFFX1 \registers_reg[429][3]  ( .D(n8198), .E(n15), .CK(clk), .Q(
        \registers[429][3] ) );
  EDFFX1 \registers_reg[429][2]  ( .D(n8152), .E(n15), .CK(clk), .Q(
        \registers[429][2] ) );
  EDFFX1 \registers_reg[429][1]  ( .D(n8096), .E(n15), .CK(clk), .Q(
        \registers[429][1] ) );
  EDFFX1 \registers_reg[429][0]  ( .D(n8039), .E(n15), .CK(clk), .Q(
        \registers[429][0] ) );
  EDFFX1 \registers_reg[425][7]  ( .D(n8424), .E(n11), .CK(clk), .Q(
        \registers[425][7] ) );
  EDFFX1 \registers_reg[425][6]  ( .D(n8366), .E(n11), .CK(clk), .Q(
        \registers[425][6] ) );
  EDFFX1 \registers_reg[425][5]  ( .D(n8308), .E(n11), .CK(clk), .Q(
        \registers[425][5] ) );
  EDFFX1 \registers_reg[425][4]  ( .D(n8250), .E(n11), .CK(clk), .Q(
        \registers[425][4] ) );
  EDFFX1 \registers_reg[425][3]  ( .D(n8199), .E(n11), .CK(clk), .Q(
        \registers[425][3] ) );
  EDFFX1 \registers_reg[425][2]  ( .D(n8153), .E(n11), .CK(clk), .Q(
        \registers[425][2] ) );
  EDFFX1 \registers_reg[425][1]  ( .D(n8097), .E(n11), .CK(clk), .Q(
        \registers[425][1] ) );
  EDFFX1 \registers_reg[425][0]  ( .D(n8037), .E(n11), .CK(clk), .Q(
        \registers[425][0] ) );
  EDFFX1 \registers_reg[421][7]  ( .D(n8422), .E(n243), .CK(clk), .Q(
        \registers[421][7] ) );
  EDFFX1 \registers_reg[421][6]  ( .D(n8364), .E(n243), .CK(clk), .Q(
        \registers[421][6] ) );
  EDFFX1 \registers_reg[421][5]  ( .D(n8306), .E(n243), .CK(clk), .Q(
        \registers[421][5] ) );
  EDFFX1 \registers_reg[421][4]  ( .D(n8248), .E(n243), .CK(clk), .Q(
        \registers[421][4] ) );
  EDFFX1 \registers_reg[421][3]  ( .D(n8194), .E(n243), .CK(clk), .Q(
        \registers[421][3] ) );
  EDFFX1 \registers_reg[421][2]  ( .D(n8732), .E(n243), .CK(clk), .Q(
        \registers[421][2] ) );
  EDFFX1 \registers_reg[421][1]  ( .D(n8704), .E(n243), .CK(clk), .Q(
        \registers[421][1] ) );
  EDFFX1 \registers_reg[421][0]  ( .D(n8035), .E(n243), .CK(clk), .Q(
        \registers[421][0] ) );
  EDFFX1 \registers_reg[417][7]  ( .D(n8423), .E(n239), .CK(clk), .Q(
        \registers[417][7] ) );
  EDFFX1 \registers_reg[417][6]  ( .D(n8365), .E(n239), .CK(clk), .Q(
        \registers[417][6] ) );
  EDFFX1 \registers_reg[417][5]  ( .D(n8307), .E(n239), .CK(clk), .Q(
        \registers[417][5] ) );
  EDFFX1 \registers_reg[417][4]  ( .D(n8249), .E(n239), .CK(clk), .Q(
        \registers[417][4] ) );
  EDFFX1 \registers_reg[417][3]  ( .D(n8195), .E(n239), .CK(clk), .Q(
        \registers[417][3] ) );
  EDFFX1 \registers_reg[417][2]  ( .D(n8150), .E(n239), .CK(clk), .Q(
        \registers[417][2] ) );
  EDFFX1 \registers_reg[417][1]  ( .D(n8094), .E(n239), .CK(clk), .Q(
        \registers[417][1] ) );
  EDFFX1 \registers_reg[417][0]  ( .D(n8036), .E(n239), .CK(clk), .Q(
        \registers[417][0] ) );
  EDFFX1 \registers_reg[413][7]  ( .D(n8424), .E(n703), .CK(clk), .Q(
        \registers[413][7] ) );
  EDFFX1 \registers_reg[413][6]  ( .D(n8366), .E(n703), .CK(clk), .Q(
        \registers[413][6] ) );
  EDFFX1 \registers_reg[413][5]  ( .D(n8308), .E(n703), .CK(clk), .Q(
        \registers[413][5] ) );
  EDFFX1 \registers_reg[413][4]  ( .D(n8250), .E(n703), .CK(clk), .Q(
        \registers[413][4] ) );
  EDFFX1 \registers_reg[413][3]  ( .D(n8196), .E(n703), .CK(clk), .Q(
        \registers[413][3] ) );
  EDFFX1 \registers_reg[413][2]  ( .D(n8151), .E(n703), .CK(clk), .Q(
        \registers[413][2] ) );
  EDFFX1 \registers_reg[413][1]  ( .D(n8095), .E(n703), .CK(clk), .Q(
        \registers[413][1] ) );
  EDFFX1 \registers_reg[413][0]  ( .D(n8034), .E(n703), .CK(clk), .Q(
        \registers[413][0] ) );
  EDFFX1 \registers_reg[409][7]  ( .D(n8422), .E(n699), .CK(clk), .Q(
        \registers[409][7] ) );
  EDFFX1 \registers_reg[409][6]  ( .D(n8364), .E(n699), .CK(clk), .Q(
        \registers[409][6] ) );
  EDFFX1 \registers_reg[409][5]  ( .D(n8306), .E(n699), .CK(clk), .Q(
        \registers[409][5] ) );
  EDFFX1 \registers_reg[409][4]  ( .D(n8248), .E(n699), .CK(clk), .Q(
        \registers[409][4] ) );
  EDFFX1 \registers_reg[409][3]  ( .D(n8194), .E(n699), .CK(clk), .Q(
        \registers[409][3] ) );
  EDFFX1 \registers_reg[409][2]  ( .D(n8731), .E(n699), .CK(clk), .Q(
        \registers[409][2] ) );
  EDFFX1 \registers_reg[409][1]  ( .D(n8703), .E(n699), .CK(clk), .Q(
        \registers[409][1] ) );
  EDFFX1 \registers_reg[409][0]  ( .D(n8035), .E(n699), .CK(clk), .Q(
        \registers[409][0] ) );
  EDFFX1 \registers_reg[405][7]  ( .D(n8421), .E(n695), .CK(clk), .Q(
        \registers[405][7] ) );
  EDFFX1 \registers_reg[405][6]  ( .D(n8363), .E(n695), .CK(clk), .Q(
        \registers[405][6] ) );
  EDFFX1 \registers_reg[405][5]  ( .D(n8305), .E(n695), .CK(clk), .Q(
        \registers[405][5] ) );
  EDFFX1 \registers_reg[405][4]  ( .D(n8247), .E(n695), .CK(clk), .Q(
        \registers[405][4] ) );
  EDFFX1 \registers_reg[405][3]  ( .D(n8195), .E(n695), .CK(clk), .Q(
        \registers[405][3] ) );
  EDFFX1 \registers_reg[405][2]  ( .D(n8150), .E(n695), .CK(clk), .Q(
        \registers[405][2] ) );
  EDFFX1 \registers_reg[405][1]  ( .D(n8094), .E(n695), .CK(clk), .Q(
        \registers[405][1] ) );
  EDFFX1 \registers_reg[405][0]  ( .D(n8036), .E(n695), .CK(clk), .Q(
        \registers[405][0] ) );
  EDFFX1 \registers_reg[401][7]  ( .D(n8419), .E(n691), .CK(clk), .Q(
        \registers[401][7] ) );
  EDFFX1 \registers_reg[401][6]  ( .D(n8361), .E(n691), .CK(clk), .Q(
        \registers[401][6] ) );
  EDFFX1 \registers_reg[401][5]  ( .D(n8303), .E(n691), .CK(clk), .Q(
        \registers[401][5] ) );
  EDFFX1 \registers_reg[401][4]  ( .D(n8245), .E(n691), .CK(clk), .Q(
        \registers[401][4] ) );
  EDFFX1 \registers_reg[401][3]  ( .D(n8196), .E(n691), .CK(clk), .Q(
        \registers[401][3] ) );
  EDFFX1 \registers_reg[401][2]  ( .D(n8151), .E(n691), .CK(clk), .Q(
        \registers[401][2] ) );
  EDFFX1 \registers_reg[401][1]  ( .D(n8095), .E(n691), .CK(clk), .Q(
        \registers[401][1] ) );
  EDFFX1 \registers_reg[401][0]  ( .D(n8034), .E(n691), .CK(clk), .Q(
        \registers[401][0] ) );
  EDFFX1 \registers_reg[397][7]  ( .D(n8420), .E(n687), .CK(clk), .Q(
        \registers[397][7] ) );
  EDFFX1 \registers_reg[397][6]  ( .D(n8362), .E(n687), .CK(clk), .Q(
        \registers[397][6] ) );
  EDFFX1 \registers_reg[397][5]  ( .D(n8304), .E(n687), .CK(clk), .Q(
        \registers[397][5] ) );
  EDFFX1 \registers_reg[397][4]  ( .D(n8246), .E(n687), .CK(clk), .Q(
        \registers[397][4] ) );
  EDFFX1 \registers_reg[397][3]  ( .D(n8194), .E(n687), .CK(clk), .Q(
        \registers[397][3] ) );
  EDFFX1 \registers_reg[397][2]  ( .D(n8727), .E(n687), .CK(clk), .Q(
        \registers[397][2] ) );
  EDFFX1 \registers_reg[397][1]  ( .D(n8699), .E(n687), .CK(clk), .Q(
        \registers[397][1] ) );
  EDFFX1 \registers_reg[397][0]  ( .D(n8035), .E(n687), .CK(clk), .Q(
        \registers[397][0] ) );
  EDFFX1 \registers_reg[393][7]  ( .D(n8421), .E(n683), .CK(clk), .Q(
        \registers[393][7] ) );
  EDFFX1 \registers_reg[393][6]  ( .D(n8363), .E(n683), .CK(clk), .Q(
        \registers[393][6] ) );
  EDFFX1 \registers_reg[393][5]  ( .D(n8305), .E(n683), .CK(clk), .Q(
        \registers[393][5] ) );
  EDFFX1 \registers_reg[393][4]  ( .D(n8247), .E(n683), .CK(clk), .Q(
        \registers[393][4] ) );
  EDFFX1 \registers_reg[393][3]  ( .D(n8195), .E(n683), .CK(clk), .Q(
        \registers[393][3] ) );
  EDFFX1 \registers_reg[393][2]  ( .D(n8150), .E(n683), .CK(clk), .Q(
        \registers[393][2] ) );
  EDFFX1 \registers_reg[393][1]  ( .D(n8094), .E(n683), .CK(clk), .Q(
        \registers[393][1] ) );
  EDFFX1 \registers_reg[393][0]  ( .D(n8036), .E(n683), .CK(clk), .Q(
        \registers[393][0] ) );
  EDFFX1 \registers_reg[389][7]  ( .D(n8419), .E(n999), .CK(clk), .Q(
        \registers[389][7] ) );
  EDFFX1 \registers_reg[389][6]  ( .D(n8361), .E(n999), .CK(clk), .Q(
        \registers[389][6] ) );
  EDFFX1 \registers_reg[389][5]  ( .D(n8303), .E(n999), .CK(clk), .Q(
        \registers[389][5] ) );
  EDFFX1 \registers_reg[389][4]  ( .D(n8245), .E(n999), .CK(clk), .Q(
        \registers[389][4] ) );
  EDFFX1 \registers_reg[389][3]  ( .D(n8196), .E(n999), .CK(clk), .Q(
        \registers[389][3] ) );
  EDFFX1 \registers_reg[389][2]  ( .D(n8151), .E(n999), .CK(clk), .Q(
        \registers[389][2] ) );
  EDFFX1 \registers_reg[389][1]  ( .D(n8095), .E(n999), .CK(clk), .Q(
        \registers[389][1] ) );
  EDFFX1 \registers_reg[389][0]  ( .D(n8034), .E(n999), .CK(clk), .Q(
        \registers[389][0] ) );
  EDFFX1 \registers_reg[385][7]  ( .D(n8420), .E(n995), .CK(clk), .Q(
        \registers[385][7] ) );
  EDFFX1 \registers_reg[385][6]  ( .D(n8362), .E(n995), .CK(clk), .Q(
        \registers[385][6] ) );
  EDFFX1 \registers_reg[385][5]  ( .D(n8304), .E(n995), .CK(clk), .Q(
        \registers[385][5] ) );
  EDFFX1 \registers_reg[385][4]  ( .D(n8246), .E(n995), .CK(clk), .Q(
        \registers[385][4] ) );
  EDFFX1 \registers_reg[385][3]  ( .D(n8194), .E(n995), .CK(clk), .Q(
        \registers[385][3] ) );
  EDFFX1 \registers_reg[385][2]  ( .D(n8744), .E(n995), .CK(clk), .Q(
        \registers[385][2] ) );
  EDFFX1 \registers_reg[385][1]  ( .D(n8716), .E(n995), .CK(clk), .Q(
        \registers[385][1] ) );
  EDFFX1 \registers_reg[385][0]  ( .D(n8035), .E(n995), .CK(clk), .Q(
        \registers[385][0] ) );
  EDFFX1 \registers_reg[381][7]  ( .D(n8412), .E(n679), .CK(clk), .Q(
        \registers[381][7] ) );
  EDFFX1 \registers_reg[381][6]  ( .D(n8354), .E(n679), .CK(clk), .Q(
        \registers[381][6] ) );
  EDFFX1 \registers_reg[381][5]  ( .D(n8296), .E(n679), .CK(clk), .Q(
        \registers[381][5] ) );
  EDFFX1 \registers_reg[381][4]  ( .D(n8238), .E(n679), .CK(clk), .Q(
        \registers[381][4] ) );
  EDFFX1 \registers_reg[381][3]  ( .D(n8199), .E(n679), .CK(clk), .Q(
        \registers[381][3] ) );
  EDFFX1 \registers_reg[381][2]  ( .D(n8116), .E(n679), .CK(clk), .Q(
        \registers[381][2] ) );
  EDFFX1 \registers_reg[381][1]  ( .D(n8060), .E(n679), .CK(clk), .Q(
        \registers[381][1] ) );
  EDFFX1 \registers_reg[381][0]  ( .D(n7996), .E(n679), .CK(clk), .Q(
        \registers[381][0] ) );
  EDFFX1 \registers_reg[377][7]  ( .D(n8433), .E(n675), .CK(clk), .Q(
        \registers[377][7] ) );
  EDFFX1 \registers_reg[377][6]  ( .D(n8375), .E(n675), .CK(clk), .Q(
        \registers[377][6] ) );
  EDFFX1 \registers_reg[377][5]  ( .D(n8317), .E(n675), .CK(clk), .Q(
        \registers[377][5] ) );
  EDFFX1 \registers_reg[377][4]  ( .D(n8259), .E(n675), .CK(clk), .Q(
        \registers[377][4] ) );
  EDFFX1 \registers_reg[377][3]  ( .D(n8194), .E(n675), .CK(clk), .Q(
        \registers[377][3] ) );
  EDFFX1 \registers_reg[377][2]  ( .D(n8145), .E(n675), .CK(clk), .Q(
        \registers[377][2] ) );
  EDFFX1 \registers_reg[377][1]  ( .D(n8089), .E(n675), .CK(clk), .Q(
        \registers[377][1] ) );
  EDFFX1 \registers_reg[377][0]  ( .D(n7997), .E(n675), .CK(clk), .Q(
        \registers[377][0] ) );
  EDFFX1 \registers_reg[373][7]  ( .D(n8434), .E(n671), .CK(clk), .Q(
        \registers[373][7] ) );
  EDFFX1 \registers_reg[373][6]  ( .D(n8376), .E(n671), .CK(clk), .Q(
        \registers[373][6] ) );
  EDFFX1 \registers_reg[373][5]  ( .D(n8318), .E(n671), .CK(clk), .Q(
        \registers[373][5] ) );
  EDFFX1 \registers_reg[373][4]  ( .D(n8260), .E(n671), .CK(clk), .Q(
        \registers[373][4] ) );
  EDFFX1 \registers_reg[373][3]  ( .D(n8195), .E(n671), .CK(clk), .Q(
        \registers[373][3] ) );
  EDFFX1 \registers_reg[373][2]  ( .D(n8151), .E(n671), .CK(clk), .Q(
        \registers[373][2] ) );
  EDFFX1 \registers_reg[373][1]  ( .D(n8095), .E(n671), .CK(clk), .Q(
        \registers[373][1] ) );
  EDFFX1 \registers_reg[373][0]  ( .D(n8688), .E(n671), .CK(clk), .Q(
        \registers[373][0] ) );
  EDFFX1 \registers_reg[369][7]  ( .D(n8406), .E(n667), .CK(clk), .Q(
        \registers[369][7] ) );
  EDFFX1 \registers_reg[369][6]  ( .D(n8348), .E(n667), .CK(clk), .Q(
        \registers[369][6] ) );
  EDFFX1 \registers_reg[369][5]  ( .D(n8290), .E(n667), .CK(clk), .Q(
        \registers[369][5] ) );
  EDFFX1 \registers_reg[369][4]  ( .D(n8232), .E(n667), .CK(clk), .Q(
        \registers[369][4] ) );
  EDFFX1 \registers_reg[369][3]  ( .D(n8196), .E(n667), .CK(clk), .Q(
        \registers[369][3] ) );
  EDFFX1 \registers_reg[369][2]  ( .D(n8725), .E(n667), .CK(clk), .Q(
        \registers[369][2] ) );
  EDFFX1 \registers_reg[369][1]  ( .D(n8697), .E(n667), .CK(clk), .Q(
        \registers[369][1] ) );
  EDFFX1 \registers_reg[369][0]  ( .D(n8047), .E(n667), .CK(clk), .Q(
        \registers[369][0] ) );
  EDFFX1 \registers_reg[365][7]  ( .D(n8433), .E(n663), .CK(clk), .Q(
        \registers[365][7] ) );
  EDFFX1 \registers_reg[365][6]  ( .D(n8375), .E(n663), .CK(clk), .Q(
        \registers[365][6] ) );
  EDFFX1 \registers_reg[365][5]  ( .D(n8317), .E(n663), .CK(clk), .Q(
        \registers[365][5] ) );
  EDFFX1 \registers_reg[365][4]  ( .D(n8259), .E(n663), .CK(clk), .Q(
        \registers[365][4] ) );
  EDFFX1 \registers_reg[365][3]  ( .D(n8191), .E(n663), .CK(clk), .Q(
        \registers[365][3] ) );
  EDFFX1 \registers_reg[365][2]  ( .D(n8136), .E(n663), .CK(clk), .Q(
        \registers[365][2] ) );
  EDFFX1 \registers_reg[365][1]  ( .D(n8080), .E(n663), .CK(clk), .Q(
        \registers[365][1] ) );
  EDFFX1 \registers_reg[365][0]  ( .D(n8048), .E(n663), .CK(clk), .Q(
        \registers[365][0] ) );
  EDFFX1 \registers_reg[361][7]  ( .D(n8434), .E(n659), .CK(clk), .Q(
        \registers[361][7] ) );
  EDFFX1 \registers_reg[361][6]  ( .D(n8376), .E(n659), .CK(clk), .Q(
        \registers[361][6] ) );
  EDFFX1 \registers_reg[361][5]  ( .D(n8318), .E(n659), .CK(clk), .Q(
        \registers[361][5] ) );
  EDFFX1 \registers_reg[361][4]  ( .D(n8260), .E(n659), .CK(clk), .Q(
        \registers[361][4] ) );
  EDFFX1 \registers_reg[361][3]  ( .D(n8192), .E(n659), .CK(clk), .Q(
        \registers[361][3] ) );
  EDFFX1 \registers_reg[361][2]  ( .D(n8723), .E(n659), .CK(clk), .Q(
        \registers[361][2] ) );
  EDFFX1 \registers_reg[361][1]  ( .D(n8695), .E(n659), .CK(clk), .Q(
        \registers[361][1] ) );
  EDFFX1 \registers_reg[361][0]  ( .D(n8046), .E(n659), .CK(clk), .Q(
        \registers[361][0] ) );
  EDFFX1 \registers_reg[357][7]  ( .D(n8403), .E(n992), .CK(clk), .Q(
        \registers[357][7] ) );
  EDFFX1 \registers_reg[357][6]  ( .D(n8345), .E(n992), .CK(clk), .Q(
        \registers[357][6] ) );
  EDFFX1 \registers_reg[357][5]  ( .D(n8287), .E(n992), .CK(clk), .Q(
        \registers[357][5] ) );
  EDFFX1 \registers_reg[357][4]  ( .D(n8229), .E(n992), .CK(clk), .Q(
        \registers[357][4] ) );
  EDFFX1 \registers_reg[357][3]  ( .D(n8188), .E(n992), .CK(clk), .Q(
        \registers[357][3] ) );
  EDFFX1 \registers_reg[357][2]  ( .D(n8126), .E(n992), .CK(clk), .Q(
        \registers[357][2] ) );
  EDFFX1 \registers_reg[357][1]  ( .D(n8070), .E(n992), .CK(clk), .Q(
        \registers[357][1] ) );
  EDFFX1 \registers_reg[357][0]  ( .D(n8047), .E(n992), .CK(clk), .Q(
        \registers[357][0] ) );
  EDFFX1 \registers_reg[353][7]  ( .D(n8433), .E(n988), .CK(clk), .Q(
        \registers[353][7] ) );
  EDFFX1 \registers_reg[353][6]  ( .D(n8375), .E(n988), .CK(clk), .Q(
        \registers[353][6] ) );
  EDFFX1 \registers_reg[353][5]  ( .D(n8317), .E(n988), .CK(clk), .Q(
        \registers[353][5] ) );
  EDFFX1 \registers_reg[353][4]  ( .D(n8259), .E(n988), .CK(clk), .Q(
        \registers[353][4] ) );
  EDFFX1 \registers_reg[353][3]  ( .D(n8162), .E(n988), .CK(clk), .Q(
        \registers[353][3] ) );
  EDFFX1 \registers_reg[353][2]  ( .D(n8137), .E(n988), .CK(clk), .Q(
        \registers[353][2] ) );
  EDFFX1 \registers_reg[353][1]  ( .D(n8081), .E(n988), .CK(clk), .Q(
        \registers[353][1] ) );
  EDFFX1 \registers_reg[353][0]  ( .D(n8048), .E(n988), .CK(clk), .Q(
        \registers[353][0] ) );
  EDFFX1 \registers_reg[349][7]  ( .D(n8432), .E(n655), .CK(clk), .Q(
        \registers[349][7] ) );
  EDFFX1 \registers_reg[349][6]  ( .D(n8374), .E(n655), .CK(clk), .Q(
        \registers[349][6] ) );
  EDFFX1 \registers_reg[349][5]  ( .D(n8316), .E(n655), .CK(clk), .Q(
        \registers[349][5] ) );
  EDFFX1 \registers_reg[349][4]  ( .D(n8258), .E(n655), .CK(clk), .Q(
        \registers[349][4] ) );
  EDFFX1 \registers_reg[349][3]  ( .D(n8163), .E(n655), .CK(clk), .Q(
        \registers[349][3] ) );
  EDFFX1 \registers_reg[349][2]  ( .D(n8730), .E(n655), .CK(clk), .Q(
        \registers[349][2] ) );
  EDFFX1 \registers_reg[349][1]  ( .D(n8702), .E(n655), .CK(clk), .Q(
        \registers[349][1] ) );
  EDFFX1 \registers_reg[349][0]  ( .D(n8046), .E(n655), .CK(clk), .Q(
        \registers[349][0] ) );
  EDFFX1 \registers_reg[345][7]  ( .D(n8430), .E(n651), .CK(clk), .Q(
        \registers[345][7] ) );
  EDFFX1 \registers_reg[345][6]  ( .D(n8372), .E(n651), .CK(clk), .Q(
        \registers[345][6] ) );
  EDFFX1 \registers_reg[345][5]  ( .D(n8314), .E(n651), .CK(clk), .Q(
        \registers[345][5] ) );
  EDFFX1 \registers_reg[345][4]  ( .D(n8256), .E(n651), .CK(clk), .Q(
        \registers[345][4] ) );
  EDFFX1 \registers_reg[345][3]  ( .D(n8189), .E(n651), .CK(clk), .Q(
        \registers[345][3] ) );
  EDFFX1 \registers_reg[345][2]  ( .D(n8127), .E(n651), .CK(clk), .Q(
        \registers[345][2] ) );
  EDFFX1 \registers_reg[345][1]  ( .D(n8071), .E(n651), .CK(clk), .Q(
        \registers[345][1] ) );
  EDFFX1 \registers_reg[345][0]  ( .D(n8047), .E(n651), .CK(clk), .Q(
        \registers[345][0] ) );
  EDFFX1 \registers_reg[341][7]  ( .D(n8431), .E(n647), .CK(clk), .Q(
        \registers[341][7] ) );
  EDFFX1 \registers_reg[341][6]  ( .D(n8373), .E(n647), .CK(clk), .Q(
        \registers[341][6] ) );
  EDFFX1 \registers_reg[341][5]  ( .D(n8315), .E(n647), .CK(clk), .Q(
        \registers[341][5] ) );
  EDFFX1 \registers_reg[341][4]  ( .D(n8257), .E(n647), .CK(clk), .Q(
        \registers[341][4] ) );
  EDFFX1 \registers_reg[341][3]  ( .D(n8163), .E(n647), .CK(clk), .Q(
        \registers[341][3] ) );
  EDFFX1 \registers_reg[341][2]  ( .D(n8135), .E(n647), .CK(clk), .Q(
        \registers[341][2] ) );
  EDFFX1 \registers_reg[341][1]  ( .D(n8079), .E(n647), .CK(clk), .Q(
        \registers[341][1] ) );
  EDFFX1 \registers_reg[341][0]  ( .D(n8048), .E(n647), .CK(clk), .Q(
        \registers[341][0] ) );
  EDFFX1 \registers_reg[337][7]  ( .D(n8432), .E(n643), .CK(clk), .Q(
        \registers[337][7] ) );
  EDFFX1 \registers_reg[337][6]  ( .D(n8374), .E(n643), .CK(clk), .Q(
        \registers[337][6] ) );
  EDFFX1 \registers_reg[337][5]  ( .D(n8316), .E(n643), .CK(clk), .Q(
        \registers[337][5] ) );
  EDFFX1 \registers_reg[337][4]  ( .D(n8258), .E(n643), .CK(clk), .Q(
        \registers[337][4] ) );
  EDFFX1 \registers_reg[337][3]  ( .D(n8163), .E(n643), .CK(clk), .Q(
        \registers[337][3] ) );
  EDFFX1 \registers_reg[337][2]  ( .D(n8744), .E(n643), .CK(clk), .Q(
        \registers[337][2] ) );
  EDFFX1 \registers_reg[337][1]  ( .D(n8716), .E(n643), .CK(clk), .Q(
        \registers[337][1] ) );
  EDFFX1 \registers_reg[337][0]  ( .D(n8046), .E(n643), .CK(clk), .Q(
        \registers[337][0] ) );
  EDFFX1 \registers_reg[333][7]  ( .D(n8430), .E(n639), .CK(clk), .Q(
        \registers[333][7] ) );
  EDFFX1 \registers_reg[333][6]  ( .D(n8372), .E(n639), .CK(clk), .Q(
        \registers[333][6] ) );
  EDFFX1 \registers_reg[333][5]  ( .D(n8314), .E(n639), .CK(clk), .Q(
        \registers[333][5] ) );
  EDFFX1 \registers_reg[333][4]  ( .D(n8256), .E(n639), .CK(clk), .Q(
        \registers[333][4] ) );
  EDFFX1 \registers_reg[333][3]  ( .D(n8190), .E(n639), .CK(clk), .Q(
        \registers[333][3] ) );
  EDFFX1 \registers_reg[333][2]  ( .D(n8128), .E(n639), .CK(clk), .Q(
        \registers[333][2] ) );
  EDFFX1 \registers_reg[333][1]  ( .D(n8072), .E(n639), .CK(clk), .Q(
        \registers[333][1] ) );
  EDFFX1 \registers_reg[333][0]  ( .D(n8047), .E(n639), .CK(clk), .Q(
        \registers[333][0] ) );
  EDFFX1 \registers_reg[329][7]  ( .D(n8431), .E(n635), .CK(clk), .Q(
        \registers[329][7] ) );
  EDFFX1 \registers_reg[329][6]  ( .D(n8373), .E(n635), .CK(clk), .Q(
        \registers[329][6] ) );
  EDFFX1 \registers_reg[329][5]  ( .D(n8315), .E(n635), .CK(clk), .Q(
        \registers[329][5] ) );
  EDFFX1 \registers_reg[329][4]  ( .D(n8257), .E(n635), .CK(clk), .Q(
        \registers[329][4] ) );
  EDFFX1 \registers_reg[329][3]  ( .D(n8165), .E(n635), .CK(clk), .Q(
        \registers[329][3] ) );
  EDFFX1 \registers_reg[329][2]  ( .D(n8132), .E(n635), .CK(clk), .Q(
        \registers[329][2] ) );
  EDFFX1 \registers_reg[329][1]  ( .D(n8076), .E(n635), .CK(clk), .Q(
        \registers[329][1] ) );
  EDFFX1 \registers_reg[329][0]  ( .D(n8048), .E(n635), .CK(clk), .Q(
        \registers[329][0] ) );
  EDFFX1 \registers_reg[325][7]  ( .D(n8432), .E(n985), .CK(clk), .Q(
        \registers[325][7] ) );
  EDFFX1 \registers_reg[325][6]  ( .D(n8374), .E(n985), .CK(clk), .Q(
        \registers[325][6] ) );
  EDFFX1 \registers_reg[325][5]  ( .D(n8316), .E(n985), .CK(clk), .Q(
        \registers[325][5] ) );
  EDFFX1 \registers_reg[325][4]  ( .D(n8258), .E(n985), .CK(clk), .Q(
        \registers[325][4] ) );
  EDFFX1 \registers_reg[325][3]  ( .D(n8170), .E(n985), .CK(clk), .Q(
        \registers[325][3] ) );
  EDFFX1 \registers_reg[325][2]  ( .D(n8744), .E(n985), .CK(clk), .Q(
        \registers[325][2] ) );
  EDFFX1 \registers_reg[325][1]  ( .D(n8716), .E(n985), .CK(clk), .Q(
        \registers[325][1] ) );
  EDFFX1 \registers_reg[325][0]  ( .D(n8046), .E(n985), .CK(clk), .Q(
        \registers[325][0] ) );
  EDFFX1 \registers_reg[321][7]  ( .D(n8430), .E(n981), .CK(clk), .Q(
        \registers[321][7] ) );
  EDFFX1 \registers_reg[321][6]  ( .D(n8372), .E(n981), .CK(clk), .Q(
        \registers[321][6] ) );
  EDFFX1 \registers_reg[321][5]  ( .D(n8314), .E(n981), .CK(clk), .Q(
        \registers[321][5] ) );
  EDFFX1 \registers_reg[321][4]  ( .D(n8256), .E(n981), .CK(clk), .Q(
        \registers[321][4] ) );
  EDFFX1 \registers_reg[321][3]  ( .D(n8185), .E(n981), .CK(clk), .Q(
        \registers[321][3] ) );
  EDFFX1 \registers_reg[321][2]  ( .D(n8129), .E(n981), .CK(clk), .Q(
        \registers[321][2] ) );
  EDFFX1 \registers_reg[321][1]  ( .D(n8073), .E(n981), .CK(clk), .Q(
        \registers[321][1] ) );
  EDFFX1 \registers_reg[321][0]  ( .D(n8047), .E(n981), .CK(clk), .Q(
        \registers[321][0] ) );
  EDFFX1 \registers_reg[317][7]  ( .D(n8432), .E(n631), .CK(clk), .Q(
        \registers[317][7] ) );
  EDFFX1 \registers_reg[317][6]  ( .D(n8374), .E(n631), .CK(clk), .Q(
        \registers[317][6] ) );
  EDFFX1 \registers_reg[317][5]  ( .D(n8316), .E(n631), .CK(clk), .Q(
        \registers[317][5] ) );
  EDFFX1 \registers_reg[317][4]  ( .D(n8258), .E(n631), .CK(clk), .Q(
        \registers[317][4] ) );
  EDFFX1 \registers_reg[317][3]  ( .D(n8171), .E(n631), .CK(clk), .Q(
        \registers[317][3] ) );
  EDFFX1 \registers_reg[317][2]  ( .D(n8159), .E(n631), .CK(clk), .Q(
        \registers[317][2] ) );
  EDFFX1 \registers_reg[317][1]  ( .D(n8103), .E(n631), .CK(clk), .Q(
        \registers[317][1] ) );
  EDFFX1 \registers_reg[317][0]  ( .D(n8043), .E(n631), .CK(clk), .Q(
        \registers[317][0] ) );
  EDFFX1 \registers_reg[313][7]  ( .D(n8430), .E(n627), .CK(clk), .Q(
        \registers[313][7] ) );
  EDFFX1 \registers_reg[313][6]  ( .D(n8372), .E(n627), .CK(clk), .Q(
        \registers[313][6] ) );
  EDFFX1 \registers_reg[313][5]  ( .D(n8314), .E(n627), .CK(clk), .Q(
        \registers[313][5] ) );
  EDFFX1 \registers_reg[313][4]  ( .D(n8256), .E(n627), .CK(clk), .Q(
        \registers[313][4] ) );
  EDFFX1 \registers_reg[313][3]  ( .D(n8186), .E(n627), .CK(clk), .Q(
        \registers[313][3] ) );
  EDFFX1 \registers_reg[313][2]  ( .D(n8160), .E(n627), .CK(clk), .Q(
        \registers[313][2] ) );
  EDFFX1 \registers_reg[313][1]  ( .D(n8104), .E(n627), .CK(clk), .Q(
        \registers[313][1] ) );
  EDFFX1 \registers_reg[313][0]  ( .D(n8044), .E(n627), .CK(clk), .Q(
        \registers[313][0] ) );
  EDFFX1 \registers_reg[309][7]  ( .D(n8431), .E(n623), .CK(clk), .Q(
        \registers[309][7] ) );
  EDFFX1 \registers_reg[309][6]  ( .D(n8373), .E(n623), .CK(clk), .Q(
        \registers[309][6] ) );
  EDFFX1 \registers_reg[309][5]  ( .D(n8315), .E(n623), .CK(clk), .Q(
        \registers[309][5] ) );
  EDFFX1 \registers_reg[309][4]  ( .D(n8257), .E(n623), .CK(clk), .Q(
        \registers[309][4] ) );
  EDFFX1 \registers_reg[309][3]  ( .D(n8199), .E(n623), .CK(clk), .Q(
        \registers[309][3] ) );
  EDFFX1 \registers_reg[309][2]  ( .D(n8158), .E(n623), .CK(clk), .Q(
        \registers[309][2] ) );
  EDFFX1 \registers_reg[309][1]  ( .D(n8102), .E(n623), .CK(clk), .Q(
        \registers[309][1] ) );
  EDFFX1 \registers_reg[309][0]  ( .D(n8045), .E(n623), .CK(clk), .Q(
        \registers[309][0] ) );
  EDFFX1 \registers_reg[305][7]  ( .D(n8432), .E(n619), .CK(clk), .Q(
        \registers[305][7] ) );
  EDFFX1 \registers_reg[305][6]  ( .D(n8374), .E(n619), .CK(clk), .Q(
        \registers[305][6] ) );
  EDFFX1 \registers_reg[305][5]  ( .D(n8316), .E(n619), .CK(clk), .Q(
        \registers[305][5] ) );
  EDFFX1 \registers_reg[305][4]  ( .D(n8258), .E(n619), .CK(clk), .Q(
        \registers[305][4] ) );
  EDFFX1 \registers_reg[305][3]  ( .D(n8172), .E(n619), .CK(clk), .Q(
        \registers[305][3] ) );
  EDFFX1 \registers_reg[305][2]  ( .D(n8159), .E(n619), .CK(clk), .Q(
        \registers[305][2] ) );
  EDFFX1 \registers_reg[305][1]  ( .D(n8103), .E(n619), .CK(clk), .Q(
        \registers[305][1] ) );
  EDFFX1 \registers_reg[305][0]  ( .D(n8043), .E(n619), .CK(clk), .Q(
        \registers[305][0] ) );
  EDFFX1 \registers_reg[301][7]  ( .D(n8429), .E(n615), .CK(clk), .Q(
        \registers[301][7] ) );
  EDFFX1 \registers_reg[301][6]  ( .D(n8371), .E(n615), .CK(clk), .Q(
        \registers[301][6] ) );
  EDFFX1 \registers_reg[301][5]  ( .D(n8313), .E(n615), .CK(clk), .Q(
        \registers[301][5] ) );
  EDFFX1 \registers_reg[301][4]  ( .D(n8255), .E(n615), .CK(clk), .Q(
        \registers[301][4] ) );
  EDFFX1 \registers_reg[301][3]  ( .D(n8187), .E(n615), .CK(clk), .Q(
        \registers[301][3] ) );
  EDFFX1 \registers_reg[301][2]  ( .D(n8160), .E(n615), .CK(clk), .Q(
        \registers[301][2] ) );
  EDFFX1 \registers_reg[301][1]  ( .D(n8104), .E(n615), .CK(clk), .Q(
        \registers[301][1] ) );
  EDFFX1 \registers_reg[301][0]  ( .D(n8044), .E(n615), .CK(clk), .Q(
        \registers[301][0] ) );
  EDFFX1 \registers_reg[297][7]  ( .D(n8403), .E(n611), .CK(clk), .Q(
        \registers[297][7] ) );
  EDFFX1 \registers_reg[297][6]  ( .D(n8345), .E(n611), .CK(clk), .Q(
        \registers[297][6] ) );
  EDFFX1 \registers_reg[297][5]  ( .D(n8287), .E(n611), .CK(clk), .Q(
        \registers[297][5] ) );
  EDFFX1 \registers_reg[297][4]  ( .D(n8229), .E(n611), .CK(clk), .Q(
        \registers[297][4] ) );
  EDFFX1 \registers_reg[297][3]  ( .D(n8194), .E(n611), .CK(clk), .Q(
        \registers[297][3] ) );
  EDFFX1 \registers_reg[297][2]  ( .D(n8158), .E(n611), .CK(clk), .Q(
        \registers[297][2] ) );
  EDFFX1 \registers_reg[297][1]  ( .D(n8102), .E(n611), .CK(clk), .Q(
        \registers[297][1] ) );
  EDFFX1 \registers_reg[297][0]  ( .D(n8045), .E(n611), .CK(clk), .Q(
        \registers[297][0] ) );
  EDFFX1 \registers_reg[293][7]  ( .D(n8428), .E(n978), .CK(clk), .Q(
        \registers[293][7] ) );
  EDFFX1 \registers_reg[293][6]  ( .D(n8370), .E(n978), .CK(clk), .Q(
        \registers[293][6] ) );
  EDFFX1 \registers_reg[293][5]  ( .D(n8312), .E(n978), .CK(clk), .Q(
        \registers[293][5] ) );
  EDFFX1 \registers_reg[293][4]  ( .D(n8254), .E(n978), .CK(clk), .Q(
        \registers[293][4] ) );
  EDFFX1 \registers_reg[293][3]  ( .D(n8202), .E(n978), .CK(clk), .Q(
        \registers[293][3] ) );
  EDFFX1 \registers_reg[293][2]  ( .D(n8159), .E(n978), .CK(clk), .Q(
        \registers[293][2] ) );
  EDFFX1 \registers_reg[293][1]  ( .D(n8103), .E(n978), .CK(clk), .Q(
        \registers[293][1] ) );
  EDFFX1 \registers_reg[293][0]  ( .D(n8043), .E(n978), .CK(clk), .Q(
        \registers[293][0] ) );
  EDFFX1 \registers_reg[289][7]  ( .D(n8429), .E(n974), .CK(clk), .Q(
        \registers[289][7] ) );
  EDFFX1 \registers_reg[289][6]  ( .D(n8371), .E(n974), .CK(clk), .Q(
        \registers[289][6] ) );
  EDFFX1 \registers_reg[289][5]  ( .D(n8313), .E(n974), .CK(clk), .Q(
        \registers[289][5] ) );
  EDFFX1 \registers_reg[289][4]  ( .D(n8255), .E(n974), .CK(clk), .Q(
        \registers[289][4] ) );
  EDFFX1 \registers_reg[289][3]  ( .D(n8200), .E(n974), .CK(clk), .Q(
        \registers[289][3] ) );
  EDFFX1 \registers_reg[289][2]  ( .D(n8160), .E(n974), .CK(clk), .Q(
        \registers[289][2] ) );
  EDFFX1 \registers_reg[289][1]  ( .D(n8104), .E(n974), .CK(clk), .Q(
        \registers[289][1] ) );
  EDFFX1 \registers_reg[289][0]  ( .D(n8044), .E(n974), .CK(clk), .Q(
        \registers[289][0] ) );
  EDFFX1 \registers_reg[285][7]  ( .D(n8401), .E(n607), .CK(clk), .Q(
        \registers[285][7] ) );
  EDFFX1 \registers_reg[285][6]  ( .D(n8343), .E(n607), .CK(clk), .Q(
        \registers[285][6] ) );
  EDFFX1 \registers_reg[285][5]  ( .D(n8285), .E(n607), .CK(clk), .Q(
        \registers[285][5] ) );
  EDFFX1 \registers_reg[285][4]  ( .D(n8227), .E(n607), .CK(clk), .Q(
        \registers[285][4] ) );
  EDFFX1 \registers_reg[285][3]  ( .D(n8201), .E(n607), .CK(clk), .Q(
        \registers[285][3] ) );
  EDFFX1 \registers_reg[285][2]  ( .D(n8158), .E(n607), .CK(clk), .Q(
        \registers[285][2] ) );
  EDFFX1 \registers_reg[285][1]  ( .D(n8102), .E(n607), .CK(clk), .Q(
        \registers[285][1] ) );
  EDFFX1 \registers_reg[285][0]  ( .D(n8045), .E(n607), .CK(clk), .Q(
        \registers[285][0] ) );
  EDFFX1 \registers_reg[281][7]  ( .D(n8428), .E(n603), .CK(clk), .Q(
        \registers[281][7] ) );
  EDFFX1 \registers_reg[281][6]  ( .D(n8370), .E(n603), .CK(clk), .Q(
        \registers[281][6] ) );
  EDFFX1 \registers_reg[281][5]  ( .D(n8312), .E(n603), .CK(clk), .Q(
        \registers[281][5] ) );
  EDFFX1 \registers_reg[281][4]  ( .D(n8254), .E(n603), .CK(clk), .Q(
        \registers[281][4] ) );
  EDFFX1 \registers_reg[281][3]  ( .D(n8202), .E(n603), .CK(clk), .Q(
        \registers[281][3] ) );
  EDFFX1 \registers_reg[281][2]  ( .D(n8159), .E(n603), .CK(clk), .Q(
        \registers[281][2] ) );
  EDFFX1 \registers_reg[281][1]  ( .D(n8103), .E(n603), .CK(clk), .Q(
        \registers[281][1] ) );
  EDFFX1 \registers_reg[281][0]  ( .D(n8043), .E(n603), .CK(clk), .Q(
        \registers[281][0] ) );
  EDFFX1 \registers_reg[277][7]  ( .D(n8429), .E(n599), .CK(clk), .Q(
        \registers[277][7] ) );
  EDFFX1 \registers_reg[277][6]  ( .D(n8371), .E(n599), .CK(clk), .Q(
        \registers[277][6] ) );
  EDFFX1 \registers_reg[277][5]  ( .D(n8313), .E(n599), .CK(clk), .Q(
        \registers[277][5] ) );
  EDFFX1 \registers_reg[277][4]  ( .D(n8255), .E(n599), .CK(clk), .Q(
        \registers[277][4] ) );
  EDFFX1 \registers_reg[277][3]  ( .D(n8200), .E(n599), .CK(clk), .Q(
        \registers[277][3] ) );
  EDFFX1 \registers_reg[277][2]  ( .D(n8160), .E(n599), .CK(clk), .Q(
        \registers[277][2] ) );
  EDFFX1 \registers_reg[277][1]  ( .D(n8104), .E(n599), .CK(clk), .Q(
        \registers[277][1] ) );
  EDFFX1 \registers_reg[277][0]  ( .D(n8044), .E(n599), .CK(clk), .Q(
        \registers[277][0] ) );
  EDFFX1 \registers_reg[273][7]  ( .D(n8402), .E(n595), .CK(clk), .Q(
        \registers[273][7] ) );
  EDFFX1 \registers_reg[273][6]  ( .D(n8344), .E(n595), .CK(clk), .Q(
        \registers[273][6] ) );
  EDFFX1 \registers_reg[273][5]  ( .D(n8286), .E(n595), .CK(clk), .Q(
        \registers[273][5] ) );
  EDFFX1 \registers_reg[273][4]  ( .D(n8228), .E(n595), .CK(clk), .Q(
        \registers[273][4] ) );
  EDFFX1 \registers_reg[273][3]  ( .D(n8201), .E(n595), .CK(clk), .Q(
        \registers[273][3] ) );
  EDFFX1 \registers_reg[273][2]  ( .D(n8158), .E(n595), .CK(clk), .Q(
        \registers[273][2] ) );
  EDFFX1 \registers_reg[273][1]  ( .D(n8102), .E(n595), .CK(clk), .Q(
        \registers[273][1] ) );
  EDFFX1 \registers_reg[273][0]  ( .D(n8045), .E(n595), .CK(clk), .Q(
        \registers[273][0] ) );
  EDFFX1 \registers_reg[269][7]  ( .D(n8428), .E(n591), .CK(clk), .Q(
        \registers[269][7] ) );
  EDFFX1 \registers_reg[269][6]  ( .D(n8370), .E(n591), .CK(clk), .Q(
        \registers[269][6] ) );
  EDFFX1 \registers_reg[269][5]  ( .D(n8312), .E(n591), .CK(clk), .Q(
        \registers[269][5] ) );
  EDFFX1 \registers_reg[269][4]  ( .D(n8254), .E(n591), .CK(clk), .Q(
        \registers[269][4] ) );
  EDFFX1 \registers_reg[269][3]  ( .D(n8202), .E(n591), .CK(clk), .Q(
        \registers[269][3] ) );
  EDFFX1 \registers_reg[269][2]  ( .D(n8156), .E(n591), .CK(clk), .Q(
        \registers[269][2] ) );
  EDFFX1 \registers_reg[269][1]  ( .D(n8100), .E(n591), .CK(clk), .Q(
        \registers[269][1] ) );
  EDFFX1 \registers_reg[269][0]  ( .D(n8040), .E(n591), .CK(clk), .Q(
        \registers[269][0] ) );
  EDFFX1 \registers_reg[265][7]  ( .D(n8429), .E(n587), .CK(clk), .Q(
        \registers[265][7] ) );
  EDFFX1 \registers_reg[265][6]  ( .D(n8371), .E(n587), .CK(clk), .Q(
        \registers[265][6] ) );
  EDFFX1 \registers_reg[265][5]  ( .D(n8313), .E(n587), .CK(clk), .Q(
        \registers[265][5] ) );
  EDFFX1 \registers_reg[265][4]  ( .D(n8255), .E(n587), .CK(clk), .Q(
        \registers[265][4] ) );
  EDFFX1 \registers_reg[265][3]  ( .D(n8200), .E(n587), .CK(clk), .Q(
        \registers[265][3] ) );
  EDFFX1 \registers_reg[265][2]  ( .D(n8157), .E(n587), .CK(clk), .Q(
        \registers[265][2] ) );
  EDFFX1 \registers_reg[265][1]  ( .D(n8101), .E(n587), .CK(clk), .Q(
        \registers[265][1] ) );
  EDFFX1 \registers_reg[265][0]  ( .D(n8041), .E(n587), .CK(clk), .Q(
        \registers[265][0] ) );
  EDFFX1 \registers_reg[261][7]  ( .D(n8412), .E(n971), .CK(clk), .Q(
        \registers[261][7] ) );
  EDFFX1 \registers_reg[261][6]  ( .D(n8354), .E(n971), .CK(clk), .Q(
        \registers[261][6] ) );
  EDFFX1 \registers_reg[261][5]  ( .D(n8296), .E(n971), .CK(clk), .Q(
        \registers[261][5] ) );
  EDFFX1 \registers_reg[261][4]  ( .D(n8238), .E(n971), .CK(clk), .Q(
        \registers[261][4] ) );
  EDFFX1 \registers_reg[261][3]  ( .D(n8201), .E(n971), .CK(clk), .Q(
        \registers[261][3] ) );
  EDFFX1 \registers_reg[261][2]  ( .D(n8155), .E(n971), .CK(clk), .Q(
        \registers[261][2] ) );
  EDFFX1 \registers_reg[261][1]  ( .D(n8099), .E(n971), .CK(clk), .Q(
        \registers[261][1] ) );
  EDFFX1 \registers_reg[261][0]  ( .D(n8042), .E(n971), .CK(clk), .Q(
        \registers[261][0] ) );
  EDFFX1 \registers_reg[257][7]  ( .D(n8431), .E(n967), .CK(clk), .Q(
        \registers[257][7] ) );
  EDFFX1 \registers_reg[257][6]  ( .D(n8373), .E(n967), .CK(clk), .Q(
        \registers[257][6] ) );
  EDFFX1 \registers_reg[257][5]  ( .D(n8315), .E(n967), .CK(clk), .Q(
        \registers[257][5] ) );
  EDFFX1 \registers_reg[257][4]  ( .D(n8257), .E(n967), .CK(clk), .Q(
        \registers[257][4] ) );
  EDFFX1 \registers_reg[257][3]  ( .D(n8195), .E(n967), .CK(clk), .Q(
        \registers[257][3] ) );
  EDFFX1 \registers_reg[257][2]  ( .D(n8158), .E(n967), .CK(clk), .Q(
        \registers[257][2] ) );
  EDFFX1 \registers_reg[257][1]  ( .D(n8102), .E(n967), .CK(clk), .Q(
        \registers[257][1] ) );
  EDFFX1 \registers_reg[257][0]  ( .D(n8040), .E(n967), .CK(clk), .Q(
        \registers[257][0] ) );
  EDFFX1 \registers_reg[253][7]  ( .D(n8411), .E(n583), .CK(clk), .Q(
        \registers[253][7] ) );
  EDFFX1 \registers_reg[253][6]  ( .D(n8353), .E(n583), .CK(clk), .Q(
        \registers[253][6] ) );
  EDFFX1 \registers_reg[253][5]  ( .D(n8295), .E(n583), .CK(clk), .Q(
        \registers[253][5] ) );
  EDFFX1 \registers_reg[253][4]  ( .D(n8237), .E(n583), .CK(clk), .Q(
        \registers[253][4] ) );
  EDFFX1 \registers_reg[253][3]  ( .D(n8188), .E(n583), .CK(clk), .Q(
        \registers[253][3] ) );
  EDFFX1 \registers_reg[253][2]  ( .D(n8143), .E(n583), .CK(clk), .Q(
        \registers[253][2] ) );
  EDFFX1 \registers_reg[253][1]  ( .D(n8087), .E(n583), .CK(clk), .Q(
        \registers[253][1] ) );
  EDFFX1 \registers_reg[253][0]  ( .D(n8026), .E(n583), .CK(clk), .Q(
        \registers[253][0] ) );
  EDFFX1 \registers_reg[249][7]  ( .D(n8412), .E(n579), .CK(clk), .Q(
        \registers[249][7] ) );
  EDFFX1 \registers_reg[249][6]  ( .D(n8354), .E(n579), .CK(clk), .Q(
        \registers[249][6] ) );
  EDFFX1 \registers_reg[249][5]  ( .D(n8296), .E(n579), .CK(clk), .Q(
        \registers[249][5] ) );
  EDFFX1 \registers_reg[249][4]  ( .D(n8238), .E(n579), .CK(clk), .Q(
        \registers[249][4] ) );
  EDFFX1 \registers_reg[249][3]  ( .D(n8189), .E(n579), .CK(clk), .Q(
        \registers[249][3] ) );
  EDFFX1 \registers_reg[249][2]  ( .D(n8141), .E(n579), .CK(clk), .Q(
        \registers[249][2] ) );
  EDFFX1 \registers_reg[249][1]  ( .D(n8085), .E(n579), .CK(clk), .Q(
        \registers[249][1] ) );
  EDFFX1 \registers_reg[249][0]  ( .D(n8027), .E(n579), .CK(clk), .Q(
        \registers[249][0] ) );
  EDFFX1 \registers_reg[245][7]  ( .D(n8410), .E(n575), .CK(clk), .Q(
        \registers[245][7] ) );
  EDFFX1 \registers_reg[245][6]  ( .D(n8352), .E(n575), .CK(clk), .Q(
        \registers[245][6] ) );
  EDFFX1 \registers_reg[245][5]  ( .D(n8294), .E(n575), .CK(clk), .Q(
        \registers[245][5] ) );
  EDFFX1 \registers_reg[245][4]  ( .D(n8236), .E(n575), .CK(clk), .Q(
        \registers[245][4] ) );
  EDFFX1 \registers_reg[245][3]  ( .D(n8190), .E(n575), .CK(clk), .Q(
        \registers[245][3] ) );
  EDFFX1 \registers_reg[245][2]  ( .D(n8142), .E(n575), .CK(clk), .Q(
        \registers[245][2] ) );
  EDFFX1 \registers_reg[245][1]  ( .D(n8086), .E(n575), .CK(clk), .Q(
        \registers[245][1] ) );
  EDFFX1 \registers_reg[245][0]  ( .D(n8025), .E(n575), .CK(clk), .Q(
        \registers[245][0] ) );
  EDFFX1 \registers_reg[241][7]  ( .D(n8411), .E(n571), .CK(clk), .Q(
        \registers[241][7] ) );
  EDFFX1 \registers_reg[241][6]  ( .D(n8353), .E(n571), .CK(clk), .Q(
        \registers[241][6] ) );
  EDFFX1 \registers_reg[241][5]  ( .D(n8295), .E(n571), .CK(clk), .Q(
        \registers[241][5] ) );
  EDFFX1 \registers_reg[241][4]  ( .D(n8237), .E(n571), .CK(clk), .Q(
        \registers[241][4] ) );
  EDFFX1 \registers_reg[241][3]  ( .D(n8188), .E(n571), .CK(clk), .Q(
        \registers[241][3] ) );
  EDFFX1 \registers_reg[241][2]  ( .D(n8143), .E(n571), .CK(clk), .Q(
        \registers[241][2] ) );
  EDFFX1 \registers_reg[241][1]  ( .D(n8087), .E(n571), .CK(clk), .Q(
        \registers[241][1] ) );
  EDFFX1 \registers_reg[241][0]  ( .D(n8026), .E(n571), .CK(clk), .Q(
        \registers[241][0] ) );
  EDFFX1 \registers_reg[237][7]  ( .D(n8412), .E(n567), .CK(clk), .Q(
        \registers[237][7] ) );
  EDFFX1 \registers_reg[237][6]  ( .D(n8354), .E(n567), .CK(clk), .Q(
        \registers[237][6] ) );
  EDFFX1 \registers_reg[237][5]  ( .D(n8296), .E(n567), .CK(clk), .Q(
        \registers[237][5] ) );
  EDFFX1 \registers_reg[237][4]  ( .D(n8238), .E(n567), .CK(clk), .Q(
        \registers[237][4] ) );
  EDFFX1 \registers_reg[237][3]  ( .D(n8189), .E(n567), .CK(clk), .Q(
        \registers[237][3] ) );
  EDFFX1 \registers_reg[237][2]  ( .D(n8141), .E(n567), .CK(clk), .Q(
        \registers[237][2] ) );
  EDFFX1 \registers_reg[237][1]  ( .D(n8085), .E(n567), .CK(clk), .Q(
        \registers[237][1] ) );
  EDFFX1 \registers_reg[237][0]  ( .D(n8027), .E(n567), .CK(clk), .Q(
        \registers[237][0] ) );
  EDFFX1 \registers_reg[233][7]  ( .D(n8410), .E(n563), .CK(clk), .Q(
        \registers[233][7] ) );
  EDFFX1 \registers_reg[233][6]  ( .D(n8352), .E(n563), .CK(clk), .Q(
        \registers[233][6] ) );
  EDFFX1 \registers_reg[233][5]  ( .D(n8294), .E(n563), .CK(clk), .Q(
        \registers[233][5] ) );
  EDFFX1 \registers_reg[233][4]  ( .D(n8236), .E(n563), .CK(clk), .Q(
        \registers[233][4] ) );
  EDFFX1 \registers_reg[233][3]  ( .D(n8187), .E(n563), .CK(clk), .Q(
        \registers[233][3] ) );
  EDFFX1 \registers_reg[233][2]  ( .D(n8142), .E(n563), .CK(clk), .Q(
        \registers[233][2] ) );
  EDFFX1 \registers_reg[233][1]  ( .D(n8086), .E(n563), .CK(clk), .Q(
        \registers[233][1] ) );
  EDFFX1 \registers_reg[233][0]  ( .D(n8025), .E(n563), .CK(clk), .Q(
        \registers[233][0] ) );
  EDFFX1 \registers_reg[229][7]  ( .D(n8411), .E(n1031), .CK(clk), .Q(
        \registers[229][7] ) );
  EDFFX1 \registers_reg[229][6]  ( .D(n8353), .E(n1031), .CK(clk), .Q(
        \registers[229][6] ) );
  EDFFX1 \registers_reg[229][5]  ( .D(n8295), .E(n1031), .CK(clk), .Q(
        \registers[229][5] ) );
  EDFFX1 \registers_reg[229][4]  ( .D(n8237), .E(n1031), .CK(clk), .Q(
        \registers[229][4] ) );
  EDFFX1 \registers_reg[229][3]  ( .D(n8185), .E(n1031), .CK(clk), .Q(
        \registers[229][3] ) );
  EDFFX1 \registers_reg[229][2]  ( .D(n8143), .E(n1031), .CK(clk), .Q(
        \registers[229][2] ) );
  EDFFX1 \registers_reg[229][1]  ( .D(n8087), .E(n1031), .CK(clk), .Q(
        \registers[229][1] ) );
  EDFFX1 \registers_reg[229][0]  ( .D(n8026), .E(n1031), .CK(clk), .Q(
        \registers[229][0] ) );
  EDFFX1 \registers_reg[225][7]  ( .D(n8412), .E(n964), .CK(clk), .Q(
        \registers[225][7] ) );
  EDFFX1 \registers_reg[225][6]  ( .D(n8354), .E(n964), .CK(clk), .Q(
        \registers[225][6] ) );
  EDFFX1 \registers_reg[225][5]  ( .D(n8296), .E(n964), .CK(clk), .Q(
        \registers[225][5] ) );
  EDFFX1 \registers_reg[225][4]  ( .D(n8238), .E(n964), .CK(clk), .Q(
        \registers[225][4] ) );
  EDFFX1 \registers_reg[225][3]  ( .D(n8186), .E(n964), .CK(clk), .Q(
        \registers[225][3] ) );
  EDFFX1 \registers_reg[225][2]  ( .D(n8141), .E(n964), .CK(clk), .Q(
        \registers[225][2] ) );
  EDFFX1 \registers_reg[225][1]  ( .D(n8085), .E(n964), .CK(clk), .Q(
        \registers[225][1] ) );
  EDFFX1 \registers_reg[225][0]  ( .D(n8027), .E(n964), .CK(clk), .Q(
        \registers[225][0] ) );
  EDFFX1 \registers_reg[221][7]  ( .D(n8410), .E(n559), .CK(clk), .Q(
        \registers[221][7] ) );
  EDFFX1 \registers_reg[221][6]  ( .D(n8352), .E(n559), .CK(clk), .Q(
        \registers[221][6] ) );
  EDFFX1 \registers_reg[221][5]  ( .D(n8294), .E(n559), .CK(clk), .Q(
        \registers[221][5] ) );
  EDFFX1 \registers_reg[221][4]  ( .D(n8236), .E(n559), .CK(clk), .Q(
        \registers[221][4] ) );
  EDFFX1 \registers_reg[221][3]  ( .D(n8187), .E(n559), .CK(clk), .Q(
        \registers[221][3] ) );
  EDFFX1 \registers_reg[221][2]  ( .D(n8142), .E(n559), .CK(clk), .Q(
        \registers[221][2] ) );
  EDFFX1 \registers_reg[221][1]  ( .D(n8086), .E(n559), .CK(clk), .Q(
        \registers[221][1] ) );
  EDFFX1 \registers_reg[221][0]  ( .D(n8025), .E(n559), .CK(clk), .Q(
        \registers[221][0] ) );
  EDFFX1 \registers_reg[217][7]  ( .D(n8411), .E(n555), .CK(clk), .Q(
        \registers[217][7] ) );
  EDFFX1 \registers_reg[217][6]  ( .D(n8353), .E(n555), .CK(clk), .Q(
        \registers[217][6] ) );
  EDFFX1 \registers_reg[217][5]  ( .D(n8295), .E(n555), .CK(clk), .Q(
        \registers[217][5] ) );
  EDFFX1 \registers_reg[217][4]  ( .D(n8237), .E(n555), .CK(clk), .Q(
        \registers[217][4] ) );
  EDFFX1 \registers_reg[217][3]  ( .D(n8185), .E(n555), .CK(clk), .Q(
        \registers[217][3] ) );
  EDFFX1 \registers_reg[217][2]  ( .D(n8140), .E(n555), .CK(clk), .Q(
        \registers[217][2] ) );
  EDFFX1 \registers_reg[217][1]  ( .D(n8084), .E(n555), .CK(clk), .Q(
        \registers[217][1] ) );
  EDFFX1 \registers_reg[217][0]  ( .D(n8023), .E(n555), .CK(clk), .Q(
        \registers[217][0] ) );
  EDFFX1 \registers_reg[213][7]  ( .D(n8412), .E(n551), .CK(clk), .Q(
        \registers[213][7] ) );
  EDFFX1 \registers_reg[213][6]  ( .D(n8354), .E(n551), .CK(clk), .Q(
        \registers[213][6] ) );
  EDFFX1 \registers_reg[213][5]  ( .D(n8296), .E(n551), .CK(clk), .Q(
        \registers[213][5] ) );
  EDFFX1 \registers_reg[213][4]  ( .D(n8238), .E(n551), .CK(clk), .Q(
        \registers[213][4] ) );
  EDFFX1 \registers_reg[213][3]  ( .D(n8186), .E(n551), .CK(clk), .Q(
        \registers[213][3] ) );
  EDFFX1 \registers_reg[213][2]  ( .D(n8138), .E(n551), .CK(clk), .Q(
        \registers[213][2] ) );
  EDFFX1 \registers_reg[213][1]  ( .D(n8082), .E(n551), .CK(clk), .Q(
        \registers[213][1] ) );
  EDFFX1 \registers_reg[213][0]  ( .D(n8024), .E(n551), .CK(clk), .Q(
        \registers[213][0] ) );
  EDFFX1 \registers_reg[209][7]  ( .D(n8410), .E(n547), .CK(clk), .Q(
        \registers[209][7] ) );
  EDFFX1 \registers_reg[209][6]  ( .D(n8352), .E(n547), .CK(clk), .Q(
        \registers[209][6] ) );
  EDFFX1 \registers_reg[209][5]  ( .D(n8294), .E(n547), .CK(clk), .Q(
        \registers[209][5] ) );
  EDFFX1 \registers_reg[209][4]  ( .D(n8236), .E(n547), .CK(clk), .Q(
        \registers[209][4] ) );
  EDFFX1 \registers_reg[209][3]  ( .D(n8187), .E(n547), .CK(clk), .Q(
        \registers[209][3] ) );
  EDFFX1 \registers_reg[209][2]  ( .D(n8139), .E(n547), .CK(clk), .Q(
        \registers[209][2] ) );
  EDFFX1 \registers_reg[209][1]  ( .D(n8083), .E(n547), .CK(clk), .Q(
        \registers[209][1] ) );
  EDFFX1 \registers_reg[209][0]  ( .D(n8022), .E(n547), .CK(clk), .Q(
        \registers[209][0] ) );
  EDFFX1 \registers_reg[205][7]  ( .D(n8409), .E(n543), .CK(clk), .Q(
        \registers[205][7] ) );
  EDFFX1 \registers_reg[205][6]  ( .D(n8351), .E(n543), .CK(clk), .Q(
        \registers[205][6] ) );
  EDFFX1 \registers_reg[205][5]  ( .D(n8293), .E(n543), .CK(clk), .Q(
        \registers[205][5] ) );
  EDFFX1 \registers_reg[205][4]  ( .D(n8235), .E(n543), .CK(clk), .Q(
        \registers[205][4] ) );
  EDFFX1 \registers_reg[205][3]  ( .D(n8185), .E(n543), .CK(clk), .Q(
        \registers[205][3] ) );
  EDFFX1 \registers_reg[205][2]  ( .D(n8140), .E(n543), .CK(clk), .Q(
        \registers[205][2] ) );
  EDFFX1 \registers_reg[205][1]  ( .D(n8084), .E(n543), .CK(clk), .Q(
        \registers[205][1] ) );
  EDFFX1 \registers_reg[205][0]  ( .D(n8023), .E(n543), .CK(clk), .Q(
        \registers[205][0] ) );
  EDFFX1 \registers_reg[201][7]  ( .D(n8407), .E(n539), .CK(clk), .Q(
        \registers[201][7] ) );
  EDFFX1 \registers_reg[201][6]  ( .D(n8349), .E(n539), .CK(clk), .Q(
        \registers[201][6] ) );
  EDFFX1 \registers_reg[201][5]  ( .D(n8291), .E(n539), .CK(clk), .Q(
        \registers[201][5] ) );
  EDFFX1 \registers_reg[201][4]  ( .D(n8233), .E(n539), .CK(clk), .Q(
        \registers[201][4] ) );
  EDFFX1 \registers_reg[201][3]  ( .D(n8186), .E(n539), .CK(clk), .Q(
        \registers[201][3] ) );
  EDFFX1 \registers_reg[201][2]  ( .D(n8138), .E(n539), .CK(clk), .Q(
        \registers[201][2] ) );
  EDFFX1 \registers_reg[201][1]  ( .D(n8082), .E(n539), .CK(clk), .Q(
        \registers[201][1] ) );
  EDFFX1 \registers_reg[201][0]  ( .D(n8024), .E(n539), .CK(clk), .Q(
        \registers[201][0] ) );
  EDFFX1 \registers_reg[197][7]  ( .D(n8408), .E(n1027), .CK(clk), .Q(
        \registers[197][7] ) );
  EDFFX1 \registers_reg[197][6]  ( .D(n8350), .E(n1027), .CK(clk), .Q(
        \registers[197][6] ) );
  EDFFX1 \registers_reg[197][5]  ( .D(n8292), .E(n1027), .CK(clk), .Q(
        \registers[197][5] ) );
  EDFFX1 \registers_reg[197][4]  ( .D(n8234), .E(n1027), .CK(clk), .Q(
        \registers[197][4] ) );
  EDFFX1 \registers_reg[197][3]  ( .D(n8187), .E(n1027), .CK(clk), .Q(
        \registers[197][3] ) );
  EDFFX1 \registers_reg[197][2]  ( .D(n8139), .E(n1027), .CK(clk), .Q(
        \registers[197][2] ) );
  EDFFX1 \registers_reg[197][1]  ( .D(n8083), .E(n1027), .CK(clk), .Q(
        \registers[197][1] ) );
  EDFFX1 \registers_reg[197][0]  ( .D(n8022), .E(n1027), .CK(clk), .Q(
        \registers[197][0] ) );
  EDFFX1 \registers_reg[193][7]  ( .D(n8409), .E(n961), .CK(clk), .Q(
        \registers[193][7] ) );
  EDFFX1 \registers_reg[193][6]  ( .D(n8351), .E(n961), .CK(clk), .Q(
        \registers[193][6] ) );
  EDFFX1 \registers_reg[193][5]  ( .D(n8293), .E(n961), .CK(clk), .Q(
        \registers[193][5] ) );
  EDFFX1 \registers_reg[193][4]  ( .D(n8235), .E(n961), .CK(clk), .Q(
        \registers[193][4] ) );
  EDFFX1 \registers_reg[193][3]  ( .D(n8185), .E(n961), .CK(clk), .Q(
        \registers[193][3] ) );
  EDFFX1 \registers_reg[193][2]  ( .D(n8140), .E(n961), .CK(clk), .Q(
        \registers[193][2] ) );
  EDFFX1 \registers_reg[193][1]  ( .D(n8084), .E(n961), .CK(clk), .Q(
        \registers[193][1] ) );
  EDFFX1 \registers_reg[193][0]  ( .D(n8023), .E(n961), .CK(clk), .Q(
        \registers[193][0] ) );
  EDFFX1 \registers_reg[189][7]  ( .D(n8408), .E(n535), .CK(clk), .Q(
        \registers[189][7] ) );
  EDFFX1 \registers_reg[189][6]  ( .D(n8350), .E(n535), .CK(clk), .Q(
        \registers[189][6] ) );
  EDFFX1 \registers_reg[189][5]  ( .D(n8292), .E(n535), .CK(clk), .Q(
        \registers[189][5] ) );
  EDFFX1 \registers_reg[189][4]  ( .D(n8234), .E(n535), .CK(clk), .Q(
        \registers[189][4] ) );
  EDFFX1 \registers_reg[189][3]  ( .D(n8187), .E(n535), .CK(clk), .Q(
        \registers[189][3] ) );
  EDFFX1 \registers_reg[189][2]  ( .D(n8139), .E(n535), .CK(clk), .Q(
        \registers[189][2] ) );
  EDFFX1 \registers_reg[189][1]  ( .D(n8083), .E(n535), .CK(clk), .Q(
        \registers[189][1] ) );
  EDFFX1 \registers_reg[189][0]  ( .D(n8022), .E(n535), .CK(clk), .Q(
        \registers[189][0] ) );
  EDFFX1 \registers_reg[185][7]  ( .D(n8409), .E(n531), .CK(clk), .Q(
        \registers[185][7] ) );
  EDFFX1 \registers_reg[185][6]  ( .D(n8351), .E(n531), .CK(clk), .Q(
        \registers[185][6] ) );
  EDFFX1 \registers_reg[185][5]  ( .D(n8293), .E(n531), .CK(clk), .Q(
        \registers[185][5] ) );
  EDFFX1 \registers_reg[185][4]  ( .D(n8235), .E(n531), .CK(clk), .Q(
        \registers[185][4] ) );
  EDFFX1 \registers_reg[185][3]  ( .D(n8185), .E(n531), .CK(clk), .Q(
        \registers[185][3] ) );
  EDFFX1 \registers_reg[185][2]  ( .D(n8140), .E(n531), .CK(clk), .Q(
        \registers[185][2] ) );
  EDFFX1 \registers_reg[185][1]  ( .D(n8084), .E(n531), .CK(clk), .Q(
        \registers[185][1] ) );
  EDFFX1 \registers_reg[185][0]  ( .D(n8023), .E(n531), .CK(clk), .Q(
        \registers[185][0] ) );
  EDFFX1 \registers_reg[181][7]  ( .D(n8407), .E(n527), .CK(clk), .Q(
        \registers[181][7] ) );
  EDFFX1 \registers_reg[181][6]  ( .D(n8349), .E(n527), .CK(clk), .Q(
        \registers[181][6] ) );
  EDFFX1 \registers_reg[181][5]  ( .D(n8291), .E(n527), .CK(clk), .Q(
        \registers[181][5] ) );
  EDFFX1 \registers_reg[181][4]  ( .D(n8233), .E(n527), .CK(clk), .Q(
        \registers[181][4] ) );
  EDFFX1 \registers_reg[181][3]  ( .D(n8186), .E(n527), .CK(clk), .Q(
        \registers[181][3] ) );
  EDFFX1 \registers_reg[181][2]  ( .D(n8138), .E(n527), .CK(clk), .Q(
        \registers[181][2] ) );
  EDFFX1 \registers_reg[181][1]  ( .D(n8082), .E(n527), .CK(clk), .Q(
        \registers[181][1] ) );
  EDFFX1 \registers_reg[181][0]  ( .D(n8024), .E(n527), .CK(clk), .Q(
        \registers[181][0] ) );
  EDFFX1 \registers_reg[177][7]  ( .D(n8408), .E(n523), .CK(clk), .Q(
        \registers[177][7] ) );
  EDFFX1 \registers_reg[177][6]  ( .D(n8350), .E(n523), .CK(clk), .Q(
        \registers[177][6] ) );
  EDFFX1 \registers_reg[177][5]  ( .D(n8292), .E(n523), .CK(clk), .Q(
        \registers[177][5] ) );
  EDFFX1 \registers_reg[177][4]  ( .D(n8234), .E(n523), .CK(clk), .Q(
        \registers[177][4] ) );
  EDFFX1 \registers_reg[177][3]  ( .D(n8187), .E(n523), .CK(clk), .Q(
        \registers[177][3] ) );
  EDFFX1 \registers_reg[177][2]  ( .D(n8139), .E(n523), .CK(clk), .Q(
        \registers[177][2] ) );
  EDFFX1 \registers_reg[177][1]  ( .D(n8083), .E(n523), .CK(clk), .Q(
        \registers[177][1] ) );
  EDFFX1 \registers_reg[177][0]  ( .D(n8022), .E(n523), .CK(clk), .Q(
        \registers[177][0] ) );
  EDFFX1 \registers_reg[173][7]  ( .D(n8409), .E(n519), .CK(clk), .Q(
        \registers[173][7] ) );
  EDFFX1 \registers_reg[173][6]  ( .D(n8351), .E(n519), .CK(clk), .Q(
        \registers[173][6] ) );
  EDFFX1 \registers_reg[173][5]  ( .D(n8293), .E(n519), .CK(clk), .Q(
        \registers[173][5] ) );
  EDFFX1 \registers_reg[173][4]  ( .D(n8235), .E(n519), .CK(clk), .Q(
        \registers[173][4] ) );
  EDFFX1 \registers_reg[173][3]  ( .D(n8182), .E(n519), .CK(clk), .Q(
        \registers[173][3] ) );
  EDFFX1 \registers_reg[173][2]  ( .D(n8140), .E(n519), .CK(clk), .Q(
        \registers[173][2] ) );
  EDFFX1 \registers_reg[173][1]  ( .D(n8084), .E(n519), .CK(clk), .Q(
        \registers[173][1] ) );
  EDFFX1 \registers_reg[173][0]  ( .D(n8023), .E(n519), .CK(clk), .Q(
        \registers[173][0] ) );
  EDFFX1 \registers_reg[169][7]  ( .D(n8407), .E(n515), .CK(clk), .Q(
        \registers[169][7] ) );
  EDFFX1 \registers_reg[169][6]  ( .D(n8349), .E(n515), .CK(clk), .Q(
        \registers[169][6] ) );
  EDFFX1 \registers_reg[169][5]  ( .D(n8291), .E(n515), .CK(clk), .Q(
        \registers[169][5] ) );
  EDFFX1 \registers_reg[169][4]  ( .D(n8233), .E(n515), .CK(clk), .Q(
        \registers[169][4] ) );
  EDFFX1 \registers_reg[169][3]  ( .D(n8183), .E(n515), .CK(clk), .Q(
        \registers[169][3] ) );
  EDFFX1 \registers_reg[169][2]  ( .D(n8135), .E(n515), .CK(clk), .Q(
        \registers[169][2] ) );
  EDFFX1 \registers_reg[169][1]  ( .D(n8079), .E(n515), .CK(clk), .Q(
        \registers[169][1] ) );
  EDFFX1 \registers_reg[169][0]  ( .D(n8024), .E(n515), .CK(clk), .Q(
        \registers[169][0] ) );
  EDFFX1 \registers_reg[165][7]  ( .D(n8408), .E(n1023), .CK(clk), .Q(
        \registers[165][7] ) );
  EDFFX1 \registers_reg[165][6]  ( .D(n8350), .E(n1023), .CK(clk), .Q(
        \registers[165][6] ) );
  EDFFX1 \registers_reg[165][5]  ( .D(n8292), .E(n1023), .CK(clk), .Q(
        \registers[165][5] ) );
  EDFFX1 \registers_reg[165][4]  ( .D(n8234), .E(n1023), .CK(clk), .Q(
        \registers[165][4] ) );
  EDFFX1 \registers_reg[165][3]  ( .D(n8184), .E(n1023), .CK(clk), .Q(
        \registers[165][3] ) );
  EDFFX1 \registers_reg[165][2]  ( .D(n8136), .E(n1023), .CK(clk), .Q(
        \registers[165][2] ) );
  EDFFX1 \registers_reg[165][1]  ( .D(n8080), .E(n1023), .CK(clk), .Q(
        \registers[165][1] ) );
  EDFFX1 \registers_reg[165][0]  ( .D(n8019), .E(n1023), .CK(clk), .Q(
        \registers[165][0] ) );
  EDFFX1 \registers_reg[161][7]  ( .D(n8409), .E(n958), .CK(clk), .Q(
        \registers[161][7] ) );
  EDFFX1 \registers_reg[161][6]  ( .D(n8351), .E(n958), .CK(clk), .Q(
        \registers[161][6] ) );
  EDFFX1 \registers_reg[161][5]  ( .D(n8293), .E(n958), .CK(clk), .Q(
        \registers[161][5] ) );
  EDFFX1 \registers_reg[161][4]  ( .D(n8235), .E(n958), .CK(clk), .Q(
        \registers[161][4] ) );
  EDFFX1 \registers_reg[161][3]  ( .D(n8182), .E(n958), .CK(clk), .Q(
        \registers[161][3] ) );
  EDFFX1 \registers_reg[161][2]  ( .D(n8137), .E(n958), .CK(clk), .Q(
        \registers[161][2] ) );
  EDFFX1 \registers_reg[161][1]  ( .D(n8081), .E(n958), .CK(clk), .Q(
        \registers[161][1] ) );
  EDFFX1 \registers_reg[161][0]  ( .D(n8020), .E(n958), .CK(clk), .Q(
        \registers[161][0] ) );
  EDFFX1 \registers_reg[157][7]  ( .D(n8405), .E(n511), .CK(clk), .Q(
        \registers[157][7] ) );
  EDFFX1 \registers_reg[157][6]  ( .D(n8347), .E(n511), .CK(clk), .Q(
        \registers[157][6] ) );
  EDFFX1 \registers_reg[157][5]  ( .D(n8289), .E(n511), .CK(clk), .Q(
        \registers[157][5] ) );
  EDFFX1 \registers_reg[157][4]  ( .D(n8231), .E(n511), .CK(clk), .Q(
        \registers[157][4] ) );
  EDFFX1 \registers_reg[157][3]  ( .D(n8183), .E(n511), .CK(clk), .Q(
        \registers[157][3] ) );
  EDFFX1 \registers_reg[157][2]  ( .D(n8135), .E(n511), .CK(clk), .Q(
        \registers[157][2] ) );
  EDFFX1 \registers_reg[157][1]  ( .D(n8079), .E(n511), .CK(clk), .Q(
        \registers[157][1] ) );
  EDFFX1 \registers_reg[157][0]  ( .D(n8021), .E(n511), .CK(clk), .Q(
        \registers[157][0] ) );
  EDFFX1 \registers_reg[153][7]  ( .D(n8406), .E(n507), .CK(clk), .Q(
        \registers[153][7] ) );
  EDFFX1 \registers_reg[153][6]  ( .D(n8348), .E(n507), .CK(clk), .Q(
        \registers[153][6] ) );
  EDFFX1 \registers_reg[153][5]  ( .D(n8290), .E(n507), .CK(clk), .Q(
        \registers[153][5] ) );
  EDFFX1 \registers_reg[153][4]  ( .D(n8232), .E(n507), .CK(clk), .Q(
        \registers[153][4] ) );
  EDFFX1 \registers_reg[153][3]  ( .D(n8184), .E(n507), .CK(clk), .Q(
        \registers[153][3] ) );
  EDFFX1 \registers_reg[153][2]  ( .D(n8136), .E(n507), .CK(clk), .Q(
        \registers[153][2] ) );
  EDFFX1 \registers_reg[153][1]  ( .D(n8080), .E(n507), .CK(clk), .Q(
        \registers[153][1] ) );
  EDFFX1 \registers_reg[153][0]  ( .D(n8019), .E(n507), .CK(clk), .Q(
        \registers[153][0] ) );
  EDFFX1 \registers_reg[149][7]  ( .D(n8404), .E(n503), .CK(clk), .Q(
        \registers[149][7] ) );
  EDFFX1 \registers_reg[149][6]  ( .D(n8346), .E(n503), .CK(clk), .Q(
        \registers[149][6] ) );
  EDFFX1 \registers_reg[149][5]  ( .D(n8288), .E(n503), .CK(clk), .Q(
        \registers[149][5] ) );
  EDFFX1 \registers_reg[149][4]  ( .D(n8230), .E(n503), .CK(clk), .Q(
        \registers[149][4] ) );
  EDFFX1 \registers_reg[149][3]  ( .D(n8182), .E(n503), .CK(clk), .Q(
        \registers[149][3] ) );
  EDFFX1 \registers_reg[149][2]  ( .D(n8137), .E(n503), .CK(clk), .Q(
        \registers[149][2] ) );
  EDFFX1 \registers_reg[149][1]  ( .D(n8081), .E(n503), .CK(clk), .Q(
        \registers[149][1] ) );
  EDFFX1 \registers_reg[149][0]  ( .D(n8020), .E(n503), .CK(clk), .Q(
        \registers[149][0] ) );
  EDFFX1 \registers_reg[145][7]  ( .D(n8405), .E(n499), .CK(clk), .Q(
        \registers[145][7] ) );
  EDFFX1 \registers_reg[145][6]  ( .D(n8347), .E(n499), .CK(clk), .Q(
        \registers[145][6] ) );
  EDFFX1 \registers_reg[145][5]  ( .D(n8289), .E(n499), .CK(clk), .Q(
        \registers[145][5] ) );
  EDFFX1 \registers_reg[145][4]  ( .D(n8231), .E(n499), .CK(clk), .Q(
        \registers[145][4] ) );
  EDFFX1 \registers_reg[145][3]  ( .D(n8183), .E(n499), .CK(clk), .Q(
        \registers[145][3] ) );
  EDFFX1 \registers_reg[145][2]  ( .D(n8135), .E(n499), .CK(clk), .Q(
        \registers[145][2] ) );
  EDFFX1 \registers_reg[145][1]  ( .D(n8079), .E(n499), .CK(clk), .Q(
        \registers[145][1] ) );
  EDFFX1 \registers_reg[145][0]  ( .D(n8021), .E(n499), .CK(clk), .Q(
        \registers[145][0] ) );
  EDFFX1 \registers_reg[141][7]  ( .D(n8406), .E(n495), .CK(clk), .Q(
        \registers[141][7] ) );
  EDFFX1 \registers_reg[141][6]  ( .D(n8348), .E(n495), .CK(clk), .Q(
        \registers[141][6] ) );
  EDFFX1 \registers_reg[141][5]  ( .D(n8290), .E(n495), .CK(clk), .Q(
        \registers[141][5] ) );
  EDFFX1 \registers_reg[141][4]  ( .D(n8232), .E(n495), .CK(clk), .Q(
        \registers[141][4] ) );
  EDFFX1 \registers_reg[141][3]  ( .D(n8184), .E(n495), .CK(clk), .Q(
        \registers[141][3] ) );
  EDFFX1 \registers_reg[141][2]  ( .D(n8136), .E(n495), .CK(clk), .Q(
        \registers[141][2] ) );
  EDFFX1 \registers_reg[141][1]  ( .D(n8080), .E(n495), .CK(clk), .Q(
        \registers[141][1] ) );
  EDFFX1 \registers_reg[141][0]  ( .D(n8019), .E(n495), .CK(clk), .Q(
        \registers[141][0] ) );
  EDFFX1 \registers_reg[137][7]  ( .D(n8404), .E(n491), .CK(clk), .Q(
        \registers[137][7] ) );
  EDFFX1 \registers_reg[137][6]  ( .D(n8346), .E(n491), .CK(clk), .Q(
        \registers[137][6] ) );
  EDFFX1 \registers_reg[137][5]  ( .D(n8288), .E(n491), .CK(clk), .Q(
        \registers[137][5] ) );
  EDFFX1 \registers_reg[137][4]  ( .D(n8230), .E(n491), .CK(clk), .Q(
        \registers[137][4] ) );
  EDFFX1 \registers_reg[137][3]  ( .D(n8182), .E(n491), .CK(clk), .Q(
        \registers[137][3] ) );
  EDFFX1 \registers_reg[137][2]  ( .D(n8137), .E(n491), .CK(clk), .Q(
        \registers[137][2] ) );
  EDFFX1 \registers_reg[137][1]  ( .D(n8081), .E(n491), .CK(clk), .Q(
        \registers[137][1] ) );
  EDFFX1 \registers_reg[137][0]  ( .D(n8020), .E(n491), .CK(clk), .Q(
        \registers[137][0] ) );
  EDFFX1 \registers_reg[133][7]  ( .D(n8405), .E(n1019), .CK(clk), .Q(
        \registers[133][7] ) );
  EDFFX1 \registers_reg[133][6]  ( .D(n8347), .E(n1019), .CK(clk), .Q(
        \registers[133][6] ) );
  EDFFX1 \registers_reg[133][5]  ( .D(n8289), .E(n1019), .CK(clk), .Q(
        \registers[133][5] ) );
  EDFFX1 \registers_reg[133][4]  ( .D(n8231), .E(n1019), .CK(clk), .Q(
        \registers[133][4] ) );
  EDFFX1 \registers_reg[133][3]  ( .D(n8183), .E(n1019), .CK(clk), .Q(
        \registers[133][3] ) );
  EDFFX1 \registers_reg[133][2]  ( .D(n8135), .E(n1019), .CK(clk), .Q(
        \registers[133][2] ) );
  EDFFX1 \registers_reg[133][1]  ( .D(n8079), .E(n1019), .CK(clk), .Q(
        \registers[133][1] ) );
  EDFFX1 \registers_reg[133][0]  ( .D(n8021), .E(n1019), .CK(clk), .Q(
        \registers[133][0] ) );
  EDFFX1 \registers_reg[129][7]  ( .D(n8407), .E(n955), .CK(clk), .Q(
        \registers[129][7] ) );
  EDFFX1 \registers_reg[129][6]  ( .D(n8349), .E(n955), .CK(clk), .Q(
        \registers[129][6] ) );
  EDFFX1 \registers_reg[129][5]  ( .D(n8291), .E(n955), .CK(clk), .Q(
        \registers[129][5] ) );
  EDFFX1 \registers_reg[129][4]  ( .D(n8233), .E(n955), .CK(clk), .Q(
        \registers[129][4] ) );
  EDFFX1 \registers_reg[129][3]  ( .D(n8186), .E(n955), .CK(clk), .Q(
        \registers[129][3] ) );
  EDFFX1 \registers_reg[129][2]  ( .D(n8138), .E(n955), .CK(clk), .Q(
        \registers[129][2] ) );
  EDFFX1 \registers_reg[129][1]  ( .D(n8082), .E(n955), .CK(clk), .Q(
        \registers[129][1] ) );
  EDFFX1 \registers_reg[129][0]  ( .D(n8022), .E(n955), .CK(clk), .Q(
        \registers[129][0] ) );
  EDFFX1 \registers_reg[125][7]  ( .D(n8421), .E(n487), .CK(clk), .Q(
        \registers[125][7] ) );
  EDFFX1 \registers_reg[125][6]  ( .D(n8363), .E(n487), .CK(clk), .Q(
        \registers[125][6] ) );
  EDFFX1 \registers_reg[125][5]  ( .D(n8305), .E(n487), .CK(clk), .Q(
        \registers[125][5] ) );
  EDFFX1 \registers_reg[125][4]  ( .D(n8247), .E(n487), .CK(clk), .Q(
        \registers[125][4] ) );
  EDFFX1 \registers_reg[125][3]  ( .D(n8195), .E(n487), .CK(clk), .Q(
        \registers[125][3] ) );
  EDFFX1 \registers_reg[125][2]  ( .D(n8150), .E(n487), .CK(clk), .Q(
        \registers[125][2] ) );
  EDFFX1 \registers_reg[125][1]  ( .D(n8094), .E(n487), .CK(clk), .Q(
        \registers[125][1] ) );
  EDFFX1 \registers_reg[125][0]  ( .D(n8034), .E(n487), .CK(clk), .Q(
        \registers[125][0] ) );
  EDFFX1 \registers_reg[121][7]  ( .D(n8419), .E(n483), .CK(clk), .Q(
        \registers[121][7] ) );
  EDFFX1 \registers_reg[121][6]  ( .D(n8361), .E(n483), .CK(clk), .Q(
        \registers[121][6] ) );
  EDFFX1 \registers_reg[121][5]  ( .D(n8303), .E(n483), .CK(clk), .Q(
        \registers[121][5] ) );
  EDFFX1 \registers_reg[121][4]  ( .D(n8245), .E(n483), .CK(clk), .Q(
        \registers[121][4] ) );
  EDFFX1 \registers_reg[121][3]  ( .D(n8196), .E(n483), .CK(clk), .Q(
        \registers[121][3] ) );
  EDFFX1 \registers_reg[121][2]  ( .D(n8151), .E(n483), .CK(clk), .Q(
        \registers[121][2] ) );
  EDFFX1 \registers_reg[121][1]  ( .D(n8095), .E(n483), .CK(clk), .Q(
        \registers[121][1] ) );
  EDFFX1 \registers_reg[121][0]  ( .D(n8035), .E(n483), .CK(clk), .Q(
        \registers[121][0] ) );
  EDFFX1 \registers_reg[117][7]  ( .D(n8420), .E(n479), .CK(clk), .Q(
        \registers[117][7] ) );
  EDFFX1 \registers_reg[117][6]  ( .D(n8362), .E(n479), .CK(clk), .Q(
        \registers[117][6] ) );
  EDFFX1 \registers_reg[117][5]  ( .D(n8304), .E(n479), .CK(clk), .Q(
        \registers[117][5] ) );
  EDFFX1 \registers_reg[117][4]  ( .D(n8246), .E(n479), .CK(clk), .Q(
        \registers[117][4] ) );
  EDFFX1 \registers_reg[117][3]  ( .D(n8194), .E(n479), .CK(clk), .Q(
        \registers[117][3] ) );
  EDFFX1 \registers_reg[117][2]  ( .D(n8736), .E(n479), .CK(clk), .Q(
        \registers[117][2] ) );
  EDFFX1 \registers_reg[117][1]  ( .D(n8708), .E(n479), .CK(clk), .Q(
        \registers[117][1] ) );
  EDFFX1 \registers_reg[117][0]  ( .D(n8036), .E(n479), .CK(clk), .Q(
        \registers[117][0] ) );
  EDFFX1 \registers_reg[113][7]  ( .D(n8421), .E(n475), .CK(clk), .Q(
        \registers[113][7] ) );
  EDFFX1 \registers_reg[113][6]  ( .D(n8363), .E(n475), .CK(clk), .Q(
        \registers[113][6] ) );
  EDFFX1 \registers_reg[113][5]  ( .D(n8305), .E(n475), .CK(clk), .Q(
        \registers[113][5] ) );
  EDFFX1 \registers_reg[113][4]  ( .D(n8247), .E(n475), .CK(clk), .Q(
        \registers[113][4] ) );
  EDFFX1 \registers_reg[113][3]  ( .D(n8195), .E(n475), .CK(clk), .Q(
        \registers[113][3] ) );
  EDFFX1 \registers_reg[113][2]  ( .D(n8147), .E(n475), .CK(clk), .Q(
        \registers[113][2] ) );
  EDFFX1 \registers_reg[113][1]  ( .D(n8091), .E(n475), .CK(clk), .Q(
        \registers[113][1] ) );
  EDFFX1 \registers_reg[113][0]  ( .D(n8031), .E(n475), .CK(clk), .Q(
        \registers[113][0] ) );
  EDFFX1 \registers_reg[109][7]  ( .D(n8419), .E(n471), .CK(clk), .Q(
        \registers[109][7] ) );
  EDFFX1 \registers_reg[109][6]  ( .D(n8361), .E(n471), .CK(clk), .Q(
        \registers[109][6] ) );
  EDFFX1 \registers_reg[109][5]  ( .D(n8303), .E(n471), .CK(clk), .Q(
        \registers[109][5] ) );
  EDFFX1 \registers_reg[109][4]  ( .D(n8245), .E(n471), .CK(clk), .Q(
        \registers[109][4] ) );
  EDFFX1 \registers_reg[109][3]  ( .D(n8196), .E(n471), .CK(clk), .Q(
        \registers[109][3] ) );
  EDFFX1 \registers_reg[109][2]  ( .D(n8148), .E(n471), .CK(clk), .Q(
        \registers[109][2] ) );
  EDFFX1 \registers_reg[109][1]  ( .D(n8092), .E(n471), .CK(clk), .Q(
        \registers[109][1] ) );
  EDFFX1 \registers_reg[109][0]  ( .D(n8032), .E(n471), .CK(clk), .Q(
        \registers[109][0] ) );
  EDFFX1 \registers_reg[105][7]  ( .D(n8420), .E(n467), .CK(clk), .Q(
        \registers[105][7] ) );
  EDFFX1 \registers_reg[105][6]  ( .D(n8362), .E(n467), .CK(clk), .Q(
        \registers[105][6] ) );
  EDFFX1 \registers_reg[105][5]  ( .D(n8304), .E(n467), .CK(clk), .Q(
        \registers[105][5] ) );
  EDFFX1 \registers_reg[105][4]  ( .D(n8246), .E(n467), .CK(clk), .Q(
        \registers[105][4] ) );
  EDFFX1 \registers_reg[105][3]  ( .D(n8191), .E(n467), .CK(clk), .Q(
        \registers[105][3] ) );
  EDFFX1 \registers_reg[105][2]  ( .D(n8149), .E(n467), .CK(clk), .Q(
        \registers[105][2] ) );
  EDFFX1 \registers_reg[105][1]  ( .D(n8093), .E(n467), .CK(clk), .Q(
        \registers[105][1] ) );
  EDFFX1 \registers_reg[105][0]  ( .D(n8033), .E(n467), .CK(clk), .Q(
        \registers[105][0] ) );
  EDFFX1 \registers_reg[101][7]  ( .D(n8416), .E(n952), .CK(clk), .Q(
        \registers[101][7] ) );
  EDFFX1 \registers_reg[101][6]  ( .D(n8358), .E(n952), .CK(clk), .Q(
        \registers[101][6] ) );
  EDFFX1 \registers_reg[101][5]  ( .D(n8300), .E(n952), .CK(clk), .Q(
        \registers[101][5] ) );
  EDFFX1 \registers_reg[101][4]  ( .D(n8242), .E(n952), .CK(clk), .Q(
        \registers[101][4] ) );
  EDFFX1 \registers_reg[101][3]  ( .D(n8192), .E(n952), .CK(clk), .Q(
        \registers[101][3] ) );
  EDFFX1 \registers_reg[101][2]  ( .D(n8147), .E(n952), .CK(clk), .Q(
        \registers[101][2] ) );
  EDFFX1 \registers_reg[101][1]  ( .D(n8091), .E(n952), .CK(clk), .Q(
        \registers[101][1] ) );
  EDFFX1 \registers_reg[101][0]  ( .D(n8031), .E(n952), .CK(clk), .Q(
        \registers[101][0] ) );
  EDFFX1 \registers_reg[97][7]  ( .D(n8417), .E(n948), .CK(clk), .Q(
        \registers[97][7] ) );
  EDFFX1 \registers_reg[97][6]  ( .D(n8359), .E(n948), .CK(clk), .Q(
        \registers[97][6] ) );
  EDFFX1 \registers_reg[97][5]  ( .D(n8301), .E(n948), .CK(clk), .Q(
        \registers[97][5] ) );
  EDFFX1 \registers_reg[97][4]  ( .D(n8243), .E(n948), .CK(clk), .Q(
        \registers[97][4] ) );
  EDFFX1 \registers_reg[97][3]  ( .D(n8193), .E(n948), .CK(clk), .Q(
        \registers[97][3] ) );
  EDFFX1 \registers_reg[97][2]  ( .D(n8148), .E(n948), .CK(clk), .Q(
        \registers[97][2] ) );
  EDFFX1 \registers_reg[97][1]  ( .D(n8092), .E(n948), .CK(clk), .Q(
        \registers[97][1] ) );
  EDFFX1 \registers_reg[97][0]  ( .D(n8032), .E(n948), .CK(clk), .Q(
        \registers[97][0] ) );
  EDFFX1 \registers_reg[93][7]  ( .D(n8418), .E(n463), .CK(clk), .Q(
        \registers[93][7] ) );
  EDFFX1 \registers_reg[93][6]  ( .D(n8360), .E(n463), .CK(clk), .Q(
        \registers[93][6] ) );
  EDFFX1 \registers_reg[93][5]  ( .D(n8302), .E(n463), .CK(clk), .Q(
        \registers[93][5] ) );
  EDFFX1 \registers_reg[93][4]  ( .D(n8244), .E(n463), .CK(clk), .Q(
        \registers[93][4] ) );
  EDFFX1 \registers_reg[93][3]  ( .D(n8191), .E(n463), .CK(clk), .Q(
        \registers[93][3] ) );
  EDFFX1 \registers_reg[93][2]  ( .D(n8149), .E(n463), .CK(clk), .Q(
        \registers[93][2] ) );
  EDFFX1 \registers_reg[93][1]  ( .D(n8093), .E(n463), .CK(clk), .Q(
        \registers[93][1] ) );
  EDFFX1 \registers_reg[93][0]  ( .D(n8033), .E(n463), .CK(clk), .Q(
        \registers[93][0] ) );
  EDFFX1 \registers_reg[89][7]  ( .D(n8416), .E(n459), .CK(clk), .Q(
        \registers[89][7] ) );
  EDFFX1 \registers_reg[89][6]  ( .D(n8358), .E(n459), .CK(clk), .Q(
        \registers[89][6] ) );
  EDFFX1 \registers_reg[89][5]  ( .D(n8300), .E(n459), .CK(clk), .Q(
        \registers[89][5] ) );
  EDFFX1 \registers_reg[89][4]  ( .D(n8242), .E(n459), .CK(clk), .Q(
        \registers[89][4] ) );
  EDFFX1 \registers_reg[89][3]  ( .D(n8192), .E(n459), .CK(clk), .Q(
        \registers[89][3] ) );
  EDFFX1 \registers_reg[89][2]  ( .D(n8147), .E(n459), .CK(clk), .Q(
        \registers[89][2] ) );
  EDFFX1 \registers_reg[89][1]  ( .D(n8091), .E(n459), .CK(clk), .Q(
        \registers[89][1] ) );
  EDFFX1 \registers_reg[89][0]  ( .D(n8031), .E(n459), .CK(clk), .Q(
        \registers[89][0] ) );
  EDFFX1 \registers_reg[85][7]  ( .D(n8417), .E(n455), .CK(clk), .Q(
        \registers[85][7] ) );
  EDFFX1 \registers_reg[85][6]  ( .D(n8359), .E(n455), .CK(clk), .Q(
        \registers[85][6] ) );
  EDFFX1 \registers_reg[85][5]  ( .D(n8301), .E(n455), .CK(clk), .Q(
        \registers[85][5] ) );
  EDFFX1 \registers_reg[85][4]  ( .D(n8243), .E(n455), .CK(clk), .Q(
        \registers[85][4] ) );
  EDFFX1 \registers_reg[85][3]  ( .D(n8193), .E(n455), .CK(clk), .Q(
        \registers[85][3] ) );
  EDFFX1 \registers_reg[85][2]  ( .D(n8148), .E(n455), .CK(clk), .Q(
        \registers[85][2] ) );
  EDFFX1 \registers_reg[85][1]  ( .D(n8092), .E(n455), .CK(clk), .Q(
        \registers[85][1] ) );
  EDFFX1 \registers_reg[85][0]  ( .D(n8032), .E(n455), .CK(clk), .Q(
        \registers[85][0] ) );
  EDFFX1 \registers_reg[81][7]  ( .D(n8418), .E(n451), .CK(clk), .Q(
        \registers[81][7] ) );
  EDFFX1 \registers_reg[81][6]  ( .D(n8360), .E(n451), .CK(clk), .Q(
        \registers[81][6] ) );
  EDFFX1 \registers_reg[81][5]  ( .D(n8302), .E(n451), .CK(clk), .Q(
        \registers[81][5] ) );
  EDFFX1 \registers_reg[81][4]  ( .D(n8244), .E(n451), .CK(clk), .Q(
        \registers[81][4] ) );
  EDFFX1 \registers_reg[81][3]  ( .D(n8191), .E(n451), .CK(clk), .Q(
        \registers[81][3] ) );
  EDFFX1 \registers_reg[81][2]  ( .D(n8149), .E(n451), .CK(clk), .Q(
        \registers[81][2] ) );
  EDFFX1 \registers_reg[81][1]  ( .D(n8093), .E(n451), .CK(clk), .Q(
        \registers[81][1] ) );
  EDFFX1 \registers_reg[81][0]  ( .D(n8033), .E(n451), .CK(clk), .Q(
        \registers[81][0] ) );
  EDFFX1 \registers_reg[77][7]  ( .D(n8416), .E(n447), .CK(clk), .Q(
        \registers[77][7] ) );
  EDFFX1 \registers_reg[77][6]  ( .D(n8358), .E(n447), .CK(clk), .Q(
        \registers[77][6] ) );
  EDFFX1 \registers_reg[77][5]  ( .D(n8300), .E(n447), .CK(clk), .Q(
        \registers[77][5] ) );
  EDFFX1 \registers_reg[77][4]  ( .D(n8242), .E(n447), .CK(clk), .Q(
        \registers[77][4] ) );
  EDFFX1 \registers_reg[77][3]  ( .D(n8192), .E(n447), .CK(clk), .Q(
        \registers[77][3] ) );
  EDFFX1 \registers_reg[77][2]  ( .D(n8147), .E(n447), .CK(clk), .Q(
        \registers[77][2] ) );
  EDFFX1 \registers_reg[77][1]  ( .D(n8091), .E(n447), .CK(clk), .Q(
        \registers[77][1] ) );
  EDFFX1 \registers_reg[77][0]  ( .D(n8031), .E(n447), .CK(clk), .Q(
        \registers[77][0] ) );
  EDFFX1 \registers_reg[73][7]  ( .D(n8417), .E(n443), .CK(clk), .Q(
        \registers[73][7] ) );
  EDFFX1 \registers_reg[73][6]  ( .D(n8359), .E(n443), .CK(clk), .Q(
        \registers[73][6] ) );
  EDFFX1 \registers_reg[73][5]  ( .D(n8301), .E(n443), .CK(clk), .Q(
        \registers[73][5] ) );
  EDFFX1 \registers_reg[73][4]  ( .D(n8243), .E(n443), .CK(clk), .Q(
        \registers[73][4] ) );
  EDFFX1 \registers_reg[73][3]  ( .D(n8193), .E(n443), .CK(clk), .Q(
        \registers[73][3] ) );
  EDFFX1 \registers_reg[73][2]  ( .D(n8148), .E(n443), .CK(clk), .Q(
        \registers[73][2] ) );
  EDFFX1 \registers_reg[73][1]  ( .D(n8092), .E(n443), .CK(clk), .Q(
        \registers[73][1] ) );
  EDFFX1 \registers_reg[73][0]  ( .D(n8032), .E(n443), .CK(clk), .Q(
        \registers[73][0] ) );
  EDFFX1 \registers_reg[69][7]  ( .D(n8418), .E(n945), .CK(clk), .Q(
        \registers[69][7] ) );
  EDFFX1 \registers_reg[69][6]  ( .D(n8360), .E(n945), .CK(clk), .Q(
        \registers[69][6] ) );
  EDFFX1 \registers_reg[69][5]  ( .D(n8302), .E(n945), .CK(clk), .Q(
        \registers[69][5] ) );
  EDFFX1 \registers_reg[69][4]  ( .D(n8244), .E(n945), .CK(clk), .Q(
        \registers[69][4] ) );
  EDFFX1 \registers_reg[69][3]  ( .D(n8191), .E(n945), .CK(clk), .Q(
        \registers[69][3] ) );
  EDFFX1 \registers_reg[69][2]  ( .D(n8149), .E(n945), .CK(clk), .Q(
        \registers[69][2] ) );
  EDFFX1 \registers_reg[69][1]  ( .D(n8093), .E(n945), .CK(clk), .Q(
        \registers[69][1] ) );
  EDFFX1 \registers_reg[69][0]  ( .D(n8033), .E(n945), .CK(clk), .Q(
        \registers[69][0] ) );
  EDFFX1 \registers_reg[65][7]  ( .D(n8416), .E(n941), .CK(clk), .Q(
        \registers[65][7] ) );
  EDFFX1 \registers_reg[65][6]  ( .D(n8358), .E(n941), .CK(clk), .Q(
        \registers[65][6] ) );
  EDFFX1 \registers_reg[65][5]  ( .D(n8300), .E(n941), .CK(clk), .Q(
        \registers[65][5] ) );
  EDFFX1 \registers_reg[65][4]  ( .D(n8242), .E(n941), .CK(clk), .Q(
        \registers[65][4] ) );
  EDFFX1 \registers_reg[65][3]  ( .D(n8192), .E(n941), .CK(clk), .Q(
        \registers[65][3] ) );
  EDFFX1 \registers_reg[65][2]  ( .D(n8144), .E(n941), .CK(clk), .Q(
        \registers[65][2] ) );
  EDFFX1 \registers_reg[65][1]  ( .D(n8088), .E(n941), .CK(clk), .Q(
        \registers[65][1] ) );
  EDFFX1 \registers_reg[65][0]  ( .D(n8028), .E(n941), .CK(clk), .Q(
        \registers[65][0] ) );
  EDFFX1 \registers_reg[61][7]  ( .D(n8418), .E(n439), .CK(clk), .Q(
        \registers[61][7] ) );
  EDFFX1 \registers_reg[61][6]  ( .D(n8360), .E(n439), .CK(clk), .Q(
        \registers[61][6] ) );
  EDFFX1 \registers_reg[61][5]  ( .D(n8302), .E(n439), .CK(clk), .Q(
        \registers[61][5] ) );
  EDFFX1 \registers_reg[61][4]  ( .D(n8244), .E(n439), .CK(clk), .Q(
        \registers[61][4] ) );
  EDFFX1 \registers_reg[61][3]  ( .D(n8191), .E(n439), .CK(clk), .Q(
        \registers[61][3] ) );
  EDFFX1 \registers_reg[61][2]  ( .D(n8146), .E(n439), .CK(clk), .Q(
        \registers[61][2] ) );
  EDFFX1 \registers_reg[61][1]  ( .D(n8090), .E(n439), .CK(clk), .Q(
        \registers[61][1] ) );
  EDFFX1 \registers_reg[61][0]  ( .D(n8030), .E(n439), .CK(clk), .Q(
        \registers[61][0] ) );
  EDFFX1 \registers_reg[57][7]  ( .D(n8416), .E(n435), .CK(clk), .Q(
        \registers[57][7] ) );
  EDFFX1 \registers_reg[57][6]  ( .D(n8358), .E(n435), .CK(clk), .Q(
        \registers[57][6] ) );
  EDFFX1 \registers_reg[57][5]  ( .D(n8300), .E(n435), .CK(clk), .Q(
        \registers[57][5] ) );
  EDFFX1 \registers_reg[57][4]  ( .D(n8242), .E(n435), .CK(clk), .Q(
        \registers[57][4] ) );
  EDFFX1 \registers_reg[57][3]  ( .D(n8192), .E(n435), .CK(clk), .Q(
        \registers[57][3] ) );
  EDFFX1 \registers_reg[57][2]  ( .D(n8144), .E(n435), .CK(clk), .Q(
        \registers[57][2] ) );
  EDFFX1 \registers_reg[57][1]  ( .D(n8088), .E(n435), .CK(clk), .Q(
        \registers[57][1] ) );
  EDFFX1 \registers_reg[57][0]  ( .D(n8028), .E(n435), .CK(clk), .Q(
        \registers[57][0] ) );
  EDFFX1 \registers_reg[53][7]  ( .D(n8417), .E(n431), .CK(clk), .Q(
        \registers[53][7] ) );
  EDFFX1 \registers_reg[53][6]  ( .D(n8359), .E(n431), .CK(clk), .Q(
        \registers[53][6] ) );
  EDFFX1 \registers_reg[53][5]  ( .D(n8301), .E(n431), .CK(clk), .Q(
        \registers[53][5] ) );
  EDFFX1 \registers_reg[53][4]  ( .D(n8243), .E(n431), .CK(clk), .Q(
        \registers[53][4] ) );
  EDFFX1 \registers_reg[53][3]  ( .D(n8193), .E(n431), .CK(clk), .Q(
        \registers[53][3] ) );
  EDFFX1 \registers_reg[53][2]  ( .D(n8145), .E(n431), .CK(clk), .Q(
        \registers[53][2] ) );
  EDFFX1 \registers_reg[53][1]  ( .D(n8089), .E(n431), .CK(clk), .Q(
        \registers[53][1] ) );
  EDFFX1 \registers_reg[53][0]  ( .D(n8029), .E(n431), .CK(clk), .Q(
        \registers[53][0] ) );
  EDFFX1 \registers_reg[49][7]  ( .D(n8413), .E(n427), .CK(clk), .Q(
        \registers[49][7] ) );
  EDFFX1 \registers_reg[49][6]  ( .D(n8355), .E(n427), .CK(clk), .Q(
        \registers[49][6] ) );
  EDFFX1 \registers_reg[49][5]  ( .D(n8297), .E(n427), .CK(clk), .Q(
        \registers[49][5] ) );
  EDFFX1 \registers_reg[49][4]  ( .D(n8239), .E(n427), .CK(clk), .Q(
        \registers[49][4] ) );
  EDFFX1 \registers_reg[49][3]  ( .D(n8191), .E(n427), .CK(clk), .Q(
        \registers[49][3] ) );
  EDFFX1 \registers_reg[49][2]  ( .D(n8146), .E(n427), .CK(clk), .Q(
        \registers[49][2] ) );
  EDFFX1 \registers_reg[49][1]  ( .D(n8090), .E(n427), .CK(clk), .Q(
        \registers[49][1] ) );
  EDFFX1 \registers_reg[49][0]  ( .D(n8030), .E(n427), .CK(clk), .Q(
        \registers[49][0] ) );
  EDFFX1 \registers_reg[45][7]  ( .D(n8414), .E(n423), .CK(clk), .Q(
        \registers[45][7] ) );
  EDFFX1 \registers_reg[45][6]  ( .D(n8356), .E(n423), .CK(clk), .Q(
        \registers[45][6] ) );
  EDFFX1 \registers_reg[45][5]  ( .D(n8298), .E(n423), .CK(clk), .Q(
        \registers[45][5] ) );
  EDFFX1 \registers_reg[45][4]  ( .D(n8240), .E(n423), .CK(clk), .Q(
        \registers[45][4] ) );
  EDFFX1 \registers_reg[45][3]  ( .D(n8192), .E(n423), .CK(clk), .Q(
        \registers[45][3] ) );
  EDFFX1 \registers_reg[45][2]  ( .D(n8144), .E(n423), .CK(clk), .Q(
        \registers[45][2] ) );
  EDFFX1 \registers_reg[45][1]  ( .D(n8088), .E(n423), .CK(clk), .Q(
        \registers[45][1] ) );
  EDFFX1 \registers_reg[45][0]  ( .D(n8028), .E(n423), .CK(clk), .Q(
        \registers[45][0] ) );
  EDFFX1 \registers_reg[41][7]  ( .D(n8415), .E(n419), .CK(clk), .Q(
        \registers[41][7] ) );
  EDFFX1 \registers_reg[41][6]  ( .D(n8357), .E(n419), .CK(clk), .Q(
        \registers[41][6] ) );
  EDFFX1 \registers_reg[41][5]  ( .D(n8299), .E(n419), .CK(clk), .Q(
        \registers[41][5] ) );
  EDFFX1 \registers_reg[41][4]  ( .D(n8241), .E(n419), .CK(clk), .Q(
        \registers[41][4] ) );
  EDFFX1 \registers_reg[41][3]  ( .D(n8190), .E(n419), .CK(clk), .Q(
        \registers[41][3] ) );
  EDFFX1 \registers_reg[41][2]  ( .D(n8145), .E(n419), .CK(clk), .Q(
        \registers[41][2] ) );
  EDFFX1 \registers_reg[41][1]  ( .D(n8089), .E(n419), .CK(clk), .Q(
        \registers[41][1] ) );
  EDFFX1 \registers_reg[41][0]  ( .D(n8029), .E(n419), .CK(clk), .Q(
        \registers[41][0] ) );
  EDFFX1 \registers_reg[37][7]  ( .D(n8413), .E(n938), .CK(clk), .Q(
        \registers[37][7] ) );
  EDFFX1 \registers_reg[37][6]  ( .D(n8355), .E(n938), .CK(clk), .Q(
        \registers[37][6] ) );
  EDFFX1 \registers_reg[37][5]  ( .D(n8297), .E(n938), .CK(clk), .Q(
        \registers[37][5] ) );
  EDFFX1 \registers_reg[37][4]  ( .D(n8239), .E(n938), .CK(clk), .Q(
        \registers[37][4] ) );
  EDFFX1 \registers_reg[37][3]  ( .D(n8188), .E(n938), .CK(clk), .Q(
        \registers[37][3] ) );
  EDFFX1 \registers_reg[37][2]  ( .D(n8146), .E(n938), .CK(clk), .Q(
        \registers[37][2] ) );
  EDFFX1 \registers_reg[37][1]  ( .D(n8090), .E(n938), .CK(clk), .Q(
        \registers[37][1] ) );
  EDFFX1 \registers_reg[37][0]  ( .D(n8030), .E(n938), .CK(clk), .Q(
        \registers[37][0] ) );
  EDFFX1 \registers_reg[33][7]  ( .D(n8414), .E(n934), .CK(clk), .Q(
        \registers[33][7] ) );
  EDFFX1 \registers_reg[33][6]  ( .D(n8356), .E(n934), .CK(clk), .Q(
        \registers[33][6] ) );
  EDFFX1 \registers_reg[33][5]  ( .D(n8298), .E(n934), .CK(clk), .Q(
        \registers[33][5] ) );
  EDFFX1 \registers_reg[33][4]  ( .D(n8240), .E(n934), .CK(clk), .Q(
        \registers[33][4] ) );
  EDFFX1 \registers_reg[33][3]  ( .D(n8189), .E(n934), .CK(clk), .Q(
        \registers[33][3] ) );
  EDFFX1 \registers_reg[33][2]  ( .D(n8144), .E(n934), .CK(clk), .Q(
        \registers[33][2] ) );
  EDFFX1 \registers_reg[33][1]  ( .D(n8088), .E(n934), .CK(clk), .Q(
        \registers[33][1] ) );
  EDFFX1 \registers_reg[33][0]  ( .D(n8028), .E(n934), .CK(clk), .Q(
        \registers[33][0] ) );
  EDFFX1 \registers_reg[29][7]  ( .D(n8415), .E(n415), .CK(clk), .Q(
        \registers[29][7] ) );
  EDFFX1 \registers_reg[29][6]  ( .D(n8357), .E(n415), .CK(clk), .Q(
        \registers[29][6] ) );
  EDFFX1 \registers_reg[29][5]  ( .D(n8299), .E(n415), .CK(clk), .Q(
        \registers[29][5] ) );
  EDFFX1 \registers_reg[29][4]  ( .D(n8241), .E(n415), .CK(clk), .Q(
        \registers[29][4] ) );
  EDFFX1 \registers_reg[29][3]  ( .D(n8190), .E(n415), .CK(clk), .Q(
        \registers[29][3] ) );
  EDFFX1 \registers_reg[29][2]  ( .D(n8145), .E(n415), .CK(clk), .Q(
        \registers[29][2] ) );
  EDFFX1 \registers_reg[29][1]  ( .D(n8089), .E(n415), .CK(clk), .Q(
        \registers[29][1] ) );
  EDFFX1 \registers_reg[29][0]  ( .D(n8029), .E(n415), .CK(clk), .Q(
        \registers[29][0] ) );
  EDFFX1 \registers_reg[25][7]  ( .D(n8413), .E(n411), .CK(clk), .Q(
        \registers[25][7] ) );
  EDFFX1 \registers_reg[25][6]  ( .D(n8355), .E(n411), .CK(clk), .Q(
        \registers[25][6] ) );
  EDFFX1 \registers_reg[25][5]  ( .D(n8297), .E(n411), .CK(clk), .Q(
        \registers[25][5] ) );
  EDFFX1 \registers_reg[25][4]  ( .D(n8239), .E(n411), .CK(clk), .Q(
        \registers[25][4] ) );
  EDFFX1 \registers_reg[25][3]  ( .D(n8188), .E(n411), .CK(clk), .Q(
        \registers[25][3] ) );
  EDFFX1 \registers_reg[25][2]  ( .D(n8146), .E(n411), .CK(clk), .Q(
        \registers[25][2] ) );
  EDFFX1 \registers_reg[25][1]  ( .D(n8090), .E(n411), .CK(clk), .Q(
        \registers[25][1] ) );
  EDFFX1 \registers_reg[25][0]  ( .D(n8030), .E(n411), .CK(clk), .Q(
        \registers[25][0] ) );
  EDFFX1 \registers_reg[21][7]  ( .D(n8414), .E(n407), .CK(clk), .Q(
        \registers[21][7] ) );
  EDFFX1 \registers_reg[21][6]  ( .D(n8356), .E(n407), .CK(clk), .Q(
        \registers[21][6] ) );
  EDFFX1 \registers_reg[21][5]  ( .D(n8298), .E(n407), .CK(clk), .Q(
        \registers[21][5] ) );
  EDFFX1 \registers_reg[21][4]  ( .D(n8240), .E(n407), .CK(clk), .Q(
        \registers[21][4] ) );
  EDFFX1 \registers_reg[21][3]  ( .D(n8189), .E(n407), .CK(clk), .Q(
        \registers[21][3] ) );
  EDFFX1 \registers_reg[21][2]  ( .D(n8144), .E(n407), .CK(clk), .Q(
        \registers[21][2] ) );
  EDFFX1 \registers_reg[21][1]  ( .D(n8088), .E(n407), .CK(clk), .Q(
        \registers[21][1] ) );
  EDFFX1 \registers_reg[21][0]  ( .D(n8028), .E(n407), .CK(clk), .Q(
        \registers[21][0] ) );
  EDFFX1 \registers_reg[17][7]  ( .D(n8415), .E(n403), .CK(clk), .Q(
        \registers[17][7] ) );
  EDFFX1 \registers_reg[17][6]  ( .D(n8357), .E(n403), .CK(clk), .Q(
        \registers[17][6] ) );
  EDFFX1 \registers_reg[17][5]  ( .D(n8299), .E(n403), .CK(clk), .Q(
        \registers[17][5] ) );
  EDFFX1 \registers_reg[17][4]  ( .D(n8241), .E(n403), .CK(clk), .Q(
        \registers[17][4] ) );
  EDFFX1 \registers_reg[17][3]  ( .D(n8190), .E(n403), .CK(clk), .Q(
        \registers[17][3] ) );
  EDFFX1 \registers_reg[17][2]  ( .D(n8145), .E(n403), .CK(clk), .Q(
        \registers[17][2] ) );
  EDFFX1 \registers_reg[17][1]  ( .D(n8089), .E(n403), .CK(clk), .Q(
        \registers[17][1] ) );
  EDFFX1 \registers_reg[17][0]  ( .D(n8029), .E(n403), .CK(clk), .Q(
        \registers[17][0] ) );
  EDFFX1 \registers_reg[13][7]  ( .D(n8413), .E(n399), .CK(clk), .Q(
        \registers[13][7] ) );
  EDFFX1 \registers_reg[13][6]  ( .D(n8355), .E(n399), .CK(clk), .Q(
        \registers[13][6] ) );
  EDFFX1 \registers_reg[13][5]  ( .D(n8297), .E(n399), .CK(clk), .Q(
        \registers[13][5] ) );
  EDFFX1 \registers_reg[13][4]  ( .D(n8239), .E(n399), .CK(clk), .Q(
        \registers[13][4] ) );
  EDFFX1 \registers_reg[13][3]  ( .D(n8188), .E(n399), .CK(clk), .Q(
        \registers[13][3] ) );
  EDFFX1 \registers_reg[13][2]  ( .D(n8143), .E(n399), .CK(clk), .Q(
        \registers[13][2] ) );
  EDFFX1 \registers_reg[13][1]  ( .D(n8087), .E(n399), .CK(clk), .Q(
        \registers[13][1] ) );
  EDFFX1 \registers_reg[13][0]  ( .D(n8027), .E(n399), .CK(clk), .Q(
        \registers[13][0] ) );
  EDFFX1 \registers_reg[9][7]  ( .D(n8414), .E(n395), .CK(clk), .Q(
        \registers[9][7] ) );
  EDFFX1 \registers_reg[9][6]  ( .D(n8356), .E(n395), .CK(clk), .Q(
        \registers[9][6] ) );
  EDFFX1 \registers_reg[9][5]  ( .D(n8298), .E(n395), .CK(clk), .Q(
        \registers[9][5] ), .QN(n1108) );
  EDFFX1 \registers_reg[9][4]  ( .D(n8240), .E(n395), .CK(clk), .Q(
        \registers[9][4] ), .QN(n1109) );
  EDFFX1 \registers_reg[9][3]  ( .D(n8189), .E(n395), .CK(clk), .Q(
        \registers[9][3] ), .QN(n1110) );
  EDFFX1 \registers_reg[9][2]  ( .D(n8141), .E(n395), .CK(clk), .Q(
        \registers[9][2] ), .QN(n1111) );
  EDFFX1 \registers_reg[9][1]  ( .D(n8085), .E(n395), .CK(clk), .Q(
        \registers[9][1] ), .QN(n1112) );
  EDFFX1 \registers_reg[9][0]  ( .D(n8025), .E(n395), .CK(clk), .Q(
        \registers[9][0] ), .QN(n1113) );
  EDFFX1 \registers_reg[5][7]  ( .D(n8415), .E(n1015), .CK(clk), .Q(
        \registers[5][7] ), .QN(n1134) );
  EDFFX1 \registers_reg[5][6]  ( .D(n8357), .E(n1015), .CK(clk), .Q(
        \registers[5][6] ), .QN(n1135) );
  EDFFX1 \registers_reg[5][5]  ( .D(n8299), .E(n1015), .CK(clk), .Q(
        \registers[5][5] ), .QN(n1136) );
  EDFFX1 \registers_reg[5][4]  ( .D(n8241), .E(n1015), .CK(clk), .Q(
        \registers[5][4] ), .QN(n1137) );
  EDFFX1 \registers_reg[5][3]  ( .D(n8190), .E(n1015), .CK(clk), .Q(
        \registers[5][3] ), .QN(n1138) );
  EDFFX1 \registers_reg[5][2]  ( .D(n8142), .E(n1015), .CK(clk), .Q(
        \registers[5][2] ), .QN(n1139) );
  EDFFX1 \registers_reg[5][1]  ( .D(n8086), .E(n1015), .CK(clk), .Q(
        \registers[5][1] ), .QN(n1140) );
  EDFFX1 \registers_reg[5][0]  ( .D(n8026), .E(n1015), .CK(clk), .Q(
        \registers[5][0] ), .QN(n1141) );
  EDFFX1 \registers_reg[1][7]  ( .D(n8417), .E(n391), .CK(clk), .Q(
        \registers[1][7] ), .QN(n1142) );
  EDFFX1 \registers_reg[1][6]  ( .D(n8359), .E(n391), .CK(clk), .Q(
        \registers[1][6] ), .QN(n1143) );
  EDFFX1 \registers_reg[1][5]  ( .D(n8301), .E(n391), .CK(clk), .Q(
        \registers[1][5] ), .QN(n1144) );
  EDFFX1 \registers_reg[1][4]  ( .D(n8243), .E(n391), .CK(clk), .Q(
        \registers[1][4] ), .QN(n1145) );
  EDFFX1 \registers_reg[1][3]  ( .D(n8193), .E(n391), .CK(clk), .Q(
        \registers[1][3] ), .QN(n1146) );
  EDFFX1 \registers_reg[1][2]  ( .D(n8145), .E(n391), .CK(clk), .Q(
        \registers[1][2] ), .QN(n1147) );
  EDFFX1 \registers_reg[1][1]  ( .D(n8089), .E(n391), .CK(clk), .Q(
        \registers[1][1] ), .QN(n1148) );
  EDFFX1 \registers_reg[1][0]  ( .D(n8029), .E(n391), .CK(clk), .Q(
        \registers[1][0] ), .QN(n1149) );
  EDFFX1 \registers_reg[1023][7]  ( .D(n8406), .E(n933), .CK(clk), .Q(
        \registers[1023][7] ) );
  EDFFX1 \registers_reg[1023][6]  ( .D(n8348), .E(n933), .CK(clk), .Q(
        \registers[1023][6] ) );
  EDFFX1 \registers_reg[1023][5]  ( .D(n8290), .E(n933), .CK(clk), .Q(
        \registers[1023][5] ) );
  EDFFX1 \registers_reg[1023][4]  ( .D(n8232), .E(n933), .CK(clk), .Q(
        \registers[1023][4] ) );
  EDFFX1 \registers_reg[1023][3]  ( .D(n8184), .E(n933), .CK(clk), .Q(
        \registers[1023][3] ) );
  EDFFX1 \registers_reg[1023][2]  ( .D(n8136), .E(n933), .CK(clk), .Q(
        \registers[1023][2] ) );
  EDFFX1 \registers_reg[1023][1]  ( .D(n8080), .E(n933), .CK(clk), .Q(
        \registers[1023][1] ) );
  EDFFX1 \registers_reg[1023][0]  ( .D(n8019), .E(n933), .CK(clk), .Q(
        \registers[1023][0] ) );
  EDFFX1 \registers_reg[1019][7]  ( .D(n8395), .E(n929), .CK(clk), .Q(
        \registers[1019][7] ) );
  EDFFX1 \registers_reg[1019][6]  ( .D(n8337), .E(n929), .CK(clk), .Q(
        \registers[1019][6] ) );
  EDFFX1 \registers_reg[1019][5]  ( .D(n8279), .E(n929), .CK(clk), .Q(
        \registers[1019][5] ) );
  EDFFX1 \registers_reg[1019][4]  ( .D(n8221), .E(n929), .CK(clk), .Q(
        \registers[1019][4] ) );
  EDFFX1 \registers_reg[1019][3]  ( .D(n8176), .E(n929), .CK(clk), .Q(
        \registers[1019][3] ) );
  EDFFX1 \registers_reg[1019][2]  ( .D(n8128), .E(n929), .CK(clk), .Q(
        \registers[1019][2] ) );
  EDFFX1 \registers_reg[1019][1]  ( .D(n8072), .E(n929), .CK(clk), .Q(
        \registers[1019][1] ) );
  EDFFX1 \registers_reg[1019][0]  ( .D(n8011), .E(n929), .CK(clk), .Q(
        \registers[1019][0] ) );
  EDFFX1 \registers_reg[1015][7]  ( .D(n8396), .E(n925), .CK(clk), .Q(
        \registers[1015][7] ) );
  EDFFX1 \registers_reg[1015][6]  ( .D(n8338), .E(n925), .CK(clk), .Q(
        \registers[1015][6] ) );
  EDFFX1 \registers_reg[1015][5]  ( .D(n8280), .E(n925), .CK(clk), .Q(
        \registers[1015][5] ) );
  EDFFX1 \registers_reg[1015][4]  ( .D(n8222), .E(n925), .CK(clk), .Q(
        \registers[1015][4] ) );
  EDFFX1 \registers_reg[1015][3]  ( .D(n8177), .E(n925), .CK(clk), .Q(
        \registers[1015][3] ) );
  EDFFX1 \registers_reg[1015][2]  ( .D(n8126), .E(n925), .CK(clk), .Q(
        \registers[1015][2] ) );
  EDFFX1 \registers_reg[1015][1]  ( .D(n8070), .E(n925), .CK(clk), .Q(
        \registers[1015][1] ) );
  EDFFX1 \registers_reg[1015][0]  ( .D(n8012), .E(n925), .CK(clk), .Q(
        \registers[1015][0] ) );
  EDFFX1 \registers_reg[1011][7]  ( .D(n8397), .E(n238), .CK(clk), .Q(
        \registers[1011][7] ) );
  EDFFX1 \registers_reg[1011][6]  ( .D(n8339), .E(n238), .CK(clk), .Q(
        \registers[1011][6] ) );
  EDFFX1 \registers_reg[1011][5]  ( .D(n8281), .E(n238), .CK(clk), .Q(
        \registers[1011][5] ) );
  EDFFX1 \registers_reg[1011][4]  ( .D(n8223), .E(n238), .CK(clk), .Q(
        \registers[1011][4] ) );
  EDFFX1 \registers_reg[1011][3]  ( .D(n8178), .E(n238), .CK(clk), .Q(
        \registers[1011][3] ) );
  EDFFX1 \registers_reg[1011][2]  ( .D(n8127), .E(n238), .CK(clk), .Q(
        \registers[1011][2] ) );
  EDFFX1 \registers_reg[1011][1]  ( .D(n8071), .E(n238), .CK(clk), .Q(
        \registers[1011][1] ) );
  EDFFX1 \registers_reg[1011][0]  ( .D(n8010), .E(n238), .CK(clk), .Q(
        \registers[1011][0] ) );
  EDFFX1 \registers_reg[1007][7]  ( .D(n8395), .E(n234), .CK(clk), .Q(
        \registers[1007][7] ) );
  EDFFX1 \registers_reg[1007][6]  ( .D(n8337), .E(n234), .CK(clk), .Q(
        \registers[1007][6] ) );
  EDFFX1 \registers_reg[1007][5]  ( .D(n8279), .E(n234), .CK(clk), .Q(
        \registers[1007][5] ) );
  EDFFX1 \registers_reg[1007][4]  ( .D(n8221), .E(n234), .CK(clk), .Q(
        \registers[1007][4] ) );
  EDFFX1 \registers_reg[1007][3]  ( .D(n8176), .E(n234), .CK(clk), .Q(
        \registers[1007][3] ) );
  EDFFX1 \registers_reg[1007][2]  ( .D(n8128), .E(n234), .CK(clk), .Q(
        \registers[1007][2] ) );
  EDFFX1 \registers_reg[1007][1]  ( .D(n8072), .E(n234), .CK(clk), .Q(
        \registers[1007][1] ) );
  EDFFX1 \registers_reg[1007][0]  ( .D(n8011), .E(n234), .CK(clk), .Q(
        \registers[1007][0] ) );
  EDFFX1 \registers_reg[1003][7]  ( .D(n8396), .E(n230), .CK(clk), .Q(
        \registers[1003][7] ) );
  EDFFX1 \registers_reg[1003][6]  ( .D(n8338), .E(n230), .CK(clk), .Q(
        \registers[1003][6] ) );
  EDFFX1 \registers_reg[1003][5]  ( .D(n8280), .E(n230), .CK(clk), .Q(
        \registers[1003][5] ) );
  EDFFX1 \registers_reg[1003][4]  ( .D(n8222), .E(n230), .CK(clk), .Q(
        \registers[1003][4] ) );
  EDFFX1 \registers_reg[1003][3]  ( .D(n8174), .E(n230), .CK(clk), .Q(
        \registers[1003][3] ) );
  EDFFX1 \registers_reg[1003][2]  ( .D(n8126), .E(n230), .CK(clk), .Q(
        \registers[1003][2] ) );
  EDFFX1 \registers_reg[1003][1]  ( .D(n8070), .E(n230), .CK(clk), .Q(
        \registers[1003][1] ) );
  EDFFX1 \registers_reg[1003][0]  ( .D(n8012), .E(n230), .CK(clk), .Q(
        \registers[1003][0] ) );
  EDFFX1 \registers_reg[999][7]  ( .D(n8397), .E(n386), .CK(clk), .Q(
        \registers[999][7] ) );
  EDFFX1 \registers_reg[999][6]  ( .D(n8339), .E(n386), .CK(clk), .Q(
        \registers[999][6] ) );
  EDFFX1 \registers_reg[999][5]  ( .D(n8281), .E(n386), .CK(clk), .Q(
        \registers[999][5] ) );
  EDFFX1 \registers_reg[999][4]  ( .D(n8223), .E(n386), .CK(clk), .Q(
        \registers[999][4] ) );
  EDFFX1 \registers_reg[999][3]  ( .D(n8175), .E(n386), .CK(clk), .Q(
        \registers[999][3] ) );
  EDFFX1 \registers_reg[999][2]  ( .D(n8127), .E(n386), .CK(clk), .Q(
        \registers[999][2] ) );
  EDFFX1 \registers_reg[999][1]  ( .D(n8071), .E(n386), .CK(clk), .Q(
        \registers[999][1] ) );
  EDFFX1 \registers_reg[999][0]  ( .D(n8010), .E(n386), .CK(clk), .Q(
        \registers[999][0] ) );
  EDFFX1 \registers_reg[995][7]  ( .D(n8395), .E(n382), .CK(clk), .Q(
        \registers[995][7] ) );
  EDFFX1 \registers_reg[995][6]  ( .D(n8337), .E(n382), .CK(clk), .Q(
        \registers[995][6] ) );
  EDFFX1 \registers_reg[995][5]  ( .D(n8279), .E(n382), .CK(clk), .Q(
        \registers[995][5] ) );
  EDFFX1 \registers_reg[995][4]  ( .D(n8221), .E(n382), .CK(clk), .Q(
        \registers[995][4] ) );
  EDFFX1 \registers_reg[995][3]  ( .D(n8173), .E(n382), .CK(clk), .Q(
        \registers[995][3] ) );
  EDFFX1 \registers_reg[995][2]  ( .D(n8128), .E(n382), .CK(clk), .Q(
        \registers[995][2] ) );
  EDFFX1 \registers_reg[995][1]  ( .D(n8072), .E(n382), .CK(clk), .Q(
        \registers[995][1] ) );
  EDFFX1 \registers_reg[995][0]  ( .D(n8011), .E(n382), .CK(clk), .Q(
        \registers[995][0] ) );
  EDFFX1 \registers_reg[991][7]  ( .D(n8396), .E(n921), .CK(clk), .Q(
        \registers[991][7] ) );
  EDFFX1 \registers_reg[991][6]  ( .D(n8338), .E(n921), .CK(clk), .Q(
        \registers[991][6] ) );
  EDFFX1 \registers_reg[991][5]  ( .D(n8280), .E(n921), .CK(clk), .Q(
        \registers[991][5] ) );
  EDFFX1 \registers_reg[991][4]  ( .D(n8222), .E(n921), .CK(clk), .Q(
        \registers[991][4] ) );
  EDFFX1 \registers_reg[991][3]  ( .D(n8174), .E(n921), .CK(clk), .Q(
        \registers[991][3] ) );
  EDFFX1 \registers_reg[991][2]  ( .D(n8126), .E(n921), .CK(clk), .Q(
        \registers[991][2] ) );
  EDFFX1 \registers_reg[991][1]  ( .D(n8070), .E(n921), .CK(clk), .Q(
        \registers[991][1] ) );
  EDFFX1 \registers_reg[991][0]  ( .D(n8012), .E(n921), .CK(clk), .Q(
        \registers[991][0] ) );
  EDFFX1 \registers_reg[987][7]  ( .D(n8397), .E(n917), .CK(clk), .Q(
        \registers[987][7] ) );
  EDFFX1 \registers_reg[987][6]  ( .D(n8339), .E(n917), .CK(clk), .Q(
        \registers[987][6] ) );
  EDFFX1 \registers_reg[987][5]  ( .D(n8281), .E(n917), .CK(clk), .Q(
        \registers[987][5] ) );
  EDFFX1 \registers_reg[987][4]  ( .D(n8223), .E(n917), .CK(clk), .Q(
        \registers[987][4] ) );
  EDFFX1 \registers_reg[987][3]  ( .D(n8175), .E(n917), .CK(clk), .Q(
        \registers[987][3] ) );
  EDFFX1 \registers_reg[987][2]  ( .D(n8127), .E(n917), .CK(clk), .Q(
        \registers[987][2] ) );
  EDFFX1 \registers_reg[987][1]  ( .D(n8071), .E(n917), .CK(clk), .Q(
        \registers[987][1] ) );
  EDFFX1 \registers_reg[987][0]  ( .D(n8010), .E(n917), .CK(clk), .Q(
        \registers[987][0] ) );
  EDFFX1 \registers_reg[983][7]  ( .D(n8395), .E(n913), .CK(clk), .Q(
        \registers[983][7] ) );
  EDFFX1 \registers_reg[983][6]  ( .D(n8337), .E(n913), .CK(clk), .Q(
        \registers[983][6] ) );
  EDFFX1 \registers_reg[983][5]  ( .D(n8279), .E(n913), .CK(clk), .Q(
        \registers[983][5] ) );
  EDFFX1 \registers_reg[983][4]  ( .D(n8221), .E(n913), .CK(clk), .Q(
        \registers[983][4] ) );
  EDFFX1 \registers_reg[983][3]  ( .D(n8173), .E(n913), .CK(clk), .Q(
        \registers[983][3] ) );
  EDFFX1 \registers_reg[983][2]  ( .D(n8125), .E(n913), .CK(clk), .Q(
        \registers[983][2] ) );
  EDFFX1 \registers_reg[983][1]  ( .D(n8069), .E(n913), .CK(clk), .Q(
        \registers[983][1] ) );
  EDFFX1 \registers_reg[983][0]  ( .D(n8008), .E(n913), .CK(clk), .Q(
        \registers[983][0] ) );
  EDFFX1 \registers_reg[979][7]  ( .D(n8396), .E(n226), .CK(clk), .Q(
        \registers[979][7] ) );
  EDFFX1 \registers_reg[979][6]  ( .D(n8338), .E(n226), .CK(clk), .Q(
        \registers[979][6] ) );
  EDFFX1 \registers_reg[979][5]  ( .D(n8280), .E(n226), .CK(clk), .Q(
        \registers[979][5] ) );
  EDFFX1 \registers_reg[979][4]  ( .D(n8222), .E(n226), .CK(clk), .Q(
        \registers[979][4] ) );
  EDFFX1 \registers_reg[979][3]  ( .D(n8174), .E(n226), .CK(clk), .Q(
        \registers[979][3] ) );
  EDFFX1 \registers_reg[979][2]  ( .D(n8123), .E(n226), .CK(clk), .Q(
        \registers[979][2] ) );
  EDFFX1 \registers_reg[979][1]  ( .D(n8067), .E(n226), .CK(clk), .Q(
        \registers[979][1] ) );
  EDFFX1 \registers_reg[979][0]  ( .D(n8009), .E(n226), .CK(clk), .Q(
        \registers[979][0] ) );
  EDFFX1 \registers_reg[975][7]  ( .D(n8392), .E(n222), .CK(clk), .Q(
        \registers[975][7] ) );
  EDFFX1 \registers_reg[975][6]  ( .D(n8334), .E(n222), .CK(clk), .Q(
        \registers[975][6] ) );
  EDFFX1 \registers_reg[975][5]  ( .D(n8276), .E(n222), .CK(clk), .Q(
        \registers[975][5] ) );
  EDFFX1 \registers_reg[975][4]  ( .D(n8218), .E(n222), .CK(clk), .Q(
        \registers[975][4] ) );
  EDFFX1 \registers_reg[975][3]  ( .D(n8175), .E(n222), .CK(clk), .Q(
        \registers[975][3] ) );
  EDFFX1 \registers_reg[975][2]  ( .D(n8124), .E(n222), .CK(clk), .Q(
        \registers[975][2] ) );
  EDFFX1 \registers_reg[975][1]  ( .D(n8068), .E(n222), .CK(clk), .Q(
        \registers[975][1] ) );
  EDFFX1 \registers_reg[975][0]  ( .D(n8007), .E(n222), .CK(clk), .Q(
        \registers[975][0] ) );
  EDFFX1 \registers_reg[971][7]  ( .D(n8393), .E(n218), .CK(clk), .Q(
        \registers[971][7] ) );
  EDFFX1 \registers_reg[971][6]  ( .D(n8335), .E(n218), .CK(clk), .Q(
        \registers[971][6] ) );
  EDFFX1 \registers_reg[971][5]  ( .D(n8277), .E(n218), .CK(clk), .Q(
        \registers[971][5] ) );
  EDFFX1 \registers_reg[971][4]  ( .D(n8219), .E(n218), .CK(clk), .Q(
        \registers[971][4] ) );
  EDFFX1 \registers_reg[971][3]  ( .D(n8173), .E(n218), .CK(clk), .Q(
        \registers[971][3] ) );
  EDFFX1 \registers_reg[971][2]  ( .D(n8125), .E(n218), .CK(clk), .Q(
        \registers[971][2] ) );
  EDFFX1 \registers_reg[971][1]  ( .D(n8069), .E(n218), .CK(clk), .Q(
        \registers[971][1] ) );
  EDFFX1 \registers_reg[971][0]  ( .D(n8008), .E(n218), .CK(clk), .Q(
        \registers[971][0] ) );
  EDFFX1 \registers_reg[967][7]  ( .D(n8394), .E(n379), .CK(clk), .Q(
        \registers[967][7] ) );
  EDFFX1 \registers_reg[967][6]  ( .D(n8336), .E(n379), .CK(clk), .Q(
        \registers[967][6] ) );
  EDFFX1 \registers_reg[967][5]  ( .D(n8278), .E(n379), .CK(clk), .Q(
        \registers[967][5] ) );
  EDFFX1 \registers_reg[967][4]  ( .D(n8220), .E(n379), .CK(clk), .Q(
        \registers[967][4] ) );
  EDFFX1 \registers_reg[967][3]  ( .D(n8174), .E(n379), .CK(clk), .Q(
        \registers[967][3] ) );
  EDFFX1 \registers_reg[967][2]  ( .D(n8123), .E(n379), .CK(clk), .Q(
        \registers[967][2] ) );
  EDFFX1 \registers_reg[967][1]  ( .D(n8067), .E(n379), .CK(clk), .Q(
        \registers[967][1] ) );
  EDFFX1 \registers_reg[967][0]  ( .D(n8009), .E(n379), .CK(clk), .Q(
        \registers[967][0] ) );
  EDFFX1 \registers_reg[963][7]  ( .D(n8392), .E(n375), .CK(clk), .Q(
        \registers[963][7] ) );
  EDFFX1 \registers_reg[963][6]  ( .D(n8334), .E(n375), .CK(clk), .Q(
        \registers[963][6] ) );
  EDFFX1 \registers_reg[963][5]  ( .D(n8276), .E(n375), .CK(clk), .Q(
        \registers[963][5] ) );
  EDFFX1 \registers_reg[963][4]  ( .D(n8218), .E(n375), .CK(clk), .Q(
        \registers[963][4] ) );
  EDFFX1 \registers_reg[963][3]  ( .D(n8175), .E(n375), .CK(clk), .Q(
        \registers[963][3] ) );
  EDFFX1 \registers_reg[963][2]  ( .D(n8124), .E(n375), .CK(clk), .Q(
        \registers[963][2] ) );
  EDFFX1 \registers_reg[963][1]  ( .D(n8068), .E(n375), .CK(clk), .Q(
        \registers[963][1] ) );
  EDFFX1 \registers_reg[963][0]  ( .D(n8007), .E(n375), .CK(clk), .Q(
        \registers[963][0] ) );
  EDFFX1 \registers_reg[959][7]  ( .D(n8393), .E(n909), .CK(clk), .Q(
        \registers[959][7] ) );
  EDFFX1 \registers_reg[959][6]  ( .D(n8335), .E(n909), .CK(clk), .Q(
        \registers[959][6] ) );
  EDFFX1 \registers_reg[959][5]  ( .D(n8277), .E(n909), .CK(clk), .Q(
        \registers[959][5] ) );
  EDFFX1 \registers_reg[959][4]  ( .D(n8219), .E(n909), .CK(clk), .Q(
        \registers[959][4] ) );
  EDFFX1 \registers_reg[959][3]  ( .D(n8173), .E(n909), .CK(clk), .Q(
        \registers[959][3] ) );
  EDFFX1 \registers_reg[959][2]  ( .D(n8125), .E(n909), .CK(clk), .Q(
        \registers[959][2] ) );
  EDFFX1 \registers_reg[959][1]  ( .D(n8069), .E(n909), .CK(clk), .Q(
        \registers[959][1] ) );
  EDFFX1 \registers_reg[959][0]  ( .D(n8008), .E(n909), .CK(clk), .Q(
        \registers[959][0] ) );
  EDFFX1 \registers_reg[955][7]  ( .D(n8392), .E(n905), .CK(clk), .Q(
        \registers[955][7] ) );
  EDFFX1 \registers_reg[955][6]  ( .D(n8334), .E(n905), .CK(clk), .Q(
        \registers[955][6] ) );
  EDFFX1 \registers_reg[955][5]  ( .D(n8276), .E(n905), .CK(clk), .Q(
        \registers[955][5] ) );
  EDFFX1 \registers_reg[955][4]  ( .D(n8218), .E(n905), .CK(clk), .Q(
        \registers[955][4] ) );
  EDFFX1 \registers_reg[955][3]  ( .D(n8175), .E(n905), .CK(clk), .Q(
        \registers[955][3] ) );
  EDFFX1 \registers_reg[955][2]  ( .D(n8124), .E(n905), .CK(clk), .Q(
        \registers[955][2] ) );
  EDFFX1 \registers_reg[955][1]  ( .D(n8068), .E(n905), .CK(clk), .Q(
        \registers[955][1] ) );
  EDFFX1 \registers_reg[955][0]  ( .D(n8007), .E(n905), .CK(clk), .Q(
        \registers[955][0] ) );
  EDFFX1 \registers_reg[951][7]  ( .D(n8393), .E(n901), .CK(clk), .Q(
        \registers[951][7] ) );
  EDFFX1 \registers_reg[951][6]  ( .D(n8335), .E(n901), .CK(clk), .Q(
        \registers[951][6] ) );
  EDFFX1 \registers_reg[951][5]  ( .D(n8277), .E(n901), .CK(clk), .Q(
        \registers[951][5] ) );
  EDFFX1 \registers_reg[951][4]  ( .D(n8219), .E(n901), .CK(clk), .Q(
        \registers[951][4] ) );
  EDFFX1 \registers_reg[951][3]  ( .D(n8173), .E(n901), .CK(clk), .Q(
        \registers[951][3] ) );
  EDFFX1 \registers_reg[951][2]  ( .D(n8125), .E(n901), .CK(clk), .Q(
        \registers[951][2] ) );
  EDFFX1 \registers_reg[951][1]  ( .D(n8069), .E(n901), .CK(clk), .Q(
        \registers[951][1] ) );
  EDFFX1 \registers_reg[951][0]  ( .D(n8008), .E(n901), .CK(clk), .Q(
        \registers[951][0] ) );
  EDFFX1 \registers_reg[947][7]  ( .D(n8394), .E(n214), .CK(clk), .Q(
        \registers[947][7] ) );
  EDFFX1 \registers_reg[947][6]  ( .D(n8336), .E(n214), .CK(clk), .Q(
        \registers[947][6] ) );
  EDFFX1 \registers_reg[947][5]  ( .D(n8278), .E(n214), .CK(clk), .Q(
        \registers[947][5] ) );
  EDFFX1 \registers_reg[947][4]  ( .D(n8220), .E(n214), .CK(clk), .Q(
        \registers[947][4] ) );
  EDFFX1 \registers_reg[947][3]  ( .D(n8174), .E(n214), .CK(clk), .Q(
        \registers[947][3] ) );
  EDFFX1 \registers_reg[947][2]  ( .D(n8123), .E(n214), .CK(clk), .Q(
        \registers[947][2] ) );
  EDFFX1 \registers_reg[947][1]  ( .D(n8067), .E(n214), .CK(clk), .Q(
        \registers[947][1] ) );
  EDFFX1 \registers_reg[947][0]  ( .D(n8009), .E(n214), .CK(clk), .Q(
        \registers[947][0] ) );
  EDFFX1 \registers_reg[943][7]  ( .D(n8392), .E(n210), .CK(clk), .Q(
        \registers[943][7] ) );
  EDFFX1 \registers_reg[943][6]  ( .D(n8334), .E(n210), .CK(clk), .Q(
        \registers[943][6] ) );
  EDFFX1 \registers_reg[943][5]  ( .D(n8276), .E(n210), .CK(clk), .Q(
        \registers[943][5] ) );
  EDFFX1 \registers_reg[943][4]  ( .D(n8218), .E(n210), .CK(clk), .Q(
        \registers[943][4] ) );
  EDFFX1 \registers_reg[943][3]  ( .D(n8175), .E(n210), .CK(clk), .Q(
        \registers[943][3] ) );
  EDFFX1 \registers_reg[943][2]  ( .D(n8124), .E(n210), .CK(clk), .Q(
        \registers[943][2] ) );
  EDFFX1 \registers_reg[943][1]  ( .D(n8068), .E(n210), .CK(clk), .Q(
        \registers[943][1] ) );
  EDFFX1 \registers_reg[943][0]  ( .D(n8007), .E(n210), .CK(clk), .Q(
        \registers[943][0] ) );
  EDFFX1 \registers_reg[939][7]  ( .D(n8393), .E(n206), .CK(clk), .Q(
        \registers[939][7] ) );
  EDFFX1 \registers_reg[939][6]  ( .D(n8335), .E(n206), .CK(clk), .Q(
        \registers[939][6] ) );
  EDFFX1 \registers_reg[939][5]  ( .D(n8277), .E(n206), .CK(clk), .Q(
        \registers[939][5] ) );
  EDFFX1 \registers_reg[939][4]  ( .D(n8219), .E(n206), .CK(clk), .Q(
        \registers[939][4] ) );
  EDFFX1 \registers_reg[939][3]  ( .D(n8170), .E(n206), .CK(clk), .Q(
        \registers[939][3] ) );
  EDFFX1 \registers_reg[939][2]  ( .D(n8125), .E(n206), .CK(clk), .Q(
        \registers[939][2] ) );
  EDFFX1 \registers_reg[939][1]  ( .D(n8069), .E(n206), .CK(clk), .Q(
        \registers[939][1] ) );
  EDFFX1 \registers_reg[939][0]  ( .D(n8008), .E(n206), .CK(clk), .Q(
        \registers[939][0] ) );
  EDFFX1 \registers_reg[935][7]  ( .D(n8394), .E(n372), .CK(clk), .Q(
        \registers[935][7] ) );
  EDFFX1 \registers_reg[935][6]  ( .D(n8336), .E(n372), .CK(clk), .Q(
        \registers[935][6] ) );
  EDFFX1 \registers_reg[935][5]  ( .D(n8278), .E(n372), .CK(clk), .Q(
        \registers[935][5] ) );
  EDFFX1 \registers_reg[935][4]  ( .D(n8220), .E(n372), .CK(clk), .Q(
        \registers[935][4] ) );
  EDFFX1 \registers_reg[935][3]  ( .D(n8171), .E(n372), .CK(clk), .Q(
        \registers[935][3] ) );
  EDFFX1 \registers_reg[935][2]  ( .D(n8120), .E(n372), .CK(clk), .Q(
        \registers[935][2] ) );
  EDFFX1 \registers_reg[935][1]  ( .D(n8064), .E(n372), .CK(clk), .Q(
        \registers[935][1] ) );
  EDFFX1 \registers_reg[935][0]  ( .D(n8009), .E(n372), .CK(clk), .Q(
        \registers[935][0] ) );
  EDFFX1 \registers_reg[931][7]  ( .D(n8392), .E(n368), .CK(clk), .Q(
        \registers[931][7] ) );
  EDFFX1 \registers_reg[931][6]  ( .D(n8334), .E(n368), .CK(clk), .Q(
        \registers[931][6] ) );
  EDFFX1 \registers_reg[931][5]  ( .D(n8276), .E(n368), .CK(clk), .Q(
        \registers[931][5] ) );
  EDFFX1 \registers_reg[931][4]  ( .D(n8218), .E(n368), .CK(clk), .Q(
        \registers[931][4] ) );
  EDFFX1 \registers_reg[931][3]  ( .D(n8172), .E(n368), .CK(clk), .Q(
        \registers[931][3] ) );
  EDFFX1 \registers_reg[931][2]  ( .D(n8121), .E(n368), .CK(clk), .Q(
        \registers[931][2] ) );
  EDFFX1 \registers_reg[931][1]  ( .D(n8065), .E(n368), .CK(clk), .Q(
        \registers[931][1] ) );
  EDFFX1 \registers_reg[931][0]  ( .D(n8004), .E(n368), .CK(clk), .Q(
        \registers[931][0] ) );
  EDFFX1 \registers_reg[927][7]  ( .D(n8391), .E(n897), .CK(clk), .Q(
        \registers[927][7] ) );
  EDFFX1 \registers_reg[927][6]  ( .D(n8333), .E(n897), .CK(clk), .Q(
        \registers[927][6] ) );
  EDFFX1 \registers_reg[927][5]  ( .D(n8275), .E(n897), .CK(clk), .Q(
        \registers[927][5] ) );
  EDFFX1 \registers_reg[927][4]  ( .D(n8217), .E(n897), .CK(clk), .Q(
        \registers[927][4] ) );
  EDFFX1 \registers_reg[927][3]  ( .D(n8170), .E(n897), .CK(clk), .Q(
        \registers[927][3] ) );
  EDFFX1 \registers_reg[927][2]  ( .D(n8122), .E(n897), .CK(clk), .Q(
        \registers[927][2] ) );
  EDFFX1 \registers_reg[927][1]  ( .D(n8066), .E(n897), .CK(clk), .Q(
        \registers[927][1] ) );
  EDFFX1 \registers_reg[927][0]  ( .D(n8005), .E(n897), .CK(clk), .Q(
        \registers[927][0] ) );
  EDFFX1 \registers_reg[923][7]  ( .D(n8389), .E(n893), .CK(clk), .Q(
        \registers[923][7] ) );
  EDFFX1 \registers_reg[923][6]  ( .D(n8331), .E(n893), .CK(clk), .Q(
        \registers[923][6] ) );
  EDFFX1 \registers_reg[923][5]  ( .D(n8273), .E(n893), .CK(clk), .Q(
        \registers[923][5] ) );
  EDFFX1 \registers_reg[923][4]  ( .D(n8215), .E(n893), .CK(clk), .Q(
        \registers[923][4] ) );
  EDFFX1 \registers_reg[923][3]  ( .D(n8171), .E(n893), .CK(clk), .Q(
        \registers[923][3] ) );
  EDFFX1 \registers_reg[923][2]  ( .D(n8120), .E(n893), .CK(clk), .Q(
        \registers[923][2] ) );
  EDFFX1 \registers_reg[923][1]  ( .D(n8064), .E(n893), .CK(clk), .Q(
        \registers[923][1] ) );
  EDFFX1 \registers_reg[923][0]  ( .D(n8006), .E(n893), .CK(clk), .Q(
        \registers[923][0] ) );
  EDFFX1 \registers_reg[919][7]  ( .D(n8390), .E(n889), .CK(clk), .Q(
        \registers[919][7] ) );
  EDFFX1 \registers_reg[919][6]  ( .D(n8332), .E(n889), .CK(clk), .Q(
        \registers[919][6] ) );
  EDFFX1 \registers_reg[919][5]  ( .D(n8274), .E(n889), .CK(clk), .Q(
        \registers[919][5] ) );
  EDFFX1 \registers_reg[919][4]  ( .D(n8216), .E(n889), .CK(clk), .Q(
        \registers[919][4] ) );
  EDFFX1 \registers_reg[919][3]  ( .D(n8172), .E(n889), .CK(clk), .Q(
        \registers[919][3] ) );
  EDFFX1 \registers_reg[919][2]  ( .D(n8121), .E(n889), .CK(clk), .Q(
        \registers[919][2] ) );
  EDFFX1 \registers_reg[919][1]  ( .D(n8065), .E(n889), .CK(clk), .Q(
        \registers[919][1] ) );
  EDFFX1 \registers_reg[919][0]  ( .D(n8004), .E(n889), .CK(clk), .Q(
        \registers[919][0] ) );
  EDFFX1 \registers_reg[915][7]  ( .D(n8391), .E(n202), .CK(clk), .Q(
        \registers[915][7] ) );
  EDFFX1 \registers_reg[915][6]  ( .D(n8333), .E(n202), .CK(clk), .Q(
        \registers[915][6] ) );
  EDFFX1 \registers_reg[915][5]  ( .D(n8275), .E(n202), .CK(clk), .Q(
        \registers[915][5] ) );
  EDFFX1 \registers_reg[915][4]  ( .D(n8217), .E(n202), .CK(clk), .Q(
        \registers[915][4] ) );
  EDFFX1 \registers_reg[915][3]  ( .D(n8170), .E(n202), .CK(clk), .Q(
        \registers[915][3] ) );
  EDFFX1 \registers_reg[915][2]  ( .D(n8122), .E(n202), .CK(clk), .Q(
        \registers[915][2] ) );
  EDFFX1 \registers_reg[915][1]  ( .D(n8066), .E(n202), .CK(clk), .Q(
        \registers[915][1] ) );
  EDFFX1 \registers_reg[915][0]  ( .D(n8005), .E(n202), .CK(clk), .Q(
        \registers[915][0] ) );
  EDFFX1 \registers_reg[911][7]  ( .D(n8389), .E(n198), .CK(clk), .Q(
        \registers[911][7] ) );
  EDFFX1 \registers_reg[911][6]  ( .D(n8331), .E(n198), .CK(clk), .Q(
        \registers[911][6] ) );
  EDFFX1 \registers_reg[911][5]  ( .D(n8273), .E(n198), .CK(clk), .Q(
        \registers[911][5] ) );
  EDFFX1 \registers_reg[911][4]  ( .D(n8215), .E(n198), .CK(clk), .Q(
        \registers[911][4] ) );
  EDFFX1 \registers_reg[911][3]  ( .D(n8171), .E(n198), .CK(clk), .Q(
        \registers[911][3] ) );
  EDFFX1 \registers_reg[911][2]  ( .D(n8120), .E(n198), .CK(clk), .Q(
        \registers[911][2] ) );
  EDFFX1 \registers_reg[911][1]  ( .D(n8064), .E(n198), .CK(clk), .Q(
        \registers[911][1] ) );
  EDFFX1 \registers_reg[911][0]  ( .D(n8006), .E(n198), .CK(clk), .Q(
        \registers[911][0] ) );
  EDFFX1 \registers_reg[907][7]  ( .D(n8390), .E(n194), .CK(clk), .Q(
        \registers[907][7] ) );
  EDFFX1 \registers_reg[907][6]  ( .D(n8332), .E(n194), .CK(clk), .Q(
        \registers[907][6] ) );
  EDFFX1 \registers_reg[907][5]  ( .D(n8274), .E(n194), .CK(clk), .Q(
        \registers[907][5] ) );
  EDFFX1 \registers_reg[907][4]  ( .D(n8216), .E(n194), .CK(clk), .Q(
        \registers[907][4] ) );
  EDFFX1 \registers_reg[907][3]  ( .D(n8172), .E(n194), .CK(clk), .Q(
        \registers[907][3] ) );
  EDFFX1 \registers_reg[907][2]  ( .D(n8121), .E(n194), .CK(clk), .Q(
        \registers[907][2] ) );
  EDFFX1 \registers_reg[907][1]  ( .D(n8065), .E(n194), .CK(clk), .Q(
        \registers[907][1] ) );
  EDFFX1 \registers_reg[907][0]  ( .D(n8004), .E(n194), .CK(clk), .Q(
        \registers[907][0] ) );
  EDFFX1 \registers_reg[903][7]  ( .D(n8391), .E(n365), .CK(clk), .Q(
        \registers[903][7] ) );
  EDFFX1 \registers_reg[903][6]  ( .D(n8333), .E(n365), .CK(clk), .Q(
        \registers[903][6] ) );
  EDFFX1 \registers_reg[903][5]  ( .D(n8275), .E(n365), .CK(clk), .Q(
        \registers[903][5] ) );
  EDFFX1 \registers_reg[903][4]  ( .D(n8217), .E(n365), .CK(clk), .Q(
        \registers[903][4] ) );
  EDFFX1 \registers_reg[903][3]  ( .D(n8170), .E(n365), .CK(clk), .Q(
        \registers[903][3] ) );
  EDFFX1 \registers_reg[903][2]  ( .D(n8122), .E(n365), .CK(clk), .Q(
        \registers[903][2] ) );
  EDFFX1 \registers_reg[903][1]  ( .D(n8066), .E(n365), .CK(clk), .Q(
        \registers[903][1] ) );
  EDFFX1 \registers_reg[903][0]  ( .D(n8005), .E(n365), .CK(clk), .Q(
        \registers[903][0] ) );
  EDFFX1 \registers_reg[899][7]  ( .D(n8389), .E(n361), .CK(clk), .Q(
        \registers[899][7] ) );
  EDFFX1 \registers_reg[899][6]  ( .D(n8331), .E(n361), .CK(clk), .Q(
        \registers[899][6] ) );
  EDFFX1 \registers_reg[899][5]  ( .D(n8273), .E(n361), .CK(clk), .Q(
        \registers[899][5] ) );
  EDFFX1 \registers_reg[899][4]  ( .D(n8215), .E(n361), .CK(clk), .Q(
        \registers[899][4] ) );
  EDFFX1 \registers_reg[899][3]  ( .D(n8171), .E(n361), .CK(clk), .Q(
        \registers[899][3] ) );
  EDFFX1 \registers_reg[899][2]  ( .D(n8120), .E(n361), .CK(clk), .Q(
        \registers[899][2] ) );
  EDFFX1 \registers_reg[899][1]  ( .D(n8064), .E(n361), .CK(clk), .Q(
        \registers[899][1] ) );
  EDFFX1 \registers_reg[899][0]  ( .D(n8006), .E(n361), .CK(clk), .Q(
        \registers[899][0] ) );
  EDFFX1 \registers_reg[895][7]  ( .D(n8390), .E(n885), .CK(clk), .Q(
        \registers[895][7] ) );
  EDFFX1 \registers_reg[895][6]  ( .D(n8332), .E(n885), .CK(clk), .Q(
        \registers[895][6] ) );
  EDFFX1 \registers_reg[895][5]  ( .D(n8274), .E(n885), .CK(clk), .Q(
        \registers[895][5] ) );
  EDFFX1 \registers_reg[895][4]  ( .D(n8216), .E(n885), .CK(clk), .Q(
        \registers[895][4] ) );
  EDFFX1 \registers_reg[895][3]  ( .D(n8172), .E(n885), .CK(clk), .Q(
        \registers[895][3] ) );
  EDFFX1 \registers_reg[895][2]  ( .D(n8121), .E(n885), .CK(clk), .Q(
        \registers[895][2] ) );
  EDFFX1 \registers_reg[895][1]  ( .D(n8065), .E(n885), .CK(clk), .Q(
        \registers[895][1] ) );
  EDFFX1 \registers_reg[895][0]  ( .D(n8004), .E(n885), .CK(clk), .Q(
        \registers[895][0] ) );
  EDFFX1 \registers_reg[891][7]  ( .D(n8406), .E(n881), .CK(clk), .Q(
        \registers[891][7] ) );
  EDFFX1 \registers_reg[891][6]  ( .D(n8348), .E(n881), .CK(clk), .Q(
        \registers[891][6] ) );
  EDFFX1 \registers_reg[891][5]  ( .D(n8290), .E(n881), .CK(clk), .Q(
        \registers[891][5] ) );
  EDFFX1 \registers_reg[891][4]  ( .D(n8232), .E(n881), .CK(clk), .Q(
        \registers[891][4] ) );
  EDFFX1 \registers_reg[891][3]  ( .D(n8184), .E(n881), .CK(clk), .Q(
        \registers[891][3] ) );
  EDFFX1 \registers_reg[891][2]  ( .D(n8136), .E(n881), .CK(clk), .Q(
        \registers[891][2] ) );
  EDFFX1 \registers_reg[891][1]  ( .D(n8080), .E(n881), .CK(clk), .Q(
        \registers[891][1] ) );
  EDFFX1 \registers_reg[891][0]  ( .D(n8019), .E(n881), .CK(clk), .Q(
        \registers[891][0] ) );
  EDFFX1 \registers_reg[887][7]  ( .D(n8404), .E(n877), .CK(clk), .Q(
        \registers[887][7] ) );
  EDFFX1 \registers_reg[887][6]  ( .D(n8346), .E(n877), .CK(clk), .Q(
        \registers[887][6] ) );
  EDFFX1 \registers_reg[887][5]  ( .D(n8288), .E(n877), .CK(clk), .Q(
        \registers[887][5] ) );
  EDFFX1 \registers_reg[887][4]  ( .D(n8230), .E(n877), .CK(clk), .Q(
        \registers[887][4] ) );
  EDFFX1 \registers_reg[887][3]  ( .D(n8182), .E(n877), .CK(clk), .Q(
        \registers[887][3] ) );
  EDFFX1 \registers_reg[887][2]  ( .D(n8137), .E(n877), .CK(clk), .Q(
        \registers[887][2] ) );
  EDFFX1 \registers_reg[887][1]  ( .D(n8081), .E(n877), .CK(clk), .Q(
        \registers[887][1] ) );
  EDFFX1 \registers_reg[887][0]  ( .D(n8020), .E(n877), .CK(clk), .Q(
        \registers[887][0] ) );
  EDFFX1 \registers_reg[883][7]  ( .D(n8405), .E(n190), .CK(clk), .Q(
        \registers[883][7] ) );
  EDFFX1 \registers_reg[883][6]  ( .D(n8347), .E(n190), .CK(clk), .Q(
        \registers[883][6] ) );
  EDFFX1 \registers_reg[883][5]  ( .D(n8289), .E(n190), .CK(clk), .Q(
        \registers[883][5] ) );
  EDFFX1 \registers_reg[883][4]  ( .D(n8231), .E(n190), .CK(clk), .Q(
        \registers[883][4] ) );
  EDFFX1 \registers_reg[883][3]  ( .D(n8183), .E(n190), .CK(clk), .Q(
        \registers[883][3] ) );
  EDFFX1 \registers_reg[883][2]  ( .D(n8132), .E(n190), .CK(clk), .Q(
        \registers[883][2] ) );
  EDFFX1 \registers_reg[883][1]  ( .D(n8076), .E(n190), .CK(clk), .Q(
        \registers[883][1] ) );
  EDFFX1 \registers_reg[883][0]  ( .D(n8021), .E(n190), .CK(clk), .Q(
        \registers[883][0] ) );
  EDFFX1 \registers_reg[879][7]  ( .D(n8406), .E(n186), .CK(clk), .Q(
        \registers[879][7] ) );
  EDFFX1 \registers_reg[879][6]  ( .D(n8348), .E(n186), .CK(clk), .Q(
        \registers[879][6] ) );
  EDFFX1 \registers_reg[879][5]  ( .D(n8290), .E(n186), .CK(clk), .Q(
        \registers[879][5] ) );
  EDFFX1 \registers_reg[879][4]  ( .D(n8232), .E(n186), .CK(clk), .Q(
        \registers[879][4] ) );
  EDFFX1 \registers_reg[879][3]  ( .D(n8184), .E(n186), .CK(clk), .Q(
        \registers[879][3] ) );
  EDFFX1 \registers_reg[879][2]  ( .D(n8133), .E(n186), .CK(clk), .Q(
        \registers[879][2] ) );
  EDFFX1 \registers_reg[879][1]  ( .D(n8077), .E(n186), .CK(clk), .Q(
        \registers[879][1] ) );
  EDFFX1 \registers_reg[879][0]  ( .D(n8016), .E(n186), .CK(clk), .Q(
        \registers[879][0] ) );
  EDFFX1 \registers_reg[875][7]  ( .D(n8404), .E(n182), .CK(clk), .Q(
        \registers[875][7] ) );
  EDFFX1 \registers_reg[875][6]  ( .D(n8346), .E(n182), .CK(clk), .Q(
        \registers[875][6] ) );
  EDFFX1 \registers_reg[875][5]  ( .D(n8288), .E(n182), .CK(clk), .Q(
        \registers[875][5] ) );
  EDFFX1 \registers_reg[875][4]  ( .D(n8230), .E(n182), .CK(clk), .Q(
        \registers[875][4] ) );
  EDFFX1 \registers_reg[875][3]  ( .D(n8179), .E(n182), .CK(clk), .Q(
        \registers[875][3] ) );
  EDFFX1 \registers_reg[875][2]  ( .D(n8134), .E(n182), .CK(clk), .Q(
        \registers[875][2] ) );
  EDFFX1 \registers_reg[875][1]  ( .D(n8078), .E(n182), .CK(clk), .Q(
        \registers[875][1] ) );
  EDFFX1 \registers_reg[875][0]  ( .D(n8017), .E(n182), .CK(clk), .Q(
        \registers[875][0] ) );
  EDFFX1 \registers_reg[871][7]  ( .D(n8403), .E(n358), .CK(clk), .Q(
        \registers[871][7] ) );
  EDFFX1 \registers_reg[871][6]  ( .D(n8345), .E(n358), .CK(clk), .Q(
        \registers[871][6] ) );
  EDFFX1 \registers_reg[871][5]  ( .D(n8287), .E(n358), .CK(clk), .Q(
        \registers[871][5] ) );
  EDFFX1 \registers_reg[871][4]  ( .D(n8229), .E(n358), .CK(clk), .Q(
        \registers[871][4] ) );
  EDFFX1 \registers_reg[871][3]  ( .D(n8180), .E(n358), .CK(clk), .Q(
        \registers[871][3] ) );
  EDFFX1 \registers_reg[871][2]  ( .D(n8132), .E(n358), .CK(clk), .Q(
        \registers[871][2] ) );
  EDFFX1 \registers_reg[871][1]  ( .D(n8076), .E(n358), .CK(clk), .Q(
        \registers[871][1] ) );
  EDFFX1 \registers_reg[871][0]  ( .D(n8018), .E(n358), .CK(clk), .Q(
        \registers[871][0] ) );
  EDFFX1 \registers_reg[867][7]  ( .D(n8401), .E(n354), .CK(clk), .Q(
        \registers[867][7] ) );
  EDFFX1 \registers_reg[867][6]  ( .D(n8343), .E(n354), .CK(clk), .Q(
        \registers[867][6] ) );
  EDFFX1 \registers_reg[867][5]  ( .D(n8285), .E(n354), .CK(clk), .Q(
        \registers[867][5] ) );
  EDFFX1 \registers_reg[867][4]  ( .D(n8227), .E(n354), .CK(clk), .Q(
        \registers[867][4] ) );
  EDFFX1 \registers_reg[867][3]  ( .D(n8181), .E(n354), .CK(clk), .Q(
        \registers[867][3] ) );
  EDFFX1 \registers_reg[867][2]  ( .D(n8133), .E(n354), .CK(clk), .Q(
        \registers[867][2] ) );
  EDFFX1 \registers_reg[867][1]  ( .D(n8077), .E(n354), .CK(clk), .Q(
        \registers[867][1] ) );
  EDFFX1 \registers_reg[867][0]  ( .D(n8016), .E(n354), .CK(clk), .Q(
        \registers[867][0] ) );
  EDFFX1 \registers_reg[863][7]  ( .D(n8402), .E(n873), .CK(clk), .Q(
        \registers[863][7] ) );
  EDFFX1 \registers_reg[863][6]  ( .D(n8344), .E(n873), .CK(clk), .Q(
        \registers[863][6] ) );
  EDFFX1 \registers_reg[863][5]  ( .D(n8286), .E(n873), .CK(clk), .Q(
        \registers[863][5] ) );
  EDFFX1 \registers_reg[863][4]  ( .D(n8228), .E(n873), .CK(clk), .Q(
        \registers[863][4] ) );
  EDFFX1 \registers_reg[863][3]  ( .D(n8179), .E(n873), .CK(clk), .Q(
        \registers[863][3] ) );
  EDFFX1 \registers_reg[863][2]  ( .D(n8134), .E(n873), .CK(clk), .Q(
        \registers[863][2] ) );
  EDFFX1 \registers_reg[863][1]  ( .D(n8078), .E(n873), .CK(clk), .Q(
        \registers[863][1] ) );
  EDFFX1 \registers_reg[863][0]  ( .D(n8017), .E(n873), .CK(clk), .Q(
        \registers[863][0] ) );
  EDFFX1 \registers_reg[859][7]  ( .D(n8403), .E(n869), .CK(clk), .Q(
        \registers[859][7] ) );
  EDFFX1 \registers_reg[859][6]  ( .D(n8345), .E(n869), .CK(clk), .Q(
        \registers[859][6] ) );
  EDFFX1 \registers_reg[859][5]  ( .D(n8287), .E(n869), .CK(clk), .Q(
        \registers[859][5] ) );
  EDFFX1 \registers_reg[859][4]  ( .D(n8229), .E(n869), .CK(clk), .Q(
        \registers[859][4] ) );
  EDFFX1 \registers_reg[859][3]  ( .D(n8180), .E(n869), .CK(clk), .Q(
        \registers[859][3] ) );
  EDFFX1 \registers_reg[859][2]  ( .D(n8132), .E(n869), .CK(clk), .Q(
        \registers[859][2] ) );
  EDFFX1 \registers_reg[859][1]  ( .D(n8076), .E(n869), .CK(clk), .Q(
        \registers[859][1] ) );
  EDFFX1 \registers_reg[859][0]  ( .D(n8018), .E(n869), .CK(clk), .Q(
        \registers[859][0] ) );
  EDFFX1 \registers_reg[855][7]  ( .D(n8401), .E(n865), .CK(clk), .Q(
        \registers[855][7] ) );
  EDFFX1 \registers_reg[855][6]  ( .D(n8343), .E(n865), .CK(clk), .Q(
        \registers[855][6] ) );
  EDFFX1 \registers_reg[855][5]  ( .D(n8285), .E(n865), .CK(clk), .Q(
        \registers[855][5] ) );
  EDFFX1 \registers_reg[855][4]  ( .D(n8227), .E(n865), .CK(clk), .Q(
        \registers[855][4] ) );
  EDFFX1 \registers_reg[855][3]  ( .D(n8181), .E(n865), .CK(clk), .Q(
        \registers[855][3] ) );
  EDFFX1 \registers_reg[855][2]  ( .D(n8133), .E(n865), .CK(clk), .Q(
        \registers[855][2] ) );
  EDFFX1 \registers_reg[855][1]  ( .D(n8077), .E(n865), .CK(clk), .Q(
        \registers[855][1] ) );
  EDFFX1 \registers_reg[855][0]  ( .D(n8016), .E(n865), .CK(clk), .Q(
        \registers[855][0] ) );
  EDFFX1 \registers_reg[851][7]  ( .D(n8402), .E(n178), .CK(clk), .Q(
        \registers[851][7] ) );
  EDFFX1 \registers_reg[851][6]  ( .D(n8344), .E(n178), .CK(clk), .Q(
        \registers[851][6] ) );
  EDFFX1 \registers_reg[851][5]  ( .D(n8286), .E(n178), .CK(clk), .Q(
        \registers[851][5] ) );
  EDFFX1 \registers_reg[851][4]  ( .D(n8228), .E(n178), .CK(clk), .Q(
        \registers[851][4] ) );
  EDFFX1 \registers_reg[851][3]  ( .D(n8179), .E(n178), .CK(clk), .Q(
        \registers[851][3] ) );
  EDFFX1 \registers_reg[851][2]  ( .D(n8134), .E(n178), .CK(clk), .Q(
        \registers[851][2] ) );
  EDFFX1 \registers_reg[851][1]  ( .D(n8078), .E(n178), .CK(clk), .Q(
        \registers[851][1] ) );
  EDFFX1 \registers_reg[851][0]  ( .D(n8017), .E(n178), .CK(clk), .Q(
        \registers[851][0] ) );
  EDFFX1 \registers_reg[847][7]  ( .D(n8403), .E(n174), .CK(clk), .Q(
        \registers[847][7] ) );
  EDFFX1 \registers_reg[847][6]  ( .D(n8345), .E(n174), .CK(clk), .Q(
        \registers[847][6] ) );
  EDFFX1 \registers_reg[847][5]  ( .D(n8287), .E(n174), .CK(clk), .Q(
        \registers[847][5] ) );
  EDFFX1 \registers_reg[847][4]  ( .D(n8229), .E(n174), .CK(clk), .Q(
        \registers[847][4] ) );
  EDFFX1 \registers_reg[847][3]  ( .D(n8180), .E(n174), .CK(clk), .Q(
        \registers[847][3] ) );
  EDFFX1 \registers_reg[847][2]  ( .D(n8132), .E(n174), .CK(clk), .Q(
        \registers[847][2] ) );
  EDFFX1 \registers_reg[847][1]  ( .D(n8076), .E(n174), .CK(clk), .Q(
        \registers[847][1] ) );
  EDFFX1 \registers_reg[847][0]  ( .D(n8018), .E(n174), .CK(clk), .Q(
        \registers[847][0] ) );
  EDFFX1 \registers_reg[843][7]  ( .D(n8401), .E(n170), .CK(clk), .Q(
        \registers[843][7] ) );
  EDFFX1 \registers_reg[843][6]  ( .D(n8343), .E(n170), .CK(clk), .Q(
        \registers[843][6] ) );
  EDFFX1 \registers_reg[843][5]  ( .D(n8285), .E(n170), .CK(clk), .Q(
        \registers[843][5] ) );
  EDFFX1 \registers_reg[843][4]  ( .D(n8227), .E(n170), .CK(clk), .Q(
        \registers[843][4] ) );
  EDFFX1 \registers_reg[843][3]  ( .D(n8181), .E(n170), .CK(clk), .Q(
        \registers[843][3] ) );
  EDFFX1 \registers_reg[843][2]  ( .D(n8133), .E(n170), .CK(clk), .Q(
        \registers[843][2] ) );
  EDFFX1 \registers_reg[843][1]  ( .D(n8077), .E(n170), .CK(clk), .Q(
        \registers[843][1] ) );
  EDFFX1 \registers_reg[843][0]  ( .D(n8016), .E(n170), .CK(clk), .Q(
        \registers[843][0] ) );
  EDFFX1 \registers_reg[839][7]  ( .D(n8402), .E(n351), .CK(clk), .Q(
        \registers[839][7] ) );
  EDFFX1 \registers_reg[839][6]  ( .D(n8344), .E(n351), .CK(clk), .Q(
        \registers[839][6] ) );
  EDFFX1 \registers_reg[839][5]  ( .D(n8286), .E(n351), .CK(clk), .Q(
        \registers[839][5] ) );
  EDFFX1 \registers_reg[839][4]  ( .D(n8228), .E(n351), .CK(clk), .Q(
        \registers[839][4] ) );
  EDFFX1 \registers_reg[839][3]  ( .D(n8179), .E(n351), .CK(clk), .Q(
        \registers[839][3] ) );
  EDFFX1 \registers_reg[839][2]  ( .D(n8134), .E(n351), .CK(clk), .Q(
        \registers[839][2] ) );
  EDFFX1 \registers_reg[839][1]  ( .D(n8078), .E(n351), .CK(clk), .Q(
        \registers[839][1] ) );
  EDFFX1 \registers_reg[839][0]  ( .D(n8017), .E(n351), .CK(clk), .Q(
        \registers[839][0] ) );
  EDFFX1 \registers_reg[835][7]  ( .D(n8403), .E(n347), .CK(clk), .Q(
        \registers[835][7] ) );
  EDFFX1 \registers_reg[835][6]  ( .D(n8345), .E(n347), .CK(clk), .Q(
        \registers[835][6] ) );
  EDFFX1 \registers_reg[835][5]  ( .D(n8287), .E(n347), .CK(clk), .Q(
        \registers[835][5] ) );
  EDFFX1 \registers_reg[835][4]  ( .D(n8229), .E(n347), .CK(clk), .Q(
        \registers[835][4] ) );
  EDFFX1 \registers_reg[835][3]  ( .D(n8180), .E(n347), .CK(clk), .Q(
        \registers[835][3] ) );
  EDFFX1 \registers_reg[835][2]  ( .D(n8132), .E(n347), .CK(clk), .Q(
        \registers[835][2] ) );
  EDFFX1 \registers_reg[835][1]  ( .D(n8076), .E(n347), .CK(clk), .Q(
        \registers[835][1] ) );
  EDFFX1 \registers_reg[835][0]  ( .D(n8018), .E(n347), .CK(clk), .Q(
        \registers[835][0] ) );
  EDFFX1 \registers_reg[831][7]  ( .D(n8401), .E(n861), .CK(clk), .Q(
        \registers[831][7] ) );
  EDFFX1 \registers_reg[831][6]  ( .D(n8343), .E(n861), .CK(clk), .Q(
        \registers[831][6] ) );
  EDFFX1 \registers_reg[831][5]  ( .D(n8285), .E(n861), .CK(clk), .Q(
        \registers[831][5] ) );
  EDFFX1 \registers_reg[831][4]  ( .D(n8227), .E(n861), .CK(clk), .Q(
        \registers[831][4] ) );
  EDFFX1 \registers_reg[831][3]  ( .D(n8181), .E(n861), .CK(clk), .Q(
        \registers[831][3] ) );
  EDFFX1 \registers_reg[831][2]  ( .D(n8130), .E(n861), .CK(clk), .Q(
        \registers[831][2] ) );
  EDFFX1 \registers_reg[831][1]  ( .D(n8074), .E(n861), .CK(clk), .Q(
        \registers[831][1] ) );
  EDFFX1 \registers_reg[831][0]  ( .D(n8013), .E(n861), .CK(clk), .Q(
        \registers[831][0] ) );
  EDFFX1 \registers_reg[827][7]  ( .D(n8403), .E(n857), .CK(clk), .Q(
        \registers[827][7] ) );
  EDFFX1 \registers_reg[827][6]  ( .D(n8345), .E(n857), .CK(clk), .Q(
        \registers[827][6] ) );
  EDFFX1 \registers_reg[827][5]  ( .D(n8287), .E(n857), .CK(clk), .Q(
        \registers[827][5] ) );
  EDFFX1 \registers_reg[827][4]  ( .D(n8229), .E(n857), .CK(clk), .Q(
        \registers[827][4] ) );
  EDFFX1 \registers_reg[827][3]  ( .D(n8180), .E(n857), .CK(clk), .Q(
        \registers[827][3] ) );
  EDFFX1 \registers_reg[827][2]  ( .D(n8129), .E(n857), .CK(clk), .Q(
        \registers[827][2] ) );
  EDFFX1 \registers_reg[827][1]  ( .D(n8073), .E(n857), .CK(clk), .Q(
        \registers[827][1] ) );
  EDFFX1 \registers_reg[827][0]  ( .D(n8015), .E(n857), .CK(clk), .Q(
        \registers[827][0] ) );
  EDFFX1 \registers_reg[823][7]  ( .D(n8399), .E(n853), .CK(clk), .Q(
        \registers[823][7] ) );
  EDFFX1 \registers_reg[823][6]  ( .D(n8341), .E(n853), .CK(clk), .Q(
        \registers[823][6] ) );
  EDFFX1 \registers_reg[823][5]  ( .D(n8283), .E(n853), .CK(clk), .Q(
        \registers[823][5] ) );
  EDFFX1 \registers_reg[823][4]  ( .D(n8225), .E(n853), .CK(clk), .Q(
        \registers[823][4] ) );
  EDFFX1 \registers_reg[823][3]  ( .D(n8181), .E(n853), .CK(clk), .Q(
        \registers[823][3] ) );
  EDFFX1 \registers_reg[823][2]  ( .D(n8130), .E(n853), .CK(clk), .Q(
        \registers[823][2] ) );
  EDFFX1 \registers_reg[823][1]  ( .D(n8074), .E(n853), .CK(clk), .Q(
        \registers[823][1] ) );
  EDFFX1 \registers_reg[823][0]  ( .D(n8013), .E(n853), .CK(clk), .Q(
        \registers[823][0] ) );
  EDFFX1 \registers_reg[819][7]  ( .D(n8400), .E(n166), .CK(clk), .Q(
        \registers[819][7] ) );
  EDFFX1 \registers_reg[819][6]  ( .D(n8342), .E(n166), .CK(clk), .Q(
        \registers[819][6] ) );
  EDFFX1 \registers_reg[819][5]  ( .D(n8284), .E(n166), .CK(clk), .Q(
        \registers[819][5] ) );
  EDFFX1 \registers_reg[819][4]  ( .D(n8226), .E(n166), .CK(clk), .Q(
        \registers[819][4] ) );
  EDFFX1 \registers_reg[819][3]  ( .D(n8179), .E(n166), .CK(clk), .Q(
        \registers[819][3] ) );
  EDFFX1 \registers_reg[819][2]  ( .D(n8131), .E(n166), .CK(clk), .Q(
        \registers[819][2] ) );
  EDFFX1 \registers_reg[819][1]  ( .D(n8075), .E(n166), .CK(clk), .Q(
        \registers[819][1] ) );
  EDFFX1 \registers_reg[819][0]  ( .D(n8014), .E(n166), .CK(clk), .Q(
        \registers[819][0] ) );
  EDFFX1 \registers_reg[815][7]  ( .D(n8398), .E(n162), .CK(clk), .Q(
        \registers[815][7] ) );
  EDFFX1 \registers_reg[815][6]  ( .D(n8340), .E(n162), .CK(clk), .Q(
        \registers[815][6] ) );
  EDFFX1 \registers_reg[815][5]  ( .D(n8282), .E(n162), .CK(clk), .Q(
        \registers[815][5] ) );
  EDFFX1 \registers_reg[815][4]  ( .D(n8224), .E(n162), .CK(clk), .Q(
        \registers[815][4] ) );
  EDFFX1 \registers_reg[815][3]  ( .D(n8180), .E(n162), .CK(clk), .Q(
        \registers[815][3] ) );
  EDFFX1 \registers_reg[815][2]  ( .D(n8129), .E(n162), .CK(clk), .Q(
        \registers[815][2] ) );
  EDFFX1 \registers_reg[815][1]  ( .D(n8073), .E(n162), .CK(clk), .Q(
        \registers[815][1] ) );
  EDFFX1 \registers_reg[815][0]  ( .D(n8015), .E(n162), .CK(clk), .Q(
        \registers[815][0] ) );
  EDFFX1 \registers_reg[811][7]  ( .D(n8399), .E(n158), .CK(clk), .Q(
        \registers[811][7] ) );
  EDFFX1 \registers_reg[811][6]  ( .D(n8341), .E(n158), .CK(clk), .Q(
        \registers[811][6] ) );
  EDFFX1 \registers_reg[811][5]  ( .D(n8283), .E(n158), .CK(clk), .Q(
        \registers[811][5] ) );
  EDFFX1 \registers_reg[811][4]  ( .D(n8225), .E(n158), .CK(clk), .Q(
        \registers[811][4] ) );
  EDFFX1 \registers_reg[811][3]  ( .D(n8178), .E(n158), .CK(clk), .Q(
        \registers[811][3] ) );
  EDFFX1 \registers_reg[811][2]  ( .D(n8130), .E(n158), .CK(clk), .Q(
        \registers[811][2] ) );
  EDFFX1 \registers_reg[811][1]  ( .D(n8074), .E(n158), .CK(clk), .Q(
        \registers[811][1] ) );
  EDFFX1 \registers_reg[811][0]  ( .D(n8013), .E(n158), .CK(clk), .Q(
        \registers[811][0] ) );
  EDFFX1 \registers_reg[807][7]  ( .D(n8400), .E(n329), .CK(clk), .Q(
        \registers[807][7] ) );
  EDFFX1 \registers_reg[807][6]  ( .D(n8342), .E(n329), .CK(clk), .Q(
        \registers[807][6] ) );
  EDFFX1 \registers_reg[807][5]  ( .D(n8284), .E(n329), .CK(clk), .Q(
        \registers[807][5] ) );
  EDFFX1 \registers_reg[807][4]  ( .D(n8226), .E(n329), .CK(clk), .Q(
        \registers[807][4] ) );
  EDFFX1 \registers_reg[807][3]  ( .D(n8176), .E(n329), .CK(clk), .Q(
        \registers[807][3] ) );
  EDFFX1 \registers_reg[807][2]  ( .D(n8131), .E(n329), .CK(clk), .Q(
        \registers[807][2] ) );
  EDFFX1 \registers_reg[807][1]  ( .D(n8075), .E(n329), .CK(clk), .Q(
        \registers[807][1] ) );
  EDFFX1 \registers_reg[807][0]  ( .D(n8014), .E(n329), .CK(clk), .Q(
        \registers[807][0] ) );
  EDFFX1 \registers_reg[803][7]  ( .D(n8398), .E(n325), .CK(clk), .Q(
        \registers[803][7] ) );
  EDFFX1 \registers_reg[803][6]  ( .D(n8340), .E(n325), .CK(clk), .Q(
        \registers[803][6] ) );
  EDFFX1 \registers_reg[803][5]  ( .D(n8282), .E(n325), .CK(clk), .Q(
        \registers[803][5] ) );
  EDFFX1 \registers_reg[803][4]  ( .D(n8224), .E(n325), .CK(clk), .Q(
        \registers[803][4] ) );
  EDFFX1 \registers_reg[803][3]  ( .D(n8177), .E(n325), .CK(clk), .Q(
        \registers[803][3] ) );
  EDFFX1 \registers_reg[803][2]  ( .D(n8129), .E(n325), .CK(clk), .Q(
        \registers[803][2] ) );
  EDFFX1 \registers_reg[803][1]  ( .D(n8073), .E(n325), .CK(clk), .Q(
        \registers[803][1] ) );
  EDFFX1 \registers_reg[803][0]  ( .D(n8015), .E(n325), .CK(clk), .Q(
        \registers[803][0] ) );
  EDFFX1 \registers_reg[799][7]  ( .D(n8399), .E(n849), .CK(clk), .Q(
        \registers[799][7] ) );
  EDFFX1 \registers_reg[799][6]  ( .D(n8341), .E(n849), .CK(clk), .Q(
        \registers[799][6] ) );
  EDFFX1 \registers_reg[799][5]  ( .D(n8283), .E(n849), .CK(clk), .Q(
        \registers[799][5] ) );
  EDFFX1 \registers_reg[799][4]  ( .D(n8225), .E(n849), .CK(clk), .Q(
        \registers[799][4] ) );
  EDFFX1 \registers_reg[799][3]  ( .D(n8178), .E(n849), .CK(clk), .Q(
        \registers[799][3] ) );
  EDFFX1 \registers_reg[799][2]  ( .D(n8130), .E(n849), .CK(clk), .Q(
        \registers[799][2] ) );
  EDFFX1 \registers_reg[799][1]  ( .D(n8074), .E(n849), .CK(clk), .Q(
        \registers[799][1] ) );
  EDFFX1 \registers_reg[799][0]  ( .D(n8013), .E(n849), .CK(clk), .Q(
        \registers[799][0] ) );
  EDFFX1 \registers_reg[795][7]  ( .D(n8400), .E(n845), .CK(clk), .Q(
        \registers[795][7] ) );
  EDFFX1 \registers_reg[795][6]  ( .D(n8342), .E(n845), .CK(clk), .Q(
        \registers[795][6] ) );
  EDFFX1 \registers_reg[795][5]  ( .D(n8284), .E(n845), .CK(clk), .Q(
        \registers[795][5] ) );
  EDFFX1 \registers_reg[795][4]  ( .D(n8226), .E(n845), .CK(clk), .Q(
        \registers[795][4] ) );
  EDFFX1 \registers_reg[795][3]  ( .D(n8176), .E(n845), .CK(clk), .Q(
        \registers[795][3] ) );
  EDFFX1 \registers_reg[795][2]  ( .D(n8131), .E(n845), .CK(clk), .Q(
        \registers[795][2] ) );
  EDFFX1 \registers_reg[795][1]  ( .D(n8075), .E(n845), .CK(clk), .Q(
        \registers[795][1] ) );
  EDFFX1 \registers_reg[795][0]  ( .D(n8014), .E(n845), .CK(clk), .Q(
        \registers[795][0] ) );
  EDFFX1 \registers_reg[791][7]  ( .D(n8398), .E(n841), .CK(clk), .Q(
        \registers[791][7] ) );
  EDFFX1 \registers_reg[791][6]  ( .D(n8340), .E(n841), .CK(clk), .Q(
        \registers[791][6] ) );
  EDFFX1 \registers_reg[791][5]  ( .D(n8282), .E(n841), .CK(clk), .Q(
        \registers[791][5] ) );
  EDFFX1 \registers_reg[791][4]  ( .D(n8224), .E(n841), .CK(clk), .Q(
        \registers[791][4] ) );
  EDFFX1 \registers_reg[791][3]  ( .D(n8177), .E(n841), .CK(clk), .Q(
        \registers[791][3] ) );
  EDFFX1 \registers_reg[791][2]  ( .D(n8129), .E(n841), .CK(clk), .Q(
        \registers[791][2] ) );
  EDFFX1 \registers_reg[791][1]  ( .D(n8073), .E(n841), .CK(clk), .Q(
        \registers[791][1] ) );
  EDFFX1 \registers_reg[791][0]  ( .D(n8015), .E(n841), .CK(clk), .Q(
        \registers[791][0] ) );
  EDFFX1 \registers_reg[787][7]  ( .D(n8399), .E(n154), .CK(clk), .Q(
        \registers[787][7] ) );
  EDFFX1 \registers_reg[787][6]  ( .D(n8341), .E(n154), .CK(clk), .Q(
        \registers[787][6] ) );
  EDFFX1 \registers_reg[787][5]  ( .D(n8283), .E(n154), .CK(clk), .Q(
        \registers[787][5] ) );
  EDFFX1 \registers_reg[787][4]  ( .D(n8225), .E(n154), .CK(clk), .Q(
        \registers[787][4] ) );
  EDFFX1 \registers_reg[787][3]  ( .D(n8178), .E(n154), .CK(clk), .Q(
        \registers[787][3] ) );
  EDFFX1 \registers_reg[787][2]  ( .D(n8130), .E(n154), .CK(clk), .Q(
        \registers[787][2] ) );
  EDFFX1 \registers_reg[787][1]  ( .D(n8074), .E(n154), .CK(clk), .Q(
        \registers[787][1] ) );
  EDFFX1 \registers_reg[787][0]  ( .D(n8013), .E(n154), .CK(clk), .Q(
        \registers[787][0] ) );
  EDFFX1 \registers_reg[783][7]  ( .D(n8400), .E(n150), .CK(clk), .Q(
        \registers[783][7] ) );
  EDFFX1 \registers_reg[783][6]  ( .D(n8342), .E(n150), .CK(clk), .Q(
        \registers[783][6] ) );
  EDFFX1 \registers_reg[783][5]  ( .D(n8284), .E(n150), .CK(clk), .Q(
        \registers[783][5] ) );
  EDFFX1 \registers_reg[783][4]  ( .D(n8226), .E(n150), .CK(clk), .Q(
        \registers[783][4] ) );
  EDFFX1 \registers_reg[783][3]  ( .D(n8176), .E(n150), .CK(clk), .Q(
        \registers[783][3] ) );
  EDFFX1 \registers_reg[783][2]  ( .D(n8131), .E(n150), .CK(clk), .Q(
        \registers[783][2] ) );
  EDFFX1 \registers_reg[783][1]  ( .D(n8075), .E(n150), .CK(clk), .Q(
        \registers[783][1] ) );
  EDFFX1 \registers_reg[783][0]  ( .D(n8014), .E(n150), .CK(clk), .Q(
        \registers[783][0] ) );
  EDFFX1 \registers_reg[779][7]  ( .D(n8398), .E(n146), .CK(clk), .Q(
        \registers[779][7] ) );
  EDFFX1 \registers_reg[779][6]  ( .D(n8340), .E(n146), .CK(clk), .Q(
        \registers[779][6] ) );
  EDFFX1 \registers_reg[779][5]  ( .D(n8282), .E(n146), .CK(clk), .Q(
        \registers[779][5] ) );
  EDFFX1 \registers_reg[779][4]  ( .D(n8224), .E(n146), .CK(clk), .Q(
        \registers[779][4] ) );
  EDFFX1 \registers_reg[779][3]  ( .D(n8177), .E(n146), .CK(clk), .Q(
        \registers[779][3] ) );
  EDFFX1 \registers_reg[779][2]  ( .D(n8126), .E(n146), .CK(clk), .Q(
        \registers[779][2] ) );
  EDFFX1 \registers_reg[779][1]  ( .D(n8070), .E(n146), .CK(clk), .Q(
        \registers[779][1] ) );
  EDFFX1 \registers_reg[779][0]  ( .D(n8012), .E(n146), .CK(clk), .Q(
        \registers[779][0] ) );
  EDFFX1 \registers_reg[775][7]  ( .D(n8399), .E(n322), .CK(clk), .Q(
        \registers[775][7] ) );
  EDFFX1 \registers_reg[775][6]  ( .D(n8341), .E(n322), .CK(clk), .Q(
        \registers[775][6] ) );
  EDFFX1 \registers_reg[775][5]  ( .D(n8283), .E(n322), .CK(clk), .Q(
        \registers[775][5] ) );
  EDFFX1 \registers_reg[775][4]  ( .D(n8225), .E(n322), .CK(clk), .Q(
        \registers[775][4] ) );
  EDFFX1 \registers_reg[775][3]  ( .D(n8178), .E(n322), .CK(clk), .Q(
        \registers[775][3] ) );
  EDFFX1 \registers_reg[775][2]  ( .D(n8127), .E(n322), .CK(clk), .Q(
        \registers[775][2] ) );
  EDFFX1 \registers_reg[775][1]  ( .D(n8071), .E(n322), .CK(clk), .Q(
        \registers[775][1] ) );
  EDFFX1 \registers_reg[775][0]  ( .D(n8010), .E(n322), .CK(clk), .Q(
        \registers[775][0] ) );
  EDFFX1 \registers_reg[771][7]  ( .D(n8395), .E(n318), .CK(clk), .Q(
        \registers[771][7] ) );
  EDFFX1 \registers_reg[771][6]  ( .D(n8337), .E(n318), .CK(clk), .Q(
        \registers[771][6] ) );
  EDFFX1 \registers_reg[771][5]  ( .D(n8279), .E(n318), .CK(clk), .Q(
        \registers[771][5] ) );
  EDFFX1 \registers_reg[771][4]  ( .D(n8221), .E(n318), .CK(clk), .Q(
        \registers[771][4] ) );
  EDFFX1 \registers_reg[771][3]  ( .D(n8176), .E(n318), .CK(clk), .Q(
        \registers[771][3] ) );
  EDFFX1 \registers_reg[771][2]  ( .D(n8128), .E(n318), .CK(clk), .Q(
        \registers[771][2] ) );
  EDFFX1 \registers_reg[771][1]  ( .D(n8072), .E(n318), .CK(clk), .Q(
        \registers[771][1] ) );
  EDFFX1 \registers_reg[771][0]  ( .D(n8011), .E(n318), .CK(clk), .Q(
        \registers[771][0] ) );
  EDFFX1 \registers_reg[767][7]  ( .D(n8402), .E(n837), .CK(clk), .Q(
        \registers[767][7] ) );
  EDFFX1 \registers_reg[767][6]  ( .D(n8344), .E(n837), .CK(clk), .Q(
        \registers[767][6] ) );
  EDFFX1 \registers_reg[767][5]  ( .D(n8286), .E(n837), .CK(clk), .Q(
        \registers[767][5] ) );
  EDFFX1 \registers_reg[767][4]  ( .D(n8228), .E(n837), .CK(clk), .Q(
        \registers[767][4] ) );
  EDFFX1 \registers_reg[767][3]  ( .D(n8179), .E(n837), .CK(clk), .Q(
        \registers[767][3] ) );
  EDFFX1 \registers_reg[767][2]  ( .D(n8131), .E(n837), .CK(clk), .Q(
        \registers[767][2] ) );
  EDFFX1 \registers_reg[767][1]  ( .D(n8075), .E(n837), .CK(clk), .Q(
        \registers[767][1] ) );
  EDFFX1 \registers_reg[767][0]  ( .D(n8014), .E(n837), .CK(clk), .Q(
        \registers[767][0] ) );
  EDFFX1 \registers_reg[763][7]  ( .D(n8382), .E(n833), .CK(clk), .Q(
        \registers[763][7] ) );
  EDFFX1 \registers_reg[763][6]  ( .D(n8324), .E(n833), .CK(clk), .Q(
        \registers[763][6] ) );
  EDFFX1 \registers_reg[763][5]  ( .D(n8266), .E(n833), .CK(clk), .Q(
        \registers[763][5] ) );
  EDFFX1 \registers_reg[763][4]  ( .D(n8208), .E(n833), .CK(clk), .Q(
        \registers[763][4] ) );
  EDFFX1 \registers_reg[763][3]  ( .D(n8166), .E(n833), .CK(clk), .Q(
        \registers[763][3] ) );
  EDFFX1 \registers_reg[763][2]  ( .D(n8112), .E(n833), .CK(clk), .Q(
        \registers[763][2] ) );
  EDFFX1 \registers_reg[763][1]  ( .D(n8056), .E(n833), .CK(clk), .Q(
        \registers[763][1] ) );
  EDFFX1 \registers_reg[763][0]  ( .D(n7996), .E(n833), .CK(clk), .Q(
        \registers[763][0] ) );
  EDFFX1 \registers_reg[759][7]  ( .D(n8383), .E(n829), .CK(clk), .Q(
        \registers[759][7] ) );
  EDFFX1 \registers_reg[759][6]  ( .D(n8325), .E(n829), .CK(clk), .Q(
        \registers[759][6] ) );
  EDFFX1 \registers_reg[759][5]  ( .D(n8267), .E(n829), .CK(clk), .Q(
        \registers[759][5] ) );
  EDFFX1 \registers_reg[759][4]  ( .D(n8209), .E(n829), .CK(clk), .Q(
        \registers[759][4] ) );
  EDFFX1 \registers_reg[759][3]  ( .D(n8164), .E(n829), .CK(clk), .Q(
        \registers[759][3] ) );
  EDFFX1 \registers_reg[759][2]  ( .D(n8113), .E(n829), .CK(clk), .Q(
        \registers[759][2] ) );
  EDFFX1 \registers_reg[759][1]  ( .D(n8057), .E(n829), .CK(clk), .Q(
        \registers[759][1] ) );
  EDFFX1 \registers_reg[759][0]  ( .D(n7997), .E(n829), .CK(clk), .Q(
        \registers[759][0] ) );
  EDFFX1 \registers_reg[755][7]  ( .D(n8381), .E(n142), .CK(clk), .Q(
        \registers[755][7] ) );
  EDFFX1 \registers_reg[755][6]  ( .D(n8323), .E(n142), .CK(clk), .Q(
        \registers[755][6] ) );
  EDFFX1 \registers_reg[755][5]  ( .D(n8265), .E(n142), .CK(clk), .Q(
        \registers[755][5] ) );
  EDFFX1 \registers_reg[755][4]  ( .D(n8207), .E(n142), .CK(clk), .Q(
        \registers[755][4] ) );
  EDFFX1 \registers_reg[755][3]  ( .D(n8165), .E(n142), .CK(clk), .Q(
        \registers[755][3] ) );
  EDFFX1 \registers_reg[755][2]  ( .D(n8111), .E(n142), .CK(clk), .Q(
        \registers[755][2] ) );
  EDFFX1 \registers_reg[755][1]  ( .D(n8055), .E(n142), .CK(clk), .Q(
        \registers[755][1] ) );
  EDFFX1 \registers_reg[755][0]  ( .D(n8689), .E(n142), .CK(clk), .Q(
        \registers[755][0] ) );
  EDFFX1 \registers_reg[751][7]  ( .D(n8382), .E(n138), .CK(clk), .Q(
        \registers[751][7] ) );
  EDFFX1 \registers_reg[751][6]  ( .D(n8324), .E(n138), .CK(clk), .Q(
        \registers[751][6] ) );
  EDFFX1 \registers_reg[751][5]  ( .D(n8266), .E(n138), .CK(clk), .Q(
        \registers[751][5] ) );
  EDFFX1 \registers_reg[751][4]  ( .D(n8208), .E(n138), .CK(clk), .Q(
        \registers[751][4] ) );
  EDFFX1 \registers_reg[751][3]  ( .D(n8163), .E(n138), .CK(clk), .Q(
        \registers[751][3] ) );
  EDFFX1 \registers_reg[751][2]  ( .D(n8112), .E(n138), .CK(clk), .Q(
        \registers[751][2] ) );
  EDFFX1 \registers_reg[751][1]  ( .D(n8056), .E(n138), .CK(clk), .Q(
        \registers[751][1] ) );
  EDFFX1 \registers_reg[751][0]  ( .D(n7996), .E(n138), .CK(clk), .Q(
        \registers[751][0] ) );
  EDFFX1 \registers_reg[747][7]  ( .D(n8383), .E(n134), .CK(clk), .Q(
        \registers[747][7] ) );
  EDFFX1 \registers_reg[747][6]  ( .D(n8325), .E(n134), .CK(clk), .Q(
        \registers[747][6] ) );
  EDFFX1 \registers_reg[747][5]  ( .D(n8267), .E(n134), .CK(clk), .Q(
        \registers[747][5] ) );
  EDFFX1 \registers_reg[747][4]  ( .D(n8209), .E(n134), .CK(clk), .Q(
        \registers[747][4] ) );
  EDFFX1 \registers_reg[747][3]  ( .D(n8752), .E(n134), .CK(clk), .Q(
        \registers[747][3] ) );
  EDFFX1 \registers_reg[747][2]  ( .D(n8113), .E(n134), .CK(clk), .Q(
        \registers[747][2] ) );
  EDFFX1 \registers_reg[747][1]  ( .D(n8057), .E(n134), .CK(clk), .Q(
        \registers[747][1] ) );
  EDFFX1 \registers_reg[747][0]  ( .D(n7997), .E(n134), .CK(clk), .Q(
        \registers[747][0] ) );
  EDFFX1 \registers_reg[743][7]  ( .D(n8381), .E(n315), .CK(clk), .Q(
        \registers[743][7] ) );
  EDFFX1 \registers_reg[743][6]  ( .D(n8323), .E(n315), .CK(clk), .Q(
        \registers[743][6] ) );
  EDFFX1 \registers_reg[743][5]  ( .D(n8265), .E(n315), .CK(clk), .Q(
        \registers[743][5] ) );
  EDFFX1 \registers_reg[743][4]  ( .D(n8207), .E(n315), .CK(clk), .Q(
        \registers[743][4] ) );
  EDFFX1 \registers_reg[743][3]  ( .D(n8162), .E(n315), .CK(clk), .Q(
        \registers[743][3] ) );
  EDFFX1 \registers_reg[743][2]  ( .D(n8111), .E(n315), .CK(clk), .Q(
        \registers[743][2] ) );
  EDFFX1 \registers_reg[743][1]  ( .D(n8055), .E(n315), .CK(clk), .Q(
        \registers[743][1] ) );
  EDFFX1 \registers_reg[743][0]  ( .D(n8689), .E(n315), .CK(clk), .Q(
        \registers[743][0] ) );
  EDFFX1 \registers_reg[739][7]  ( .D(n8382), .E(n311), .CK(clk), .Q(
        \registers[739][7] ) );
  EDFFX1 \registers_reg[739][6]  ( .D(n8324), .E(n311), .CK(clk), .Q(
        \registers[739][6] ) );
  EDFFX1 \registers_reg[739][5]  ( .D(n8266), .E(n311), .CK(clk), .Q(
        \registers[739][5] ) );
  EDFFX1 \registers_reg[739][4]  ( .D(n8208), .E(n311), .CK(clk), .Q(
        \registers[739][4] ) );
  EDFFX1 \registers_reg[739][3]  ( .D(n8163), .E(n311), .CK(clk), .Q(
        \registers[739][3] ) );
  EDFFX1 \registers_reg[739][2]  ( .D(n8112), .E(n311), .CK(clk), .Q(
        \registers[739][2] ) );
  EDFFX1 \registers_reg[739][1]  ( .D(n8056), .E(n311), .CK(clk), .Q(
        \registers[739][1] ) );
  EDFFX1 \registers_reg[739][0]  ( .D(n7996), .E(n311), .CK(clk), .Q(
        \registers[739][0] ) );
  EDFFX1 \registers_reg[735][7]  ( .D(n8383), .E(n825), .CK(clk), .Q(
        \registers[735][7] ) );
  EDFFX1 \registers_reg[735][6]  ( .D(n8325), .E(n825), .CK(clk), .Q(
        \registers[735][6] ) );
  EDFFX1 \registers_reg[735][5]  ( .D(n8267), .E(n825), .CK(clk), .Q(
        \registers[735][5] ) );
  EDFFX1 \registers_reg[735][4]  ( .D(n8209), .E(n825), .CK(clk), .Q(
        \registers[735][4] ) );
  EDFFX1 \registers_reg[735][3]  ( .D(n8757), .E(n825), .CK(clk), .Q(
        \registers[735][3] ) );
  EDFFX1 \registers_reg[735][2]  ( .D(n8113), .E(n825), .CK(clk), .Q(
        \registers[735][2] ) );
  EDFFX1 \registers_reg[735][1]  ( .D(n8057), .E(n825), .CK(clk), .Q(
        \registers[735][1] ) );
  EDFFX1 \registers_reg[735][0]  ( .D(n7997), .E(n825), .CK(clk), .Q(
        \registers[735][0] ) );
  EDFFX1 \registers_reg[731][7]  ( .D(n8381), .E(n821), .CK(clk), .Q(
        \registers[731][7] ) );
  EDFFX1 \registers_reg[731][6]  ( .D(n8323), .E(n821), .CK(clk), .Q(
        \registers[731][6] ) );
  EDFFX1 \registers_reg[731][5]  ( .D(n8265), .E(n821), .CK(clk), .Q(
        \registers[731][5] ) );
  EDFFX1 \registers_reg[731][4]  ( .D(n8207), .E(n821), .CK(clk), .Q(
        \registers[731][4] ) );
  EDFFX1 \registers_reg[731][3]  ( .D(n8162), .E(n821), .CK(clk), .Q(
        \registers[731][3] ) );
  EDFFX1 \registers_reg[731][2]  ( .D(n8108), .E(n821), .CK(clk), .Q(
        \registers[731][2] ) );
  EDFFX1 \registers_reg[731][1]  ( .D(n8052), .E(n821), .CK(clk), .Q(
        \registers[731][1] ) );
  EDFFX1 \registers_reg[731][0]  ( .D(n8687), .E(n821), .CK(clk), .Q(
        \registers[731][0] ) );
  EDFFX1 \registers_reg[727][7]  ( .D(n8380), .E(n817), .CK(clk), .Q(
        \registers[727][7] ) );
  EDFFX1 \registers_reg[727][6]  ( .D(n8322), .E(n817), .CK(clk), .Q(
        \registers[727][6] ) );
  EDFFX1 \registers_reg[727][5]  ( .D(n8264), .E(n817), .CK(clk), .Q(
        \registers[727][5] ) );
  EDFFX1 \registers_reg[727][4]  ( .D(n8206), .E(n817), .CK(clk), .Q(
        \registers[727][4] ) );
  EDFFX1 \registers_reg[727][3]  ( .D(n8163), .E(n817), .CK(clk), .Q(
        \registers[727][3] ) );
  EDFFX1 \registers_reg[727][2]  ( .D(n8109), .E(n817), .CK(clk), .Q(
        \registers[727][2] ) );
  EDFFX1 \registers_reg[727][1]  ( .D(n8053), .E(n817), .CK(clk), .Q(
        \registers[727][1] ) );
  EDFFX1 \registers_reg[727][0]  ( .D(n7995), .E(n817), .CK(clk), .Q(
        \registers[727][0] ) );
  EDFFX1 \registers_reg[723][7]  ( .D(n8378), .E(n130), .CK(clk), .Q(
        \registers[723][7] ) );
  EDFFX1 \registers_reg[723][6]  ( .D(n8320), .E(n130), .CK(clk), .Q(
        \registers[723][6] ) );
  EDFFX1 \registers_reg[723][5]  ( .D(n8262), .E(n130), .CK(clk), .Q(
        \registers[723][5] ) );
  EDFFX1 \registers_reg[723][4]  ( .D(n8204), .E(n130), .CK(clk), .Q(
        \registers[723][4] ) );
  EDFFX1 \registers_reg[723][3]  ( .D(n8754), .E(n130), .CK(clk), .Q(
        \registers[723][3] ) );
  EDFFX1 \registers_reg[723][2]  ( .D(n8110), .E(n130), .CK(clk), .Q(
        \registers[723][2] ) );
  EDFFX1 \registers_reg[723][1]  ( .D(n8054), .E(n130), .CK(clk), .Q(
        \registers[723][1] ) );
  EDFFX1 \registers_reg[723][0]  ( .D(n8019), .E(n130), .CK(clk), .Q(
        \registers[723][0] ) );
  EDFFX1 \registers_reg[719][7]  ( .D(n8379), .E(n126), .CK(clk), .Q(
        \registers[719][7] ) );
  EDFFX1 \registers_reg[719][6]  ( .D(n8321), .E(n126), .CK(clk), .Q(
        \registers[719][6] ) );
  EDFFX1 \registers_reg[719][5]  ( .D(n8263), .E(n126), .CK(clk), .Q(
        \registers[719][5] ) );
  EDFFX1 \registers_reg[719][4]  ( .D(n8205), .E(n126), .CK(clk), .Q(
        \registers[719][4] ) );
  EDFFX1 \registers_reg[719][3]  ( .D(n8162), .E(n126), .CK(clk), .Q(
        \registers[719][3] ) );
  EDFFX1 \registers_reg[719][2]  ( .D(n8108), .E(n126), .CK(clk), .Q(
        \registers[719][2] ) );
  EDFFX1 \registers_reg[719][1]  ( .D(n8052), .E(n126), .CK(clk), .Q(
        \registers[719][1] ) );
  EDFFX1 \registers_reg[719][0]  ( .D(n8677), .E(n126), .CK(clk), .Q(
        \registers[719][0] ) );
  EDFFX1 \registers_reg[715][7]  ( .D(n8380), .E(n122), .CK(clk), .Q(
        \registers[715][7] ) );
  EDFFX1 \registers_reg[715][6]  ( .D(n8322), .E(n122), .CK(clk), .Q(
        \registers[715][6] ) );
  EDFFX1 \registers_reg[715][5]  ( .D(n8264), .E(n122), .CK(clk), .Q(
        \registers[715][5] ) );
  EDFFX1 \registers_reg[715][4]  ( .D(n8206), .E(n122), .CK(clk), .Q(
        \registers[715][4] ) );
  EDFFX1 \registers_reg[715][3]  ( .D(n8163), .E(n122), .CK(clk), .Q(
        \registers[715][3] ) );
  EDFFX1 \registers_reg[715][2]  ( .D(n8109), .E(n122), .CK(clk), .Q(
        \registers[715][2] ) );
  EDFFX1 \registers_reg[715][1]  ( .D(n8053), .E(n122), .CK(clk), .Q(
        \registers[715][1] ) );
  EDFFX1 \registers_reg[715][0]  ( .D(n7995), .E(n122), .CK(clk), .Q(
        \registers[715][0] ) );
  EDFFX1 \registers_reg[711][7]  ( .D(n8378), .E(n308), .CK(clk), .Q(
        \registers[711][7] ) );
  EDFFX1 \registers_reg[711][6]  ( .D(n8320), .E(n308), .CK(clk), .Q(
        \registers[711][6] ) );
  EDFFX1 \registers_reg[711][5]  ( .D(n8262), .E(n308), .CK(clk), .Q(
        \registers[711][5] ) );
  EDFFX1 \registers_reg[711][4]  ( .D(n8204), .E(n308), .CK(clk), .Q(
        \registers[711][4] ) );
  EDFFX1 \registers_reg[711][3]  ( .D(n8756), .E(n308), .CK(clk), .Q(
        \registers[711][3] ) );
  EDFFX1 \registers_reg[711][2]  ( .D(n8110), .E(n308), .CK(clk), .Q(
        \registers[711][2] ) );
  EDFFX1 \registers_reg[711][1]  ( .D(n8054), .E(n308), .CK(clk), .Q(
        \registers[711][1] ) );
  EDFFX1 \registers_reg[711][0]  ( .D(n8020), .E(n308), .CK(clk), .Q(
        \registers[711][0] ) );
  EDFFX1 \registers_reg[707][7]  ( .D(n8379), .E(n304), .CK(clk), .Q(
        \registers[707][7] ) );
  EDFFX1 \registers_reg[707][6]  ( .D(n8321), .E(n304), .CK(clk), .Q(
        \registers[707][6] ) );
  EDFFX1 \registers_reg[707][5]  ( .D(n8263), .E(n304), .CK(clk), .Q(
        \registers[707][5] ) );
  EDFFX1 \registers_reg[707][4]  ( .D(n8205), .E(n304), .CK(clk), .Q(
        \registers[707][4] ) );
  EDFFX1 \registers_reg[707][3]  ( .D(n8162), .E(n304), .CK(clk), .Q(
        \registers[707][3] ) );
  EDFFX1 \registers_reg[707][2]  ( .D(n8108), .E(n304), .CK(clk), .Q(
        \registers[707][2] ) );
  EDFFX1 \registers_reg[707][1]  ( .D(n8052), .E(n304), .CK(clk), .Q(
        \registers[707][1] ) );
  EDFFX1 \registers_reg[707][0]  ( .D(n8676), .E(n304), .CK(clk), .Q(
        \registers[707][0] ) );
  EDFFX1 \registers_reg[703][7]  ( .D(n8380), .E(n813), .CK(clk), .Q(
        \registers[703][7] ) );
  EDFFX1 \registers_reg[703][6]  ( .D(n8322), .E(n813), .CK(clk), .Q(
        \registers[703][6] ) );
  EDFFX1 \registers_reg[703][5]  ( .D(n8264), .E(n813), .CK(clk), .Q(
        \registers[703][5] ) );
  EDFFX1 \registers_reg[703][4]  ( .D(n8206), .E(n813), .CK(clk), .Q(
        \registers[703][4] ) );
  EDFFX1 \registers_reg[703][3]  ( .D(n8163), .E(n813), .CK(clk), .Q(
        \registers[703][3] ) );
  EDFFX1 \registers_reg[703][2]  ( .D(n8109), .E(n813), .CK(clk), .Q(
        \registers[703][2] ) );
  EDFFX1 \registers_reg[703][1]  ( .D(n8053), .E(n813), .CK(clk), .Q(
        \registers[703][1] ) );
  EDFFX1 \registers_reg[703][0]  ( .D(n7995), .E(n813), .CK(clk), .Q(
        \registers[703][0] ) );
  EDFFX1 \registers_reg[699][7]  ( .D(n8379), .E(n809), .CK(clk), .Q(
        \registers[699][7] ) );
  EDFFX1 \registers_reg[699][6]  ( .D(n8321), .E(n809), .CK(clk), .Q(
        \registers[699][6] ) );
  EDFFX1 \registers_reg[699][5]  ( .D(n8263), .E(n809), .CK(clk), .Q(
        \registers[699][5] ) );
  EDFFX1 \registers_reg[699][4]  ( .D(n8205), .E(n809), .CK(clk), .Q(
        \registers[699][4] ) );
  EDFFX1 \registers_reg[699][3]  ( .D(n8162), .E(n809), .CK(clk), .Q(
        \registers[699][3] ) );
  EDFFX1 \registers_reg[699][2]  ( .D(n8108), .E(n809), .CK(clk), .Q(
        \registers[699][2] ) );
  EDFFX1 \registers_reg[699][1]  ( .D(n8052), .E(n809), .CK(clk), .Q(
        \registers[699][1] ) );
  EDFFX1 \registers_reg[699][0]  ( .D(n8041), .E(n809), .CK(clk), .Q(
        \registers[699][0] ) );
  EDFFX1 \registers_reg[695][7]  ( .D(n8380), .E(n805), .CK(clk), .Q(
        \registers[695][7] ) );
  EDFFX1 \registers_reg[695][6]  ( .D(n8322), .E(n805), .CK(clk), .Q(
        \registers[695][6] ) );
  EDFFX1 \registers_reg[695][5]  ( .D(n8264), .E(n805), .CK(clk), .Q(
        \registers[695][5] ) );
  EDFFX1 \registers_reg[695][4]  ( .D(n8206), .E(n805), .CK(clk), .Q(
        \registers[695][4] ) );
  EDFFX1 \registers_reg[695][3]  ( .D(n8163), .E(n805), .CK(clk), .Q(
        \registers[695][3] ) );
  EDFFX1 \registers_reg[695][2]  ( .D(n8109), .E(n805), .CK(clk), .Q(
        \registers[695][2] ) );
  EDFFX1 \registers_reg[695][1]  ( .D(n8053), .E(n805), .CK(clk), .Q(
        \registers[695][1] ) );
  EDFFX1 \registers_reg[695][0]  ( .D(n7995), .E(n805), .CK(clk), .Q(
        \registers[695][0] ) );
  EDFFX1 \registers_reg[691][7]  ( .D(n8378), .E(n118), .CK(clk), .Q(
        \registers[691][7] ) );
  EDFFX1 \registers_reg[691][6]  ( .D(n8320), .E(n118), .CK(clk), .Q(
        \registers[691][6] ) );
  EDFFX1 \registers_reg[691][5]  ( .D(n8262), .E(n118), .CK(clk), .Q(
        \registers[691][5] ) );
  EDFFX1 \registers_reg[691][4]  ( .D(n8204), .E(n118), .CK(clk), .Q(
        \registers[691][4] ) );
  EDFFX1 \registers_reg[691][3]  ( .D(n8161), .E(n118), .CK(clk), .Q(
        \registers[691][3] ) );
  EDFFX1 \registers_reg[691][2]  ( .D(n8110), .E(n118), .CK(clk), .Q(
        \registers[691][2] ) );
  EDFFX1 \registers_reg[691][1]  ( .D(n8054), .E(n118), .CK(clk), .Q(
        \registers[691][1] ) );
  EDFFX1 \registers_reg[691][0]  ( .D(n8021), .E(n118), .CK(clk), .Q(
        \registers[691][0] ) );
  EDFFX1 \registers_reg[687][7]  ( .D(n8379), .E(n114), .CK(clk), .Q(
        \registers[687][7] ) );
  EDFFX1 \registers_reg[687][6]  ( .D(n8321), .E(n114), .CK(clk), .Q(
        \registers[687][6] ) );
  EDFFX1 \registers_reg[687][5]  ( .D(n8263), .E(n114), .CK(clk), .Q(
        \registers[687][5] ) );
  EDFFX1 \registers_reg[687][4]  ( .D(n8205), .E(n114), .CK(clk), .Q(
        \registers[687][4] ) );
  EDFFX1 \registers_reg[687][3]  ( .D(n8161), .E(n114), .CK(clk), .Q(
        \registers[687][3] ) );
  EDFFX1 \registers_reg[687][2]  ( .D(n8108), .E(n114), .CK(clk), .Q(
        \registers[687][2] ) );
  EDFFX1 \registers_reg[687][1]  ( .D(n8052), .E(n114), .CK(clk), .Q(
        \registers[687][1] ) );
  EDFFX1 \registers_reg[687][0]  ( .D(n8042), .E(n114), .CK(clk), .Q(
        \registers[687][0] ) );
  EDFFX1 \registers_reg[683][7]  ( .D(n8380), .E(n110), .CK(clk), .Q(
        \registers[683][7] ) );
  EDFFX1 \registers_reg[683][6]  ( .D(n8322), .E(n110), .CK(clk), .Q(
        \registers[683][6] ) );
  EDFFX1 \registers_reg[683][5]  ( .D(n8264), .E(n110), .CK(clk), .Q(
        \registers[683][5] ) );
  EDFFX1 \registers_reg[683][4]  ( .D(n8206), .E(n110), .CK(clk), .Q(
        \registers[683][4] ) );
  EDFFX1 \registers_reg[683][3]  ( .D(n8161), .E(n110), .CK(clk), .Q(
        \registers[683][3] ) );
  EDFFX1 \registers_reg[683][2]  ( .D(n8109), .E(n110), .CK(clk), .Q(
        \registers[683][2] ) );
  EDFFX1 \registers_reg[683][1]  ( .D(n8053), .E(n110), .CK(clk), .Q(
        \registers[683][1] ) );
  EDFFX1 \registers_reg[683][0]  ( .D(n7995), .E(n110), .CK(clk), .Q(
        \registers[683][0] ) );
  EDFFX1 \registers_reg[679][7]  ( .D(n8377), .E(n301), .CK(clk), .Q(
        \registers[679][7] ) );
  EDFFX1 \registers_reg[679][6]  ( .D(n8319), .E(n301), .CK(clk), .Q(
        \registers[679][6] ) );
  EDFFX1 \registers_reg[679][5]  ( .D(n8261), .E(n301), .CK(clk), .Q(
        \registers[679][5] ) );
  EDFFX1 \registers_reg[679][4]  ( .D(n8203), .E(n301), .CK(clk), .Q(
        \registers[679][4] ) );
  EDFFX1 \registers_reg[679][3]  ( .D(n8161), .E(n301), .CK(clk), .Q(
        \registers[679][3] ) );
  EDFFX1 \registers_reg[679][2]  ( .D(n8107), .E(n301), .CK(clk), .Q(
        \registers[679][2] ) );
  EDFFX1 \registers_reg[679][1]  ( .D(n8051), .E(n301), .CK(clk), .Q(
        \registers[679][1] ) );
  EDFFX1 \registers_reg[679][0]  ( .D(n7994), .E(n301), .CK(clk), .Q(
        \registers[679][0] ) );
  EDFFX1 \registers_reg[675][7]  ( .D(n8377), .E(n297), .CK(clk), .Q(
        \registers[675][7] ) );
  EDFFX1 \registers_reg[675][6]  ( .D(n8319), .E(n297), .CK(clk), .Q(
        \registers[675][6] ) );
  EDFFX1 \registers_reg[675][5]  ( .D(n8261), .E(n297), .CK(clk), .Q(
        \registers[675][5] ) );
  EDFFX1 \registers_reg[675][4]  ( .D(n8203), .E(n297), .CK(clk), .Q(
        \registers[675][4] ) );
  EDFFX1 \registers_reg[675][3]  ( .D(n8173), .E(n297), .CK(clk), .Q(
        \registers[675][3] ) );
  EDFFX1 \registers_reg[675][2]  ( .D(n8105), .E(n297), .CK(clk), .Q(
        \registers[675][2] ) );
  EDFFX1 \registers_reg[675][1]  ( .D(n8049), .E(n297), .CK(clk), .Q(
        \registers[675][1] ) );
  EDFFX1 \registers_reg[675][0]  ( .D(n7994), .E(n297), .CK(clk), .Q(
        \registers[675][0] ) );
  EDFFX1 \registers_reg[671][7]  ( .D(n8377), .E(n801), .CK(clk), .Q(
        \registers[671][7] ) );
  EDFFX1 \registers_reg[671][6]  ( .D(n8319), .E(n801), .CK(clk), .Q(
        \registers[671][6] ) );
  EDFFX1 \registers_reg[671][5]  ( .D(n8261), .E(n801), .CK(clk), .Q(
        \registers[671][5] ) );
  EDFFX1 \registers_reg[671][4]  ( .D(n8203), .E(n801), .CK(clk), .Q(
        \registers[671][4] ) );
  EDFFX1 \registers_reg[671][3]  ( .D(n8174), .E(n801), .CK(clk), .Q(
        \registers[671][3] ) );
  EDFFX1 \registers_reg[671][2]  ( .D(n8106), .E(n801), .CK(clk), .Q(
        \registers[671][2] ) );
  EDFFX1 \registers_reg[671][1]  ( .D(n8050), .E(n801), .CK(clk), .Q(
        \registers[671][1] ) );
  EDFFX1 \registers_reg[671][0]  ( .D(n7994), .E(n801), .CK(clk), .Q(
        \registers[671][0] ) );
  EDFFX1 \registers_reg[667][7]  ( .D(n8394), .E(n797), .CK(clk), .Q(
        \registers[667][7] ) );
  EDFFX1 \registers_reg[667][6]  ( .D(n8336), .E(n797), .CK(clk), .Q(
        \registers[667][6] ) );
  EDFFX1 \registers_reg[667][5]  ( .D(n8278), .E(n797), .CK(clk), .Q(
        \registers[667][5] ) );
  EDFFX1 \registers_reg[667][4]  ( .D(n8220), .E(n797), .CK(clk), .Q(
        \registers[667][4] ) );
  EDFFX1 \registers_reg[667][3]  ( .D(n8175), .E(n797), .CK(clk), .Q(
        \registers[667][3] ) );
  EDFFX1 \registers_reg[667][2]  ( .D(n8107), .E(n797), .CK(clk), .Q(
        \registers[667][2] ) );
  EDFFX1 \registers_reg[667][1]  ( .D(n8051), .E(n797), .CK(clk), .Q(
        \registers[667][1] ) );
  EDFFX1 \registers_reg[667][0]  ( .D(n8010), .E(n797), .CK(clk), .Q(
        \registers[667][0] ) );
  EDFFX1 \registers_reg[663][7]  ( .D(n8391), .E(n793), .CK(clk), .Q(
        \registers[663][7] ) );
  EDFFX1 \registers_reg[663][6]  ( .D(n8333), .E(n793), .CK(clk), .Q(
        \registers[663][6] ) );
  EDFFX1 \registers_reg[663][5]  ( .D(n8275), .E(n793), .CK(clk), .Q(
        \registers[663][5] ) );
  EDFFX1 \registers_reg[663][4]  ( .D(n8217), .E(n793), .CK(clk), .Q(
        \registers[663][4] ) );
  EDFFX1 \registers_reg[663][3]  ( .D(n8179), .E(n793), .CK(clk), .Q(
        \registers[663][3] ) );
  EDFFX1 \registers_reg[663][2]  ( .D(n8105), .E(n793), .CK(clk), .Q(
        \registers[663][2] ) );
  EDFFX1 \registers_reg[663][1]  ( .D(n8049), .E(n793), .CK(clk), .Q(
        \registers[663][1] ) );
  EDFFX1 \registers_reg[663][0]  ( .D(n8011), .E(n793), .CK(clk), .Q(
        \registers[663][0] ) );
  EDFFX1 \registers_reg[659][7]  ( .D(n8388), .E(n106), .CK(clk), .Q(
        \registers[659][7] ) );
  EDFFX1 \registers_reg[659][6]  ( .D(n8330), .E(n106), .CK(clk), .Q(
        \registers[659][6] ) );
  EDFFX1 \registers_reg[659][5]  ( .D(n8272), .E(n106), .CK(clk), .Q(
        \registers[659][5] ) );
  EDFFX1 \registers_reg[659][4]  ( .D(n8214), .E(n106), .CK(clk), .Q(
        \registers[659][4] ) );
  EDFFX1 \registers_reg[659][3]  ( .D(n8180), .E(n106), .CK(clk), .Q(
        \registers[659][3] ) );
  EDFFX1 \registers_reg[659][2]  ( .D(n8106), .E(n106), .CK(clk), .Q(
        \registers[659][2] ) );
  EDFFX1 \registers_reg[659][1]  ( .D(n8050), .E(n106), .CK(clk), .Q(
        \registers[659][1] ) );
  EDFFX1 \registers_reg[659][0]  ( .D(n8013), .E(n106), .CK(clk), .Q(
        \registers[659][0] ) );
  EDFFX1 \registers_reg[655][7]  ( .D(n8385), .E(n102), .CK(clk), .Q(
        \registers[655][7] ) );
  EDFFX1 \registers_reg[655][6]  ( .D(n8327), .E(n102), .CK(clk), .Q(
        \registers[655][6] ) );
  EDFFX1 \registers_reg[655][5]  ( .D(n8269), .E(n102), .CK(clk), .Q(
        \registers[655][5] ) );
  EDFFX1 \registers_reg[655][4]  ( .D(n8211), .E(n102), .CK(clk), .Q(
        \registers[655][4] ) );
  EDFFX1 \registers_reg[655][3]  ( .D(n8181), .E(n102), .CK(clk), .Q(
        \registers[655][3] ) );
  EDFFX1 \registers_reg[655][2]  ( .D(n8107), .E(n102), .CK(clk), .Q(
        \registers[655][2] ) );
  EDFFX1 \registers_reg[655][1]  ( .D(n8051), .E(n102), .CK(clk), .Q(
        \registers[655][1] ) );
  EDFFX1 \registers_reg[655][0]  ( .D(n8015), .E(n102), .CK(clk), .Q(
        \registers[655][0] ) );
  EDFFX1 \registers_reg[651][7]  ( .D(n8387), .E(n98), .CK(clk), .Q(
        \registers[651][7] ) );
  EDFFX1 \registers_reg[651][6]  ( .D(n8329), .E(n98), .CK(clk), .Q(
        \registers[651][6] ) );
  EDFFX1 \registers_reg[651][5]  ( .D(n8271), .E(n98), .CK(clk), .Q(
        \registers[651][5] ) );
  EDFFX1 \registers_reg[651][4]  ( .D(n8213), .E(n98), .CK(clk), .Q(
        \registers[651][4] ) );
  EDFFX1 \registers_reg[651][3]  ( .D(n8177), .E(n98), .CK(clk), .Q(
        \registers[651][3] ) );
  EDFFX1 \registers_reg[651][2]  ( .D(n8105), .E(n98), .CK(clk), .Q(
        \registers[651][2] ) );
  EDFFX1 \registers_reg[651][1]  ( .D(n8049), .E(n98), .CK(clk), .Q(
        \registers[651][1] ) );
  EDFFX1 \registers_reg[651][0]  ( .D(n8014), .E(n98), .CK(clk), .Q(
        \registers[651][0] ) );
  EDFFX1 \registers_reg[647][7]  ( .D(n8384), .E(n294), .CK(clk), .Q(
        \registers[647][7] ) );
  EDFFX1 \registers_reg[647][6]  ( .D(n8326), .E(n294), .CK(clk), .Q(
        \registers[647][6] ) );
  EDFFX1 \registers_reg[647][5]  ( .D(n8268), .E(n294), .CK(clk), .Q(
        \registers[647][5] ) );
  EDFFX1 \registers_reg[647][4]  ( .D(n8210), .E(n294), .CK(clk), .Q(
        \registers[647][4] ) );
  EDFFX1 \registers_reg[647][3]  ( .D(n8178), .E(n294), .CK(clk), .Q(
        \registers[647][3] ) );
  EDFFX1 \registers_reg[647][2]  ( .D(n8106), .E(n294), .CK(clk), .Q(
        \registers[647][2] ) );
  EDFFX1 \registers_reg[647][1]  ( .D(n8050), .E(n294), .CK(clk), .Q(
        \registers[647][1] ) );
  EDFFX1 \registers_reg[647][0]  ( .D(n8007), .E(n294), .CK(clk), .Q(
        \registers[647][0] ) );
  EDFFX1 \registers_reg[643][7]  ( .D(n8421), .E(n290), .CK(clk), .Q(
        \registers[643][7] ) );
  EDFFX1 \registers_reg[643][6]  ( .D(n8363), .E(n290), .CK(clk), .Q(
        \registers[643][6] ) );
  EDFFX1 \registers_reg[643][5]  ( .D(n8305), .E(n290), .CK(clk), .Q(
        \registers[643][5] ) );
  EDFFX1 \registers_reg[643][4]  ( .D(n8247), .E(n290), .CK(clk), .Q(
        \registers[643][4] ) );
  EDFFX1 \registers_reg[643][3]  ( .D(n8176), .E(n290), .CK(clk), .Q(
        \registers[643][3] ) );
  EDFFX1 \registers_reg[643][2]  ( .D(n8107), .E(n290), .CK(clk), .Q(
        \registers[643][2] ) );
  EDFFX1 \registers_reg[643][1]  ( .D(n8051), .E(n290), .CK(clk), .Q(
        \registers[643][1] ) );
  EDFFX1 \registers_reg[643][0]  ( .D(n8008), .E(n290), .CK(clk), .Q(
        \registers[643][0] ) );
  EDFFX1 \registers_reg[639][7]  ( .D(n8389), .E(n789), .CK(clk), .Q(
        \registers[639][7] ) );
  EDFFX1 \registers_reg[639][6]  ( .D(n8331), .E(n789), .CK(clk), .Q(
        \registers[639][6] ) );
  EDFFX1 \registers_reg[639][5]  ( .D(n8273), .E(n789), .CK(clk), .Q(
        \registers[639][5] ) );
  EDFFX1 \registers_reg[639][4]  ( .D(n8215), .E(n789), .CK(clk), .Q(
        \registers[639][4] ) );
  EDFFX1 \registers_reg[639][3]  ( .D(n8171), .E(n789), .CK(clk), .Q(
        \registers[639][3] ) );
  EDFFX1 \registers_reg[639][2]  ( .D(n8120), .E(n789), .CK(clk), .Q(
        \registers[639][2] ) );
  EDFFX1 \registers_reg[639][1]  ( .D(n8064), .E(n789), .CK(clk), .Q(
        \registers[639][1] ) );
  EDFFX1 \registers_reg[639][0]  ( .D(n8016), .E(n789), .CK(clk), .Q(
        \registers[639][0] ) );
  EDFFX1 \registers_reg[635][7]  ( .D(n8390), .E(n785), .CK(clk), .Q(
        \registers[635][7] ) );
  EDFFX1 \registers_reg[635][6]  ( .D(n8332), .E(n785), .CK(clk), .Q(
        \registers[635][6] ) );
  EDFFX1 \registers_reg[635][5]  ( .D(n8274), .E(n785), .CK(clk), .Q(
        \registers[635][5] ) );
  EDFFX1 \registers_reg[635][4]  ( .D(n8216), .E(n785), .CK(clk), .Q(
        \registers[635][4] ) );
  EDFFX1 \registers_reg[635][3]  ( .D(n8172), .E(n785), .CK(clk), .Q(
        \registers[635][3] ) );
  EDFFX1 \registers_reg[635][2]  ( .D(n8121), .E(n785), .CK(clk), .Q(
        \registers[635][2] ) );
  EDFFX1 \registers_reg[635][1]  ( .D(n8065), .E(n785), .CK(clk), .Q(
        \registers[635][1] ) );
  EDFFX1 \registers_reg[635][0]  ( .D(n8006), .E(n785), .CK(clk), .Q(
        \registers[635][0] ) );
  EDFFX1 \registers_reg[631][7]  ( .D(n8391), .E(n781), .CK(clk), .Q(
        \registers[631][7] ) );
  EDFFX1 \registers_reg[631][6]  ( .D(n8333), .E(n781), .CK(clk), .Q(
        \registers[631][6] ) );
  EDFFX1 \registers_reg[631][5]  ( .D(n8275), .E(n781), .CK(clk), .Q(
        \registers[631][5] ) );
  EDFFX1 \registers_reg[631][4]  ( .D(n8217), .E(n781), .CK(clk), .Q(
        \registers[631][4] ) );
  EDFFX1 \registers_reg[631][3]  ( .D(n8170), .E(n781), .CK(clk), .Q(
        \registers[631][3] ) );
  EDFFX1 \registers_reg[631][2]  ( .D(n8122), .E(n781), .CK(clk), .Q(
        \registers[631][2] ) );
  EDFFX1 \registers_reg[631][1]  ( .D(n8066), .E(n781), .CK(clk), .Q(
        \registers[631][1] ) );
  EDFFX1 \registers_reg[631][0]  ( .D(n8004), .E(n781), .CK(clk), .Q(
        \registers[631][0] ) );
  EDFFX1 \registers_reg[627][7]  ( .D(n8389), .E(n94), .CK(clk), .Q(
        \registers[627][7] ) );
  EDFFX1 \registers_reg[627][6]  ( .D(n8331), .E(n94), .CK(clk), .Q(
        \registers[627][6] ) );
  EDFFX1 \registers_reg[627][5]  ( .D(n8273), .E(n94), .CK(clk), .Q(
        \registers[627][5] ) );
  EDFFX1 \registers_reg[627][4]  ( .D(n8215), .E(n94), .CK(clk), .Q(
        \registers[627][4] ) );
  EDFFX1 \registers_reg[627][3]  ( .D(n8171), .E(n94), .CK(clk), .Q(
        \registers[627][3] ) );
  EDFFX1 \registers_reg[627][2]  ( .D(n8117), .E(n94), .CK(clk), .Q(
        \registers[627][2] ) );
  EDFFX1 \registers_reg[627][1]  ( .D(n8061), .E(n94), .CK(clk), .Q(
        \registers[627][1] ) );
  EDFFX1 \registers_reg[627][0]  ( .D(n8002), .E(n94), .CK(clk), .Q(
        \registers[627][0] ) );
  EDFFX1 \registers_reg[623][7]  ( .D(n8388), .E(n90), .CK(clk), .Q(
        \registers[623][7] ) );
  EDFFX1 \registers_reg[623][6]  ( .D(n8330), .E(n90), .CK(clk), .Q(
        \registers[623][6] ) );
  EDFFX1 \registers_reg[623][5]  ( .D(n8272), .E(n90), .CK(clk), .Q(
        \registers[623][5] ) );
  EDFFX1 \registers_reg[623][4]  ( .D(n8214), .E(n90), .CK(clk), .Q(
        \registers[623][4] ) );
  EDFFX1 \registers_reg[623][3]  ( .D(n8169), .E(n90), .CK(clk), .Q(
        \registers[623][3] ) );
  EDFFX1 \registers_reg[623][2]  ( .D(n8118), .E(n90), .CK(clk), .Q(
        \registers[623][2] ) );
  EDFFX1 \registers_reg[623][1]  ( .D(n8062), .E(n90), .CK(clk), .Q(
        \registers[623][1] ) );
  EDFFX1 \registers_reg[623][0]  ( .D(n8003), .E(n90), .CK(clk), .Q(
        \registers[623][0] ) );
  EDFFX1 \registers_reg[619][7]  ( .D(n8386), .E(n86), .CK(clk), .Q(
        \registers[619][7] ) );
  EDFFX1 \registers_reg[619][6]  ( .D(n8328), .E(n86), .CK(clk), .Q(
        \registers[619][6] ) );
  EDFFX1 \registers_reg[619][5]  ( .D(n8270), .E(n86), .CK(clk), .Q(
        \registers[619][5] ) );
  EDFFX1 \registers_reg[619][4]  ( .D(n8212), .E(n86), .CK(clk), .Q(
        \registers[619][4] ) );
  EDFFX1 \registers_reg[619][3]  ( .D(n8167), .E(n86), .CK(clk), .Q(
        \registers[619][3] ) );
  EDFFX1 \registers_reg[619][2]  ( .D(n8119), .E(n86), .CK(clk), .Q(
        \registers[619][2] ) );
  EDFFX1 \registers_reg[619][1]  ( .D(n8063), .E(n86), .CK(clk), .Q(
        \registers[619][1] ) );
  EDFFX1 \registers_reg[619][0]  ( .D(n8001), .E(n86), .CK(clk), .Q(
        \registers[619][0] ) );
  EDFFX1 \registers_reg[615][7]  ( .D(n8387), .E(n287), .CK(clk), .Q(
        \registers[615][7] ) );
  EDFFX1 \registers_reg[615][6]  ( .D(n8329), .E(n287), .CK(clk), .Q(
        \registers[615][6] ) );
  EDFFX1 \registers_reg[615][5]  ( .D(n8271), .E(n287), .CK(clk), .Q(
        \registers[615][5] ) );
  EDFFX1 \registers_reg[615][4]  ( .D(n8213), .E(n287), .CK(clk), .Q(
        \registers[615][4] ) );
  EDFFX1 \registers_reg[615][3]  ( .D(n8168), .E(n287), .CK(clk), .Q(
        \registers[615][3] ) );
  EDFFX1 \registers_reg[615][2]  ( .D(n8117), .E(n287), .CK(clk), .Q(
        \registers[615][2] ) );
  EDFFX1 \registers_reg[615][1]  ( .D(n8061), .E(n287), .CK(clk), .Q(
        \registers[615][1] ) );
  EDFFX1 \registers_reg[615][0]  ( .D(n8002), .E(n287), .CK(clk), .Q(
        \registers[615][0] ) );
  EDFFX1 \registers_reg[611][7]  ( .D(n8388), .E(n283), .CK(clk), .Q(
        \registers[611][7] ) );
  EDFFX1 \registers_reg[611][6]  ( .D(n8330), .E(n283), .CK(clk), .Q(
        \registers[611][6] ) );
  EDFFX1 \registers_reg[611][5]  ( .D(n8272), .E(n283), .CK(clk), .Q(
        \registers[611][5] ) );
  EDFFX1 \registers_reg[611][4]  ( .D(n8214), .E(n283), .CK(clk), .Q(
        \registers[611][4] ) );
  EDFFX1 \registers_reg[611][3]  ( .D(n8169), .E(n283), .CK(clk), .Q(
        \registers[611][3] ) );
  EDFFX1 \registers_reg[611][2]  ( .D(n8118), .E(n283), .CK(clk), .Q(
        \registers[611][2] ) );
  EDFFX1 \registers_reg[611][1]  ( .D(n8062), .E(n283), .CK(clk), .Q(
        \registers[611][1] ) );
  EDFFX1 \registers_reg[611][0]  ( .D(n8003), .E(n283), .CK(clk), .Q(
        \registers[611][0] ) );
  EDFFX1 \registers_reg[607][7]  ( .D(n8386), .E(n777), .CK(clk), .Q(
        \registers[607][7] ) );
  EDFFX1 \registers_reg[607][6]  ( .D(n8328), .E(n777), .CK(clk), .Q(
        \registers[607][6] ) );
  EDFFX1 \registers_reg[607][5]  ( .D(n8270), .E(n777), .CK(clk), .Q(
        \registers[607][5] ) );
  EDFFX1 \registers_reg[607][4]  ( .D(n8212), .E(n777), .CK(clk), .Q(
        \registers[607][4] ) );
  EDFFX1 \registers_reg[607][3]  ( .D(n8167), .E(n777), .CK(clk), .Q(
        \registers[607][3] ) );
  EDFFX1 \registers_reg[607][2]  ( .D(n8119), .E(n777), .CK(clk), .Q(
        \registers[607][2] ) );
  EDFFX1 \registers_reg[607][1]  ( .D(n8063), .E(n777), .CK(clk), .Q(
        \registers[607][1] ) );
  EDFFX1 \registers_reg[607][0]  ( .D(n8001), .E(n777), .CK(clk), .Q(
        \registers[607][0] ) );
  EDFFX1 \registers_reg[603][7]  ( .D(n8387), .E(n773), .CK(clk), .Q(
        \registers[603][7] ) );
  EDFFX1 \registers_reg[603][6]  ( .D(n8329), .E(n773), .CK(clk), .Q(
        \registers[603][6] ) );
  EDFFX1 \registers_reg[603][5]  ( .D(n8271), .E(n773), .CK(clk), .Q(
        \registers[603][5] ) );
  EDFFX1 \registers_reg[603][4]  ( .D(n8213), .E(n773), .CK(clk), .Q(
        \registers[603][4] ) );
  EDFFX1 \registers_reg[603][3]  ( .D(n8168), .E(n773), .CK(clk), .Q(
        \registers[603][3] ) );
  EDFFX1 \registers_reg[603][2]  ( .D(n8117), .E(n773), .CK(clk), .Q(
        \registers[603][2] ) );
  EDFFX1 \registers_reg[603][1]  ( .D(n8061), .E(n773), .CK(clk), .Q(
        \registers[603][1] ) );
  EDFFX1 \registers_reg[603][0]  ( .D(n8002), .E(n773), .CK(clk), .Q(
        \registers[603][0] ) );
  EDFFX1 \registers_reg[599][7]  ( .D(n8388), .E(n769), .CK(clk), .Q(
        \registers[599][7] ) );
  EDFFX1 \registers_reg[599][6]  ( .D(n8330), .E(n769), .CK(clk), .Q(
        \registers[599][6] ) );
  EDFFX1 \registers_reg[599][5]  ( .D(n8272), .E(n769), .CK(clk), .Q(
        \registers[599][5] ) );
  EDFFX1 \registers_reg[599][4]  ( .D(n8214), .E(n769), .CK(clk), .Q(
        \registers[599][4] ) );
  EDFFX1 \registers_reg[599][3]  ( .D(n8169), .E(n769), .CK(clk), .Q(
        \registers[599][3] ) );
  EDFFX1 \registers_reg[599][2]  ( .D(n8118), .E(n769), .CK(clk), .Q(
        \registers[599][2] ) );
  EDFFX1 \registers_reg[599][1]  ( .D(n8062), .E(n769), .CK(clk), .Q(
        \registers[599][1] ) );
  EDFFX1 \registers_reg[599][0]  ( .D(n8003), .E(n769), .CK(clk), .Q(
        \registers[599][0] ) );
  EDFFX1 \registers_reg[595][7]  ( .D(n8386), .E(n82), .CK(clk), .Q(
        \registers[595][7] ) );
  EDFFX1 \registers_reg[595][6]  ( .D(n8328), .E(n82), .CK(clk), .Q(
        \registers[595][6] ) );
  EDFFX1 \registers_reg[595][5]  ( .D(n8270), .E(n82), .CK(clk), .Q(
        \registers[595][5] ) );
  EDFFX1 \registers_reg[595][4]  ( .D(n8212), .E(n82), .CK(clk), .Q(
        \registers[595][4] ) );
  EDFFX1 \registers_reg[595][3]  ( .D(n8167), .E(n82), .CK(clk), .Q(
        \registers[595][3] ) );
  EDFFX1 \registers_reg[595][2]  ( .D(n8119), .E(n82), .CK(clk), .Q(
        \registers[595][2] ) );
  EDFFX1 \registers_reg[595][1]  ( .D(n8063), .E(n82), .CK(clk), .Q(
        \registers[595][1] ) );
  EDFFX1 \registers_reg[595][0]  ( .D(n8001), .E(n82), .CK(clk), .Q(
        \registers[595][0] ) );
  EDFFX1 \registers_reg[591][7]  ( .D(n8387), .E(n78), .CK(clk), .Q(
        \registers[591][7] ) );
  EDFFX1 \registers_reg[591][6]  ( .D(n8329), .E(n78), .CK(clk), .Q(
        \registers[591][6] ) );
  EDFFX1 \registers_reg[591][5]  ( .D(n8271), .E(n78), .CK(clk), .Q(
        \registers[591][5] ) );
  EDFFX1 \registers_reg[591][4]  ( .D(n8213), .E(n78), .CK(clk), .Q(
        \registers[591][4] ) );
  EDFFX1 \registers_reg[591][3]  ( .D(n8168), .E(n78), .CK(clk), .Q(
        \registers[591][3] ) );
  EDFFX1 \registers_reg[591][2]  ( .D(n8117), .E(n78), .CK(clk), .Q(
        \registers[591][2] ) );
  EDFFX1 \registers_reg[591][1]  ( .D(n8061), .E(n78), .CK(clk), .Q(
        \registers[591][1] ) );
  EDFFX1 \registers_reg[591][0]  ( .D(n8002), .E(n78), .CK(clk), .Q(
        \registers[591][0] ) );
  EDFFX1 \registers_reg[587][7]  ( .D(n8388), .E(n74), .CK(clk), .Q(
        \registers[587][7] ) );
  EDFFX1 \registers_reg[587][6]  ( .D(n8330), .E(n74), .CK(clk), .Q(
        \registers[587][6] ) );
  EDFFX1 \registers_reg[587][5]  ( .D(n8272), .E(n74), .CK(clk), .Q(
        \registers[587][5] ) );
  EDFFX1 \registers_reg[587][4]  ( .D(n8214), .E(n74), .CK(clk), .Q(
        \registers[587][4] ) );
  EDFFX1 \registers_reg[587][3]  ( .D(n8169), .E(n74), .CK(clk), .Q(
        \registers[587][3] ) );
  EDFFX1 \registers_reg[587][2]  ( .D(n8118), .E(n74), .CK(clk), .Q(
        \registers[587][2] ) );
  EDFFX1 \registers_reg[587][1]  ( .D(n8062), .E(n74), .CK(clk), .Q(
        \registers[587][1] ) );
  EDFFX1 \registers_reg[587][0]  ( .D(n8003), .E(n74), .CK(clk), .Q(
        \registers[587][0] ) );
  EDFFX1 \registers_reg[583][7]  ( .D(n8386), .E(n280), .CK(clk), .Q(
        \registers[583][7] ) );
  EDFFX1 \registers_reg[583][6]  ( .D(n8328), .E(n280), .CK(clk), .Q(
        \registers[583][6] ) );
  EDFFX1 \registers_reg[583][5]  ( .D(n8270), .E(n280), .CK(clk), .Q(
        \registers[583][5] ) );
  EDFFX1 \registers_reg[583][4]  ( .D(n8212), .E(n280), .CK(clk), .Q(
        \registers[583][4] ) );
  EDFFX1 \registers_reg[583][3]  ( .D(n8167), .E(n280), .CK(clk), .Q(
        \registers[583][3] ) );
  EDFFX1 \registers_reg[583][2]  ( .D(n8119), .E(n280), .CK(clk), .Q(
        \registers[583][2] ) );
  EDFFX1 \registers_reg[583][1]  ( .D(n8063), .E(n280), .CK(clk), .Q(
        \registers[583][1] ) );
  EDFFX1 \registers_reg[583][0]  ( .D(n8001), .E(n280), .CK(clk), .Q(
        \registers[583][0] ) );
  EDFFX1 \registers_reg[579][7]  ( .D(n8387), .E(n276), .CK(clk), .Q(
        \registers[579][7] ) );
  EDFFX1 \registers_reg[579][6]  ( .D(n8329), .E(n276), .CK(clk), .Q(
        \registers[579][6] ) );
  EDFFX1 \registers_reg[579][5]  ( .D(n8271), .E(n276), .CK(clk), .Q(
        \registers[579][5] ) );
  EDFFX1 \registers_reg[579][4]  ( .D(n8213), .E(n276), .CK(clk), .Q(
        \registers[579][4] ) );
  EDFFX1 \registers_reg[579][3]  ( .D(n8168), .E(n276), .CK(clk), .Q(
        \registers[579][3] ) );
  EDFFX1 \registers_reg[579][2]  ( .D(n8114), .E(n276), .CK(clk), .Q(
        \registers[579][2] ) );
  EDFFX1 \registers_reg[579][1]  ( .D(n8058), .E(n276), .CK(clk), .Q(
        \registers[579][1] ) );
  EDFFX1 \registers_reg[579][0]  ( .D(n8002), .E(n276), .CK(clk), .Q(
        \registers[579][0] ) );
  EDFFX1 \registers_reg[575][7]  ( .D(n8422), .E(n765), .CK(clk), .Q(
        \registers[575][7] ) );
  EDFFX1 \registers_reg[575][6]  ( .D(n8364), .E(n765), .CK(clk), .Q(
        \registers[575][6] ) );
  EDFFX1 \registers_reg[575][5]  ( .D(n8306), .E(n765), .CK(clk), .Q(
        \registers[575][5] ) );
  EDFFX1 \registers_reg[575][4]  ( .D(n8248), .E(n765), .CK(clk), .Q(
        \registers[575][4] ) );
  EDFFX1 \registers_reg[575][3]  ( .D(n8167), .E(n765), .CK(clk), .Q(
        \registers[575][3] ) );
  EDFFX1 \registers_reg[575][2]  ( .D(n8116), .E(n765), .CK(clk), .Q(
        \registers[575][2] ) );
  EDFFX1 \registers_reg[575][1]  ( .D(n8060), .E(n765), .CK(clk), .Q(
        \registers[575][1] ) );
  EDFFX1 \registers_reg[575][0]  ( .D(n7998), .E(n765), .CK(clk), .Q(
        \registers[575][0] ) );
  EDFFX1 \registers_reg[571][7]  ( .D(n8385), .E(n761), .CK(clk), .Q(
        \registers[571][7] ) );
  EDFFX1 \registers_reg[571][6]  ( .D(n8327), .E(n761), .CK(clk), .Q(
        \registers[571][6] ) );
  EDFFX1 \registers_reg[571][5]  ( .D(n8269), .E(n761), .CK(clk), .Q(
        \registers[571][5] ) );
  EDFFX1 \registers_reg[571][4]  ( .D(n8211), .E(n761), .CK(clk), .Q(
        \registers[571][4] ) );
  EDFFX1 \registers_reg[571][3]  ( .D(n8168), .E(n761), .CK(clk), .Q(
        \registers[571][3] ) );
  EDFFX1 \registers_reg[571][2]  ( .D(n8114), .E(n761), .CK(clk), .Q(
        \registers[571][2] ) );
  EDFFX1 \registers_reg[571][1]  ( .D(n8058), .E(n761), .CK(clk), .Q(
        \registers[571][1] ) );
  EDFFX1 \registers_reg[571][0]  ( .D(n7999), .E(n761), .CK(clk), .Q(
        \registers[571][0] ) );
  EDFFX1 \registers_reg[567][7]  ( .D(n8384), .E(n757), .CK(clk), .Q(
        \registers[567][7] ) );
  EDFFX1 \registers_reg[567][6]  ( .D(n8326), .E(n757), .CK(clk), .Q(
        \registers[567][6] ) );
  EDFFX1 \registers_reg[567][5]  ( .D(n8268), .E(n757), .CK(clk), .Q(
        \registers[567][5] ) );
  EDFFX1 \registers_reg[567][4]  ( .D(n8210), .E(n757), .CK(clk), .Q(
        \registers[567][4] ) );
  EDFFX1 \registers_reg[567][3]  ( .D(n8169), .E(n757), .CK(clk), .Q(
        \registers[567][3] ) );
  EDFFX1 \registers_reg[567][2]  ( .D(n8115), .E(n757), .CK(clk), .Q(
        \registers[567][2] ) );
  EDFFX1 \registers_reg[567][1]  ( .D(n8059), .E(n757), .CK(clk), .Q(
        \registers[567][1] ) );
  EDFFX1 \registers_reg[567][0]  ( .D(n8000), .E(n757), .CK(clk), .Q(
        \registers[567][0] ) );
  EDFFX1 \registers_reg[563][7]  ( .D(n8423), .E(n70), .CK(clk), .Q(
        \registers[563][7] ) );
  EDFFX1 \registers_reg[563][6]  ( .D(n8365), .E(n70), .CK(clk), .Q(
        \registers[563][6] ) );
  EDFFX1 \registers_reg[563][5]  ( .D(n8307), .E(n70), .CK(clk), .Q(
        \registers[563][5] ) );
  EDFFX1 \registers_reg[563][4]  ( .D(n8249), .E(n70), .CK(clk), .Q(
        \registers[563][4] ) );
  EDFFX1 \registers_reg[563][3]  ( .D(n8164), .E(n70), .CK(clk), .Q(
        \registers[563][3] ) );
  EDFFX1 \registers_reg[563][2]  ( .D(n8116), .E(n70), .CK(clk), .Q(
        \registers[563][2] ) );
  EDFFX1 \registers_reg[563][1]  ( .D(n8060), .E(n70), .CK(clk), .Q(
        \registers[563][1] ) );
  EDFFX1 \registers_reg[563][0]  ( .D(n7998), .E(n70), .CK(clk), .Q(
        \registers[563][0] ) );
  EDFFX1 \registers_reg[559][7]  ( .D(n8385), .E(n66), .CK(clk), .Q(
        \registers[559][7] ) );
  EDFFX1 \registers_reg[559][6]  ( .D(n8327), .E(n66), .CK(clk), .Q(
        \registers[559][6] ) );
  EDFFX1 \registers_reg[559][5]  ( .D(n8269), .E(n66), .CK(clk), .Q(
        \registers[559][5] ) );
  EDFFX1 \registers_reg[559][4]  ( .D(n8211), .E(n66), .CK(clk), .Q(
        \registers[559][4] ) );
  EDFFX1 \registers_reg[559][3]  ( .D(n8165), .E(n66), .CK(clk), .Q(
        \registers[559][3] ) );
  EDFFX1 \registers_reg[559][2]  ( .D(n8114), .E(n66), .CK(clk), .Q(
        \registers[559][2] ) );
  EDFFX1 \registers_reg[559][1]  ( .D(n8058), .E(n66), .CK(clk), .Q(
        \registers[559][1] ) );
  EDFFX1 \registers_reg[559][0]  ( .D(n7999), .E(n66), .CK(clk), .Q(
        \registers[559][0] ) );
  EDFFX1 \registers_reg[555][7]  ( .D(n8384), .E(n62), .CK(clk), .Q(
        \registers[555][7] ) );
  EDFFX1 \registers_reg[555][6]  ( .D(n8326), .E(n62), .CK(clk), .Q(
        \registers[555][6] ) );
  EDFFX1 \registers_reg[555][5]  ( .D(n8268), .E(n62), .CK(clk), .Q(
        \registers[555][5] ) );
  EDFFX1 \registers_reg[555][4]  ( .D(n8210), .E(n62), .CK(clk), .Q(
        \registers[555][4] ) );
  EDFFX1 \registers_reg[555][3]  ( .D(n8166), .E(n62), .CK(clk), .Q(
        \registers[555][3] ) );
  EDFFX1 \registers_reg[555][2]  ( .D(n8115), .E(n62), .CK(clk), .Q(
        \registers[555][2] ) );
  EDFFX1 \registers_reg[555][1]  ( .D(n8059), .E(n62), .CK(clk), .Q(
        \registers[555][1] ) );
  EDFFX1 \registers_reg[555][0]  ( .D(n8000), .E(n62), .CK(clk), .Q(
        \registers[555][0] ) );
  EDFFX1 \registers_reg[551][7]  ( .D(n8419), .E(n273), .CK(clk), .Q(
        \registers[551][7] ) );
  EDFFX1 \registers_reg[551][6]  ( .D(n8361), .E(n273), .CK(clk), .Q(
        \registers[551][6] ) );
  EDFFX1 \registers_reg[551][5]  ( .D(n8303), .E(n273), .CK(clk), .Q(
        \registers[551][5] ) );
  EDFFX1 \registers_reg[551][4]  ( .D(n8245), .E(n273), .CK(clk), .Q(
        \registers[551][4] ) );
  EDFFX1 \registers_reg[551][3]  ( .D(n8164), .E(n273), .CK(clk), .Q(
        \registers[551][3] ) );
  EDFFX1 \registers_reg[551][2]  ( .D(n8116), .E(n273), .CK(clk), .Q(
        \registers[551][2] ) );
  EDFFX1 \registers_reg[551][1]  ( .D(n8060), .E(n273), .CK(clk), .Q(
        \registers[551][1] ) );
  EDFFX1 \registers_reg[551][0]  ( .D(n7998), .E(n273), .CK(clk), .Q(
        \registers[551][0] ) );
  EDFFX1 \registers_reg[547][7]  ( .D(n8385), .E(n269), .CK(clk), .Q(
        \registers[547][7] ) );
  EDFFX1 \registers_reg[547][6]  ( .D(n8327), .E(n269), .CK(clk), .Q(
        \registers[547][6] ) );
  EDFFX1 \registers_reg[547][5]  ( .D(n8269), .E(n269), .CK(clk), .Q(
        \registers[547][5] ) );
  EDFFX1 \registers_reg[547][4]  ( .D(n8211), .E(n269), .CK(clk), .Q(
        \registers[547][4] ) );
  EDFFX1 \registers_reg[547][3]  ( .D(n8165), .E(n269), .CK(clk), .Q(
        \registers[547][3] ) );
  EDFFX1 \registers_reg[547][2]  ( .D(n8114), .E(n269), .CK(clk), .Q(
        \registers[547][2] ) );
  EDFFX1 \registers_reg[547][1]  ( .D(n8058), .E(n269), .CK(clk), .Q(
        \registers[547][1] ) );
  EDFFX1 \registers_reg[547][0]  ( .D(n7999), .E(n269), .CK(clk), .Q(
        \registers[547][0] ) );
  EDFFX1 \registers_reg[543][7]  ( .D(n8384), .E(n753), .CK(clk), .Q(
        \registers[543][7] ) );
  EDFFX1 \registers_reg[543][6]  ( .D(n8326), .E(n753), .CK(clk), .Q(
        \registers[543][6] ) );
  EDFFX1 \registers_reg[543][5]  ( .D(n8268), .E(n753), .CK(clk), .Q(
        \registers[543][5] ) );
  EDFFX1 \registers_reg[543][4]  ( .D(n8210), .E(n753), .CK(clk), .Q(
        \registers[543][4] ) );
  EDFFX1 \registers_reg[543][3]  ( .D(n8166), .E(n753), .CK(clk), .Q(
        \registers[543][3] ) );
  EDFFX1 \registers_reg[543][2]  ( .D(n8115), .E(n753), .CK(clk), .Q(
        \registers[543][2] ) );
  EDFFX1 \registers_reg[543][1]  ( .D(n8059), .E(n753), .CK(clk), .Q(
        \registers[543][1] ) );
  EDFFX1 \registers_reg[543][0]  ( .D(n8000), .E(n753), .CK(clk), .Q(
        \registers[543][0] ) );
  EDFFX1 \registers_reg[539][7]  ( .D(n8420), .E(n749), .CK(clk), .Q(
        \registers[539][7] ) );
  EDFFX1 \registers_reg[539][6]  ( .D(n8362), .E(n749), .CK(clk), .Q(
        \registers[539][6] ) );
  EDFFX1 \registers_reg[539][5]  ( .D(n8304), .E(n749), .CK(clk), .Q(
        \registers[539][5] ) );
  EDFFX1 \registers_reg[539][4]  ( .D(n8246), .E(n749), .CK(clk), .Q(
        \registers[539][4] ) );
  EDFFX1 \registers_reg[539][3]  ( .D(n8164), .E(n749), .CK(clk), .Q(
        \registers[539][3] ) );
  EDFFX1 \registers_reg[539][2]  ( .D(n8116), .E(n749), .CK(clk), .Q(
        \registers[539][2] ) );
  EDFFX1 \registers_reg[539][1]  ( .D(n8060), .E(n749), .CK(clk), .Q(
        \registers[539][1] ) );
  EDFFX1 \registers_reg[539][0]  ( .D(n7998), .E(n749), .CK(clk), .Q(
        \registers[539][0] ) );
  EDFFX1 \registers_reg[535][7]  ( .D(n8385), .E(n745), .CK(clk), .Q(
        \registers[535][7] ) );
  EDFFX1 \registers_reg[535][6]  ( .D(n8327), .E(n745), .CK(clk), .Q(
        \registers[535][6] ) );
  EDFFX1 \registers_reg[535][5]  ( .D(n8269), .E(n745), .CK(clk), .Q(
        \registers[535][5] ) );
  EDFFX1 \registers_reg[535][4]  ( .D(n8211), .E(n745), .CK(clk), .Q(
        \registers[535][4] ) );
  EDFFX1 \registers_reg[535][3]  ( .D(n8165), .E(n745), .CK(clk), .Q(
        \registers[535][3] ) );
  EDFFX1 \registers_reg[535][2]  ( .D(n8114), .E(n745), .CK(clk), .Q(
        \registers[535][2] ) );
  EDFFX1 \registers_reg[535][1]  ( .D(n8058), .E(n745), .CK(clk), .Q(
        \registers[535][1] ) );
  EDFFX1 \registers_reg[535][0]  ( .D(n7999), .E(n745), .CK(clk), .Q(
        \registers[535][0] ) );
  EDFFX1 \registers_reg[531][7]  ( .D(n8384), .E(n58), .CK(clk), .Q(
        \registers[531][7] ) );
  EDFFX1 \registers_reg[531][6]  ( .D(n8326), .E(n58), .CK(clk), .Q(
        \registers[531][6] ) );
  EDFFX1 \registers_reg[531][5]  ( .D(n8268), .E(n58), .CK(clk), .Q(
        \registers[531][5] ) );
  EDFFX1 \registers_reg[531][4]  ( .D(n8210), .E(n58), .CK(clk), .Q(
        \registers[531][4] ) );
  EDFFX1 \registers_reg[531][3]  ( .D(n8166), .E(n58), .CK(clk), .Q(
        \registers[531][3] ) );
  EDFFX1 \registers_reg[531][2]  ( .D(n8115), .E(n58), .CK(clk), .Q(
        \registers[531][2] ) );
  EDFFX1 \registers_reg[531][1]  ( .D(n8059), .E(n58), .CK(clk), .Q(
        \registers[531][1] ) );
  EDFFX1 \registers_reg[531][0]  ( .D(n8000), .E(n58), .CK(clk), .Q(
        \registers[531][0] ) );
  EDFFX1 \registers_reg[527][7]  ( .D(n8432), .E(n53), .CK(clk), .Q(
        \registers[527][7] ) );
  EDFFX1 \registers_reg[527][6]  ( .D(n8374), .E(n53), .CK(clk), .Q(
        \registers[527][6] ) );
  EDFFX1 \registers_reg[527][5]  ( .D(n8316), .E(n53), .CK(clk), .Q(
        \registers[527][5] ) );
  EDFFX1 \registers_reg[527][4]  ( .D(n8258), .E(n53), .CK(clk), .Q(
        \registers[527][4] ) );
  EDFFX1 \registers_reg[527][3]  ( .D(n8164), .E(n53), .CK(clk), .Q(
        \registers[527][3] ) );
  EDFFX1 \registers_reg[527][2]  ( .D(n8113), .E(n53), .CK(clk), .Q(
        \registers[527][2] ) );
  EDFFX1 \registers_reg[527][1]  ( .D(n8057), .E(n53), .CK(clk), .Q(
        \registers[527][1] ) );
  EDFFX1 \registers_reg[527][0]  ( .D(n7996), .E(n53), .CK(clk), .Q(
        \registers[527][0] ) );
  EDFFX1 \registers_reg[523][7]  ( .D(n8381), .E(n49), .CK(clk), .Q(
        \registers[523][7] ) );
  EDFFX1 \registers_reg[523][6]  ( .D(n8323), .E(n49), .CK(clk), .Q(
        \registers[523][6] ) );
  EDFFX1 \registers_reg[523][5]  ( .D(n8265), .E(n49), .CK(clk), .Q(
        \registers[523][5] ) );
  EDFFX1 \registers_reg[523][4]  ( .D(n8207), .E(n49), .CK(clk), .Q(
        \registers[523][4] ) );
  EDFFX1 \registers_reg[523][3]  ( .D(n8165), .E(n49), .CK(clk), .Q(
        \registers[523][3] ) );
  EDFFX1 \registers_reg[523][2]  ( .D(n8111), .E(n49), .CK(clk), .Q(
        \registers[523][2] ) );
  EDFFX1 \registers_reg[523][1]  ( .D(n8055), .E(n49), .CK(clk), .Q(
        \registers[523][1] ) );
  EDFFX1 \registers_reg[523][0]  ( .D(n7997), .E(n49), .CK(clk), .Q(
        \registers[523][0] ) );
  EDFFX1 \registers_reg[519][7]  ( .D(n8382), .E(n266), .CK(clk), .Q(
        \registers[519][7] ) );
  EDFFX1 \registers_reg[519][6]  ( .D(n8324), .E(n266), .CK(clk), .Q(
        \registers[519][6] ) );
  EDFFX1 \registers_reg[519][5]  ( .D(n8266), .E(n266), .CK(clk), .Q(
        \registers[519][5] ) );
  EDFFX1 \registers_reg[519][4]  ( .D(n8208), .E(n266), .CK(clk), .Q(
        \registers[519][4] ) );
  EDFFX1 \registers_reg[519][3]  ( .D(n8166), .E(n266), .CK(clk), .Q(
        \registers[519][3] ) );
  EDFFX1 \registers_reg[519][2]  ( .D(n8112), .E(n266), .CK(clk), .Q(
        \registers[519][2] ) );
  EDFFX1 \registers_reg[519][1]  ( .D(n8056), .E(n266), .CK(clk), .Q(
        \registers[519][1] ) );
  EDFFX1 \registers_reg[519][0]  ( .D(n8678), .E(n266), .CK(clk), .Q(
        \registers[519][0] ) );
  EDFFX1 \registers_reg[515][7]  ( .D(n8383), .E(n262), .CK(clk), .Q(
        \registers[515][7] ) );
  EDFFX1 \registers_reg[515][6]  ( .D(n8325), .E(n262), .CK(clk), .Q(
        \registers[515][6] ) );
  EDFFX1 \registers_reg[515][5]  ( .D(n8267), .E(n262), .CK(clk), .Q(
        \registers[515][5] ) );
  EDFFX1 \registers_reg[515][4]  ( .D(n8209), .E(n262), .CK(clk), .Q(
        \registers[515][4] ) );
  EDFFX1 \registers_reg[515][3]  ( .D(n8164), .E(n262), .CK(clk), .Q(
        \registers[515][3] ) );
  EDFFX1 \registers_reg[515][2]  ( .D(n8113), .E(n262), .CK(clk), .Q(
        \registers[515][2] ) );
  EDFFX1 \registers_reg[515][1]  ( .D(n8057), .E(n262), .CK(clk), .Q(
        \registers[515][1] ) );
  EDFFX1 \registers_reg[515][0]  ( .D(n7996), .E(n262), .CK(clk), .Q(
        \registers[515][0] ) );
  EDFFX1 \registers_reg[511][7]  ( .D(n8428), .E(n741), .CK(clk), .Q(
        \registers[511][7] ) );
  EDFFX1 \registers_reg[511][6]  ( .D(n8370), .E(n741), .CK(clk), .Q(
        \registers[511][6] ) );
  EDFFX1 \registers_reg[511][5]  ( .D(n8312), .E(n741), .CK(clk), .Q(
        \registers[511][5] ) );
  EDFFX1 \registers_reg[511][4]  ( .D(n8254), .E(n741), .CK(clk), .Q(
        \registers[511][4] ) );
  EDFFX1 \registers_reg[511][3]  ( .D(n8202), .E(n741), .CK(clk), .Q(
        \registers[511][3] ) );
  EDFFX1 \registers_reg[511][2]  ( .D(n8156), .E(n741), .CK(clk), .Q(
        \registers[511][2] ) );
  EDFFX1 \registers_reg[511][1]  ( .D(n8100), .E(n741), .CK(clk), .Q(
        \registers[511][1] ) );
  EDFFX1 \registers_reg[511][0]  ( .D(n8005), .E(n741), .CK(clk), .Q(
        \registers[511][0] ) );
  EDFFX1 \registers_reg[507][7]  ( .D(n8429), .E(n737), .CK(clk), .Q(
        \registers[507][7] ) );
  EDFFX1 \registers_reg[507][6]  ( .D(n8371), .E(n737), .CK(clk), .Q(
        \registers[507][6] ) );
  EDFFX1 \registers_reg[507][5]  ( .D(n8313), .E(n737), .CK(clk), .Q(
        \registers[507][5] ) );
  EDFFX1 \registers_reg[507][4]  ( .D(n8255), .E(n737), .CK(clk), .Q(
        \registers[507][4] ) );
  EDFFX1 \registers_reg[507][3]  ( .D(n8200), .E(n737), .CK(clk), .Q(
        \registers[507][3] ) );
  EDFFX1 \registers_reg[507][2]  ( .D(n8157), .E(n737), .CK(clk), .Q(
        \registers[507][2] ) );
  EDFFX1 \registers_reg[507][1]  ( .D(n8101), .E(n737), .CK(clk), .Q(
        \registers[507][1] ) );
  EDFFX1 \registers_reg[507][0]  ( .D(n8041), .E(n737), .CK(clk), .Q(
        \registers[507][0] ) );
  EDFFX1 \registers_reg[503][7]  ( .D(n8425), .E(n733), .CK(clk), .Q(
        \registers[503][7] ) );
  EDFFX1 \registers_reg[503][6]  ( .D(n8367), .E(n733), .CK(clk), .Q(
        \registers[503][6] ) );
  EDFFX1 \registers_reg[503][5]  ( .D(n8309), .E(n733), .CK(clk), .Q(
        \registers[503][5] ) );
  EDFFX1 \registers_reg[503][4]  ( .D(n8251), .E(n733), .CK(clk), .Q(
        \registers[503][4] ) );
  EDFFX1 \registers_reg[503][3]  ( .D(n8201), .E(n733), .CK(clk), .Q(
        \registers[503][3] ) );
  EDFFX1 \registers_reg[503][2]  ( .D(n8155), .E(n733), .CK(clk), .Q(
        \registers[503][2] ) );
  EDFFX1 \registers_reg[503][1]  ( .D(n8099), .E(n733), .CK(clk), .Q(
        \registers[503][1] ) );
  EDFFX1 \registers_reg[503][0]  ( .D(n8042), .E(n733), .CK(clk), .Q(
        \registers[503][0] ) );
  EDFFX1 \registers_reg[499][7]  ( .D(n8426), .E(n45), .CK(clk), .Q(
        \registers[499][7] ) );
  EDFFX1 \registers_reg[499][6]  ( .D(n8368), .E(n45), .CK(clk), .Q(
        \registers[499][6] ) );
  EDFFX1 \registers_reg[499][5]  ( .D(n8310), .E(n45), .CK(clk), .Q(
        \registers[499][5] ) );
  EDFFX1 \registers_reg[499][4]  ( .D(n8252), .E(n45), .CK(clk), .Q(
        \registers[499][4] ) );
  EDFFX1 \registers_reg[499][3]  ( .D(n8202), .E(n45), .CK(clk), .Q(
        \registers[499][3] ) );
  EDFFX1 \registers_reg[499][2]  ( .D(n8156), .E(n45), .CK(clk), .Q(
        \registers[499][2] ) );
  EDFFX1 \registers_reg[499][1]  ( .D(n8100), .E(n45), .CK(clk), .Q(
        \registers[499][1] ) );
  EDFFX1 \registers_reg[499][0]  ( .D(n8040), .E(n45), .CK(clk), .Q(
        \registers[499][0] ) );
  EDFFX1 \registers_reg[495][7]  ( .D(n8427), .E(n41), .CK(clk), .Q(
        \registers[495][7] ) );
  EDFFX1 \registers_reg[495][6]  ( .D(n8369), .E(n41), .CK(clk), .Q(
        \registers[495][6] ) );
  EDFFX1 \registers_reg[495][5]  ( .D(n8311), .E(n41), .CK(clk), .Q(
        \registers[495][5] ) );
  EDFFX1 \registers_reg[495][4]  ( .D(n8253), .E(n41), .CK(clk), .Q(
        \registers[495][4] ) );
  EDFFX1 \registers_reg[495][3]  ( .D(n8200), .E(n41), .CK(clk), .Q(
        \registers[495][3] ) );
  EDFFX1 \registers_reg[495][2]  ( .D(n8157), .E(n41), .CK(clk), .Q(
        \registers[495][2] ) );
  EDFFX1 \registers_reg[495][1]  ( .D(n8101), .E(n41), .CK(clk), .Q(
        \registers[495][1] ) );
  EDFFX1 \registers_reg[495][0]  ( .D(n8041), .E(n41), .CK(clk), .Q(
        \registers[495][0] ) );
  EDFFX1 \registers_reg[491][7]  ( .D(n8425), .E(n37), .CK(clk), .Q(
        \registers[491][7] ) );
  EDFFX1 \registers_reg[491][6]  ( .D(n8367), .E(n37), .CK(clk), .Q(
        \registers[491][6] ) );
  EDFFX1 \registers_reg[491][5]  ( .D(n8309), .E(n37), .CK(clk), .Q(
        \registers[491][5] ) );
  EDFFX1 \registers_reg[491][4]  ( .D(n8251), .E(n37), .CK(clk), .Q(
        \registers[491][4] ) );
  EDFFX1 \registers_reg[491][3]  ( .D(n8201), .E(n37), .CK(clk), .Q(
        \registers[491][3] ) );
  EDFFX1 \registers_reg[491][2]  ( .D(n8155), .E(n37), .CK(clk), .Q(
        \registers[491][2] ) );
  EDFFX1 \registers_reg[491][1]  ( .D(n8099), .E(n37), .CK(clk), .Q(
        \registers[491][1] ) );
  EDFFX1 \registers_reg[491][0]  ( .D(n8042), .E(n37), .CK(clk), .Q(
        \registers[491][0] ) );
  EDFFX1 \registers_reg[487][7]  ( .D(n8426), .E(n259), .CK(clk), .Q(
        \registers[487][7] ) );
  EDFFX1 \registers_reg[487][6]  ( .D(n8368), .E(n259), .CK(clk), .Q(
        \registers[487][6] ) );
  EDFFX1 \registers_reg[487][5]  ( .D(n8310), .E(n259), .CK(clk), .Q(
        \registers[487][5] ) );
  EDFFX1 \registers_reg[487][4]  ( .D(n8252), .E(n259), .CK(clk), .Q(
        \registers[487][4] ) );
  EDFFX1 \registers_reg[487][3]  ( .D(n8202), .E(n259), .CK(clk), .Q(
        \registers[487][3] ) );
  EDFFX1 \registers_reg[487][2]  ( .D(n8156), .E(n259), .CK(clk), .Q(
        \registers[487][2] ) );
  EDFFX1 \registers_reg[487][1]  ( .D(n8100), .E(n259), .CK(clk), .Q(
        \registers[487][1] ) );
  EDFFX1 \registers_reg[487][0]  ( .D(n8040), .E(n259), .CK(clk), .Q(
        \registers[487][0] ) );
  EDFFX1 \registers_reg[483][7]  ( .D(n8427), .E(n255), .CK(clk), .Q(
        \registers[483][7] ) );
  EDFFX1 \registers_reg[483][6]  ( .D(n8369), .E(n255), .CK(clk), .Q(
        \registers[483][6] ) );
  EDFFX1 \registers_reg[483][5]  ( .D(n8311), .E(n255), .CK(clk), .Q(
        \registers[483][5] ) );
  EDFFX1 \registers_reg[483][4]  ( .D(n8253), .E(n255), .CK(clk), .Q(
        \registers[483][4] ) );
  EDFFX1 \registers_reg[483][3]  ( .D(n8197), .E(n255), .CK(clk), .Q(
        \registers[483][3] ) );
  EDFFX1 \registers_reg[483][2]  ( .D(n8157), .E(n255), .CK(clk), .Q(
        \registers[483][2] ) );
  EDFFX1 \registers_reg[483][1]  ( .D(n8101), .E(n255), .CK(clk), .Q(
        \registers[483][1] ) );
  EDFFX1 \registers_reg[483][0]  ( .D(n8041), .E(n255), .CK(clk), .Q(
        \registers[483][0] ) );
  EDFFX1 \registers_reg[479][7]  ( .D(n8425), .E(n729), .CK(clk), .Q(
        \registers[479][7] ) );
  EDFFX1 \registers_reg[479][6]  ( .D(n8367), .E(n729), .CK(clk), .Q(
        \registers[479][6] ) );
  EDFFX1 \registers_reg[479][5]  ( .D(n8309), .E(n729), .CK(clk), .Q(
        \registers[479][5] ) );
  EDFFX1 \registers_reg[479][4]  ( .D(n8251), .E(n729), .CK(clk), .Q(
        \registers[479][4] ) );
  EDFFX1 \registers_reg[479][3]  ( .D(n8198), .E(n729), .CK(clk), .Q(
        \registers[479][3] ) );
  EDFFX1 \registers_reg[479][2]  ( .D(n8155), .E(n729), .CK(clk), .Q(
        \registers[479][2] ) );
  EDFFX1 \registers_reg[479][1]  ( .D(n8099), .E(n729), .CK(clk), .Q(
        \registers[479][1] ) );
  EDFFX1 \registers_reg[479][0]  ( .D(n8042), .E(n729), .CK(clk), .Q(
        \registers[479][0] ) );
  EDFFX1 \registers_reg[475][7]  ( .D(n8426), .E(n725), .CK(clk), .Q(
        \registers[475][7] ) );
  EDFFX1 \registers_reg[475][6]  ( .D(n8368), .E(n725), .CK(clk), .Q(
        \registers[475][6] ) );
  EDFFX1 \registers_reg[475][5]  ( .D(n8310), .E(n725), .CK(clk), .Q(
        \registers[475][5] ) );
  EDFFX1 \registers_reg[475][4]  ( .D(n8252), .E(n725), .CK(clk), .Q(
        \registers[475][4] ) );
  EDFFX1 \registers_reg[475][3]  ( .D(n8199), .E(n725), .CK(clk), .Q(
        \registers[475][3] ) );
  EDFFX1 \registers_reg[475][2]  ( .D(n8156), .E(n725), .CK(clk), .Q(
        \registers[475][2] ) );
  EDFFX1 \registers_reg[475][1]  ( .D(n8100), .E(n725), .CK(clk), .Q(
        \registers[475][1] ) );
  EDFFX1 \registers_reg[475][0]  ( .D(n8040), .E(n725), .CK(clk), .Q(
        \registers[475][0] ) );
  EDFFX1 \registers_reg[471][7]  ( .D(n8427), .E(n721), .CK(clk), .Q(
        \registers[471][7] ) );
  EDFFX1 \registers_reg[471][6]  ( .D(n8369), .E(n721), .CK(clk), .Q(
        \registers[471][6] ) );
  EDFFX1 \registers_reg[471][5]  ( .D(n8311), .E(n721), .CK(clk), .Q(
        \registers[471][5] ) );
  EDFFX1 \registers_reg[471][4]  ( .D(n8253), .E(n721), .CK(clk), .Q(
        \registers[471][4] ) );
  EDFFX1 \registers_reg[471][3]  ( .D(n8197), .E(n721), .CK(clk), .Q(
        \registers[471][3] ) );
  EDFFX1 \registers_reg[471][2]  ( .D(n8154), .E(n721), .CK(clk), .Q(
        \registers[471][2] ) );
  EDFFX1 \registers_reg[471][1]  ( .D(n8098), .E(n721), .CK(clk), .Q(
        \registers[471][1] ) );
  EDFFX1 \registers_reg[471][0]  ( .D(n8038), .E(n721), .CK(clk), .Q(
        \registers[471][0] ) );
  EDFFX1 \registers_reg[467][7]  ( .D(n8425), .E(n33), .CK(clk), .Q(
        \registers[467][7] ) );
  EDFFX1 \registers_reg[467][6]  ( .D(n8367), .E(n33), .CK(clk), .Q(
        \registers[467][6] ) );
  EDFFX1 \registers_reg[467][5]  ( .D(n8309), .E(n33), .CK(clk), .Q(
        \registers[467][5] ) );
  EDFFX1 \registers_reg[467][4]  ( .D(n8251), .E(n33), .CK(clk), .Q(
        \registers[467][4] ) );
  EDFFX1 \registers_reg[467][3]  ( .D(n8198), .E(n33), .CK(clk), .Q(
        \registers[467][3] ) );
  EDFFX1 \registers_reg[467][2]  ( .D(n8152), .E(n33), .CK(clk), .Q(
        \registers[467][2] ) );
  EDFFX1 \registers_reg[467][1]  ( .D(n8096), .E(n33), .CK(clk), .Q(
        \registers[467][1] ) );
  EDFFX1 \registers_reg[467][0]  ( .D(n8039), .E(n33), .CK(clk), .Q(
        \registers[467][0] ) );
  EDFFX1 \registers_reg[463][7]  ( .D(n8426), .E(n29), .CK(clk), .Q(
        \registers[463][7] ) );
  EDFFX1 \registers_reg[463][6]  ( .D(n8368), .E(n29), .CK(clk), .Q(
        \registers[463][6] ) );
  EDFFX1 \registers_reg[463][5]  ( .D(n8310), .E(n29), .CK(clk), .Q(
        \registers[463][5] ) );
  EDFFX1 \registers_reg[463][4]  ( .D(n8252), .E(n29), .CK(clk), .Q(
        \registers[463][4] ) );
  EDFFX1 \registers_reg[463][3]  ( .D(n8199), .E(n29), .CK(clk), .Q(
        \registers[463][3] ) );
  EDFFX1 \registers_reg[463][2]  ( .D(n8153), .E(n29), .CK(clk), .Q(
        \registers[463][2] ) );
  EDFFX1 \registers_reg[463][1]  ( .D(n8097), .E(n29), .CK(clk), .Q(
        \registers[463][1] ) );
  EDFFX1 \registers_reg[463][0]  ( .D(n8037), .E(n29), .CK(clk), .Q(
        \registers[463][0] ) );
  EDFFX1 \registers_reg[459][7]  ( .D(n8427), .E(n25), .CK(clk), .Q(
        \registers[459][7] ) );
  EDFFX1 \registers_reg[459][6]  ( .D(n8369), .E(n25), .CK(clk), .Q(
        \registers[459][6] ) );
  EDFFX1 \registers_reg[459][5]  ( .D(n8311), .E(n25), .CK(clk), .Q(
        \registers[459][5] ) );
  EDFFX1 \registers_reg[459][4]  ( .D(n8253), .E(n25), .CK(clk), .Q(
        \registers[459][4] ) );
  EDFFX1 \registers_reg[459][3]  ( .D(n8197), .E(n25), .CK(clk), .Q(
        \registers[459][3] ) );
  EDFFX1 \registers_reg[459][2]  ( .D(n8154), .E(n25), .CK(clk), .Q(
        \registers[459][2] ) );
  EDFFX1 \registers_reg[459][1]  ( .D(n8098), .E(n25), .CK(clk), .Q(
        \registers[459][1] ) );
  EDFFX1 \registers_reg[459][0]  ( .D(n8038), .E(n25), .CK(clk), .Q(
        \registers[459][0] ) );
  EDFFX1 \registers_reg[455][7]  ( .D(n8423), .E(n252), .CK(clk), .Q(
        \registers[455][7] ) );
  EDFFX1 \registers_reg[455][6]  ( .D(n8365), .E(n252), .CK(clk), .Q(
        \registers[455][6] ) );
  EDFFX1 \registers_reg[455][5]  ( .D(n8307), .E(n252), .CK(clk), .Q(
        \registers[455][5] ) );
  EDFFX1 \registers_reg[455][4]  ( .D(n8249), .E(n252), .CK(clk), .Q(
        \registers[455][4] ) );
  EDFFX1 \registers_reg[455][3]  ( .D(n8198), .E(n252), .CK(clk), .Q(
        \registers[455][3] ) );
  EDFFX1 \registers_reg[455][2]  ( .D(n8152), .E(n252), .CK(clk), .Q(
        \registers[455][2] ) );
  EDFFX1 \registers_reg[455][1]  ( .D(n8096), .E(n252), .CK(clk), .Q(
        \registers[455][1] ) );
  EDFFX1 \registers_reg[455][0]  ( .D(n8039), .E(n252), .CK(clk), .Q(
        \registers[455][0] ) );
  EDFFX1 \registers_reg[451][7]  ( .D(n8424), .E(n248), .CK(clk), .Q(
        \registers[451][7] ) );
  EDFFX1 \registers_reg[451][6]  ( .D(n8366), .E(n248), .CK(clk), .Q(
        \registers[451][6] ) );
  EDFFX1 \registers_reg[451][5]  ( .D(n8308), .E(n248), .CK(clk), .Q(
        \registers[451][5] ) );
  EDFFX1 \registers_reg[451][4]  ( .D(n8250), .E(n248), .CK(clk), .Q(
        \registers[451][4] ) );
  EDFFX1 \registers_reg[451][3]  ( .D(n8199), .E(n248), .CK(clk), .Q(
        \registers[451][3] ) );
  EDFFX1 \registers_reg[451][2]  ( .D(n8153), .E(n248), .CK(clk), .Q(
        \registers[451][2] ) );
  EDFFX1 \registers_reg[451][1]  ( .D(n8097), .E(n248), .CK(clk), .Q(
        \registers[451][1] ) );
  EDFFX1 \registers_reg[451][0]  ( .D(n8037), .E(n248), .CK(clk), .Q(
        \registers[451][0] ) );
  EDFFX1 \registers_reg[447][7]  ( .D(n8423), .E(n717), .CK(clk), .Q(
        \registers[447][7] ) );
  EDFFX1 \registers_reg[447][6]  ( .D(n8365), .E(n717), .CK(clk), .Q(
        \registers[447][6] ) );
  EDFFX1 \registers_reg[447][5]  ( .D(n8307), .E(n717), .CK(clk), .Q(
        \registers[447][5] ) );
  EDFFX1 \registers_reg[447][4]  ( .D(n8249), .E(n717), .CK(clk), .Q(
        \registers[447][4] ) );
  EDFFX1 \registers_reg[447][3]  ( .D(n8198), .E(n717), .CK(clk), .Q(
        \registers[447][3] ) );
  EDFFX1 \registers_reg[447][2]  ( .D(n8152), .E(n717), .CK(clk), .Q(
        \registers[447][2] ) );
  EDFFX1 \registers_reg[447][1]  ( .D(n8096), .E(n717), .CK(clk), .Q(
        \registers[447][1] ) );
  EDFFX1 \registers_reg[447][0]  ( .D(n8038), .E(n717), .CK(clk), .Q(
        \registers[447][0] ) );
  EDFFX1 \registers_reg[443][7]  ( .D(n8424), .E(n713), .CK(clk), .Q(
        \registers[443][7] ) );
  EDFFX1 \registers_reg[443][6]  ( .D(n8366), .E(n713), .CK(clk), .Q(
        \registers[443][6] ) );
  EDFFX1 \registers_reg[443][5]  ( .D(n8308), .E(n713), .CK(clk), .Q(
        \registers[443][5] ) );
  EDFFX1 \registers_reg[443][4]  ( .D(n8250), .E(n713), .CK(clk), .Q(
        \registers[443][4] ) );
  EDFFX1 \registers_reg[443][3]  ( .D(n8199), .E(n713), .CK(clk), .Q(
        \registers[443][3] ) );
  EDFFX1 \registers_reg[443][2]  ( .D(n8153), .E(n713), .CK(clk), .Q(
        \registers[443][2] ) );
  EDFFX1 \registers_reg[443][1]  ( .D(n8097), .E(n713), .CK(clk), .Q(
        \registers[443][1] ) );
  EDFFX1 \registers_reg[443][0]  ( .D(n8037), .E(n713), .CK(clk), .Q(
        \registers[443][0] ) );
  EDFFX1 \registers_reg[439][7]  ( .D(n8422), .E(n709), .CK(clk), .Q(
        \registers[439][7] ) );
  EDFFX1 \registers_reg[439][6]  ( .D(n8364), .E(n709), .CK(clk), .Q(
        \registers[439][6] ) );
  EDFFX1 \registers_reg[439][5]  ( .D(n8306), .E(n709), .CK(clk), .Q(
        \registers[439][5] ) );
  EDFFX1 \registers_reg[439][4]  ( .D(n8248), .E(n709), .CK(clk), .Q(
        \registers[439][4] ) );
  EDFFX1 \registers_reg[439][3]  ( .D(n8197), .E(n709), .CK(clk), .Q(
        \registers[439][3] ) );
  EDFFX1 \registers_reg[439][2]  ( .D(n8154), .E(n709), .CK(clk), .Q(
        \registers[439][2] ) );
  EDFFX1 \registers_reg[439][1]  ( .D(n8098), .E(n709), .CK(clk), .Q(
        \registers[439][1] ) );
  EDFFX1 \registers_reg[439][0]  ( .D(n8038), .E(n709), .CK(clk), .Q(
        \registers[439][0] ) );
  EDFFX1 \registers_reg[435][7]  ( .D(n8423), .E(n21), .CK(clk), .Q(
        \registers[435][7] ) );
  EDFFX1 \registers_reg[435][6]  ( .D(n8365), .E(n21), .CK(clk), .Q(
        \registers[435][6] ) );
  EDFFX1 \registers_reg[435][5]  ( .D(n8307), .E(n21), .CK(clk), .Q(
        \registers[435][5] ) );
  EDFFX1 \registers_reg[435][4]  ( .D(n8249), .E(n21), .CK(clk), .Q(
        \registers[435][4] ) );
  EDFFX1 \registers_reg[435][3]  ( .D(n8198), .E(n21), .CK(clk), .Q(
        \registers[435][3] ) );
  EDFFX1 \registers_reg[435][2]  ( .D(n8152), .E(n21), .CK(clk), .Q(
        \registers[435][2] ) );
  EDFFX1 \registers_reg[435][1]  ( .D(n8096), .E(n21), .CK(clk), .Q(
        \registers[435][1] ) );
  EDFFX1 \registers_reg[435][0]  ( .D(n8039), .E(n21), .CK(clk), .Q(
        \registers[435][0] ) );
  EDFFX1 \registers_reg[431][7]  ( .D(n8424), .E(n17), .CK(clk), .Q(
        \registers[431][7] ) );
  EDFFX1 \registers_reg[431][6]  ( .D(n8366), .E(n17), .CK(clk), .Q(
        \registers[431][6] ) );
  EDFFX1 \registers_reg[431][5]  ( .D(n8308), .E(n17), .CK(clk), .Q(
        \registers[431][5] ) );
  EDFFX1 \registers_reg[431][4]  ( .D(n8250), .E(n17), .CK(clk), .Q(
        \registers[431][4] ) );
  EDFFX1 \registers_reg[431][3]  ( .D(n8199), .E(n17), .CK(clk), .Q(
        \registers[431][3] ) );
  EDFFX1 \registers_reg[431][2]  ( .D(n8153), .E(n17), .CK(clk), .Q(
        \registers[431][2] ) );
  EDFFX1 \registers_reg[431][1]  ( .D(n8097), .E(n17), .CK(clk), .Q(
        \registers[431][1] ) );
  EDFFX1 \registers_reg[431][0]  ( .D(n8037), .E(n17), .CK(clk), .Q(
        \registers[431][0] ) );
  EDFFX1 \registers_reg[427][7]  ( .D(n8422), .E(n13), .CK(clk), .Q(
        \registers[427][7] ) );
  EDFFX1 \registers_reg[427][6]  ( .D(n8364), .E(n13), .CK(clk), .Q(
        \registers[427][6] ) );
  EDFFX1 \registers_reg[427][5]  ( .D(n8306), .E(n13), .CK(clk), .Q(
        \registers[427][5] ) );
  EDFFX1 \registers_reg[427][4]  ( .D(n8248), .E(n13), .CK(clk), .Q(
        \registers[427][4] ) );
  EDFFX1 \registers_reg[427][3]  ( .D(n8197), .E(n13), .CK(clk), .Q(
        \registers[427][3] ) );
  EDFFX1 \registers_reg[427][2]  ( .D(n8154), .E(n13), .CK(clk), .Q(
        \registers[427][2] ) );
  EDFFX1 \registers_reg[427][1]  ( .D(n8098), .E(n13), .CK(clk), .Q(
        \registers[427][1] ) );
  EDFFX1 \registers_reg[427][0]  ( .D(n8038), .E(n13), .CK(clk), .Q(
        \registers[427][0] ) );
  EDFFX1 \registers_reg[423][7]  ( .D(n8423), .E(n245), .CK(clk), .Q(
        \registers[423][7] ) );
  EDFFX1 \registers_reg[423][6]  ( .D(n8365), .E(n245), .CK(clk), .Q(
        \registers[423][6] ) );
  EDFFX1 \registers_reg[423][5]  ( .D(n8307), .E(n245), .CK(clk), .Q(
        \registers[423][5] ) );
  EDFFX1 \registers_reg[423][4]  ( .D(n8249), .E(n245), .CK(clk), .Q(
        \registers[423][4] ) );
  EDFFX1 \registers_reg[423][3]  ( .D(n8195), .E(n245), .CK(clk), .Q(
        \registers[423][3] ) );
  EDFFX1 \registers_reg[423][2]  ( .D(n8150), .E(n245), .CK(clk), .Q(
        \registers[423][2] ) );
  EDFFX1 \registers_reg[423][1]  ( .D(n8094), .E(n245), .CK(clk), .Q(
        \registers[423][1] ) );
  EDFFX1 \registers_reg[423][0]  ( .D(n8039), .E(n245), .CK(clk), .Q(
        \registers[423][0] ) );
  EDFFX1 \registers_reg[419][7]  ( .D(n8424), .E(n241), .CK(clk), .Q(
        \registers[419][7] ) );
  EDFFX1 \registers_reg[419][6]  ( .D(n8366), .E(n241), .CK(clk), .Q(
        \registers[419][6] ) );
  EDFFX1 \registers_reg[419][5]  ( .D(n8308), .E(n241), .CK(clk), .Q(
        \registers[419][5] ) );
  EDFFX1 \registers_reg[419][4]  ( .D(n8250), .E(n241), .CK(clk), .Q(
        \registers[419][4] ) );
  EDFFX1 \registers_reg[419][3]  ( .D(n8196), .E(n241), .CK(clk), .Q(
        \registers[419][3] ) );
  EDFFX1 \registers_reg[419][2]  ( .D(n8151), .E(n241), .CK(clk), .Q(
        \registers[419][2] ) );
  EDFFX1 \registers_reg[419][1]  ( .D(n8095), .E(n241), .CK(clk), .Q(
        \registers[419][1] ) );
  EDFFX1 \registers_reg[419][0]  ( .D(n8034), .E(n241), .CK(clk), .Q(
        \registers[419][0] ) );
  EDFFX1 \registers_reg[415][7]  ( .D(n8422), .E(n705), .CK(clk), .Q(
        \registers[415][7] ) );
  EDFFX1 \registers_reg[415][6]  ( .D(n8364), .E(n705), .CK(clk), .Q(
        \registers[415][6] ) );
  EDFFX1 \registers_reg[415][5]  ( .D(n8306), .E(n705), .CK(clk), .Q(
        \registers[415][5] ) );
  EDFFX1 \registers_reg[415][4]  ( .D(n8248), .E(n705), .CK(clk), .Q(
        \registers[415][4] ) );
  EDFFX1 \registers_reg[415][3]  ( .D(n8194), .E(n705), .CK(clk), .Q(
        \registers[415][3] ) );
  EDFFX1 \registers_reg[415][2]  ( .D(n8733), .E(n705), .CK(clk), .Q(
        \registers[415][2] ) );
  EDFFX1 \registers_reg[415][1]  ( .D(n8705), .E(n705), .CK(clk), .Q(
        \registers[415][1] ) );
  EDFFX1 \registers_reg[415][0]  ( .D(n8035), .E(n705), .CK(clk), .Q(
        \registers[415][0] ) );
  EDFFX1 \registers_reg[411][7]  ( .D(n8423), .E(n701), .CK(clk), .Q(
        \registers[411][7] ) );
  EDFFX1 \registers_reg[411][6]  ( .D(n8365), .E(n701), .CK(clk), .Q(
        \registers[411][6] ) );
  EDFFX1 \registers_reg[411][5]  ( .D(n8307), .E(n701), .CK(clk), .Q(
        \registers[411][5] ) );
  EDFFX1 \registers_reg[411][4]  ( .D(n8249), .E(n701), .CK(clk), .Q(
        \registers[411][4] ) );
  EDFFX1 \registers_reg[411][3]  ( .D(n8195), .E(n701), .CK(clk), .Q(
        \registers[411][3] ) );
  EDFFX1 \registers_reg[411][2]  ( .D(n8150), .E(n701), .CK(clk), .Q(
        \registers[411][2] ) );
  EDFFX1 \registers_reg[411][1]  ( .D(n8094), .E(n701), .CK(clk), .Q(
        \registers[411][1] ) );
  EDFFX1 \registers_reg[411][0]  ( .D(n8036), .E(n701), .CK(clk), .Q(
        \registers[411][0] ) );
  EDFFX1 \registers_reg[407][7]  ( .D(n8419), .E(n697), .CK(clk), .Q(
        \registers[407][7] ) );
  EDFFX1 \registers_reg[407][6]  ( .D(n8361), .E(n697), .CK(clk), .Q(
        \registers[407][6] ) );
  EDFFX1 \registers_reg[407][5]  ( .D(n8303), .E(n697), .CK(clk), .Q(
        \registers[407][5] ) );
  EDFFX1 \registers_reg[407][4]  ( .D(n8245), .E(n697), .CK(clk), .Q(
        \registers[407][4] ) );
  EDFFX1 \registers_reg[407][3]  ( .D(n8196), .E(n697), .CK(clk), .Q(
        \registers[407][3] ) );
  EDFFX1 \registers_reg[407][2]  ( .D(n8151), .E(n697), .CK(clk), .Q(
        \registers[407][2] ) );
  EDFFX1 \registers_reg[407][1]  ( .D(n8095), .E(n697), .CK(clk), .Q(
        \registers[407][1] ) );
  EDFFX1 \registers_reg[407][0]  ( .D(n8034), .E(n697), .CK(clk), .Q(
        \registers[407][0] ) );
  EDFFX1 \registers_reg[403][7]  ( .D(n8420), .E(n693), .CK(clk), .Q(
        \registers[403][7] ) );
  EDFFX1 \registers_reg[403][6]  ( .D(n8362), .E(n693), .CK(clk), .Q(
        \registers[403][6] ) );
  EDFFX1 \registers_reg[403][5]  ( .D(n8304), .E(n693), .CK(clk), .Q(
        \registers[403][5] ) );
  EDFFX1 \registers_reg[403][4]  ( .D(n8246), .E(n693), .CK(clk), .Q(
        \registers[403][4] ) );
  EDFFX1 \registers_reg[403][3]  ( .D(n8194), .E(n693), .CK(clk), .Q(
        \registers[403][3] ) );
  EDFFX1 \registers_reg[403][2]  ( .D(n8732), .E(n693), .CK(clk), .Q(
        \registers[403][2] ) );
  EDFFX1 \registers_reg[403][1]  ( .D(n8704), .E(n693), .CK(clk), .Q(
        \registers[403][1] ) );
  EDFFX1 \registers_reg[403][0]  ( .D(n8035), .E(n693), .CK(clk), .Q(
        \registers[403][0] ) );
  EDFFX1 \registers_reg[399][7]  ( .D(n8421), .E(n689), .CK(clk), .Q(
        \registers[399][7] ) );
  EDFFX1 \registers_reg[399][6]  ( .D(n8363), .E(n689), .CK(clk), .Q(
        \registers[399][6] ) );
  EDFFX1 \registers_reg[399][5]  ( .D(n8305), .E(n689), .CK(clk), .Q(
        \registers[399][5] ) );
  EDFFX1 \registers_reg[399][4]  ( .D(n8247), .E(n689), .CK(clk), .Q(
        \registers[399][4] ) );
  EDFFX1 \registers_reg[399][3]  ( .D(n8195), .E(n689), .CK(clk), .Q(
        \registers[399][3] ) );
  EDFFX1 \registers_reg[399][2]  ( .D(n8150), .E(n689), .CK(clk), .Q(
        \registers[399][2] ) );
  EDFFX1 \registers_reg[399][1]  ( .D(n8094), .E(n689), .CK(clk), .Q(
        \registers[399][1] ) );
  EDFFX1 \registers_reg[399][0]  ( .D(n8036), .E(n689), .CK(clk), .Q(
        \registers[399][0] ) );
  EDFFX1 \registers_reg[395][7]  ( .D(n8419), .E(n685), .CK(clk), .Q(
        \registers[395][7] ) );
  EDFFX1 \registers_reg[395][6]  ( .D(n8361), .E(n685), .CK(clk), .Q(
        \registers[395][6] ) );
  EDFFX1 \registers_reg[395][5]  ( .D(n8303), .E(n685), .CK(clk), .Q(
        \registers[395][5] ) );
  EDFFX1 \registers_reg[395][4]  ( .D(n8245), .E(n685), .CK(clk), .Q(
        \registers[395][4] ) );
  EDFFX1 \registers_reg[395][3]  ( .D(n8196), .E(n685), .CK(clk), .Q(
        \registers[395][3] ) );
  EDFFX1 \registers_reg[395][2]  ( .D(n8151), .E(n685), .CK(clk), .Q(
        \registers[395][2] ) );
  EDFFX1 \registers_reg[395][1]  ( .D(n8095), .E(n685), .CK(clk), .Q(
        \registers[395][1] ) );
  EDFFX1 \registers_reg[395][0]  ( .D(n8034), .E(n685), .CK(clk), .Q(
        \registers[395][0] ) );
  EDFFX1 \registers_reg[391][7]  ( .D(n8420), .E(n1001), .CK(clk), .Q(
        \registers[391][7] ) );
  EDFFX1 \registers_reg[391][6]  ( .D(n8362), .E(n1001), .CK(clk), .Q(
        \registers[391][6] ) );
  EDFFX1 \registers_reg[391][5]  ( .D(n8304), .E(n1001), .CK(clk), .Q(
        \registers[391][5] ) );
  EDFFX1 \registers_reg[391][4]  ( .D(n8246), .E(n1001), .CK(clk), .Q(
        \registers[391][4] ) );
  EDFFX1 \registers_reg[391][3]  ( .D(n8194), .E(n1001), .CK(clk), .Q(
        \registers[391][3] ) );
  EDFFX1 \registers_reg[391][2]  ( .D(n8731), .E(n1001), .CK(clk), .Q(
        \registers[391][2] ) );
  EDFFX1 \registers_reg[391][1]  ( .D(n8703), .E(n1001), .CK(clk), .Q(
        \registers[391][1] ) );
  EDFFX1 \registers_reg[391][0]  ( .D(n8035), .E(n1001), .CK(clk), .Q(
        \registers[391][0] ) );
  EDFFX1 \registers_reg[387][7]  ( .D(n8421), .E(n997), .CK(clk), .Q(
        \registers[387][7] ) );
  EDFFX1 \registers_reg[387][6]  ( .D(n8363), .E(n997), .CK(clk), .Q(
        \registers[387][6] ) );
  EDFFX1 \registers_reg[387][5]  ( .D(n8305), .E(n997), .CK(clk), .Q(
        \registers[387][5] ) );
  EDFFX1 \registers_reg[387][4]  ( .D(n8247), .E(n997), .CK(clk), .Q(
        \registers[387][4] ) );
  EDFFX1 \registers_reg[387][3]  ( .D(n8195), .E(n997), .CK(clk), .Q(
        \registers[387][3] ) );
  EDFFX1 \registers_reg[387][2]  ( .D(n8150), .E(n997), .CK(clk), .Q(
        \registers[387][2] ) );
  EDFFX1 \registers_reg[387][1]  ( .D(n8094), .E(n997), .CK(clk), .Q(
        \registers[387][1] ) );
  EDFFX1 \registers_reg[387][0]  ( .D(n8036), .E(n997), .CK(clk), .Q(
        \registers[387][0] ) );
  EDFFX1 \registers_reg[383][7]  ( .D(n8433), .E(n681), .CK(clk), .Q(
        \registers[383][7] ) );
  EDFFX1 \registers_reg[383][6]  ( .D(n8375), .E(n681), .CK(clk), .Q(
        \registers[383][6] ) );
  EDFFX1 \registers_reg[383][5]  ( .D(n8317), .E(n681), .CK(clk), .Q(
        \registers[383][5] ) );
  EDFFX1 \registers_reg[383][4]  ( .D(n8259), .E(n681), .CK(clk), .Q(
        \registers[383][4] ) );
  EDFFX1 \registers_reg[383][3]  ( .D(n8193), .E(n681), .CK(clk), .Q(
        \registers[383][3] ) );
  EDFFX1 \registers_reg[383][2]  ( .D(n8115), .E(n681), .CK(clk), .Q(
        \registers[383][2] ) );
  EDFFX1 \registers_reg[383][1]  ( .D(n8059), .E(n681), .CK(clk), .Q(
        \registers[383][1] ) );
  EDFFX1 \registers_reg[383][0]  ( .D(n8039), .E(n681), .CK(clk), .Q(
        \registers[383][0] ) );
  EDFFX1 \registers_reg[379][7]  ( .D(n8434), .E(n677), .CK(clk), .Q(
        \registers[379][7] ) );
  EDFFX1 \registers_reg[379][6]  ( .D(n8376), .E(n677), .CK(clk), .Q(
        \registers[379][6] ) );
  EDFFX1 \registers_reg[379][5]  ( .D(n8318), .E(n677), .CK(clk), .Q(
        \registers[379][5] ) );
  EDFFX1 \registers_reg[379][4]  ( .D(n8260), .E(n677), .CK(clk), .Q(
        \registers[379][4] ) );
  EDFFX1 \registers_reg[379][3]  ( .D(n8202), .E(n677), .CK(clk), .Q(
        \registers[379][3] ) );
  EDFFX1 \registers_reg[379][2]  ( .D(n8723), .E(n677), .CK(clk), .Q(
        \registers[379][2] ) );
  EDFFX1 \registers_reg[379][1]  ( .D(n8695), .E(n677), .CK(clk), .Q(
        \registers[379][1] ) );
  EDFFX1 \registers_reg[379][0]  ( .D(n7995), .E(n677), .CK(clk), .Q(
        \registers[379][0] ) );
  EDFFX1 \registers_reg[375][7]  ( .D(n8432), .E(n673), .CK(clk), .Q(
        \registers[375][7] ) );
  EDFFX1 \registers_reg[375][6]  ( .D(n8374), .E(n673), .CK(clk), .Q(
        \registers[375][6] ) );
  EDFFX1 \registers_reg[375][5]  ( .D(n8316), .E(n673), .CK(clk), .Q(
        \registers[375][5] ) );
  EDFFX1 \registers_reg[375][4]  ( .D(n8258), .E(n673), .CK(clk), .Q(
        \registers[375][4] ) );
  EDFFX1 \registers_reg[375][3]  ( .D(n8200), .E(n673), .CK(clk), .Q(
        \registers[375][3] ) );
  EDFFX1 \registers_reg[375][2]  ( .D(n8734), .E(n673), .CK(clk), .Q(
        \registers[375][2] ) );
  EDFFX1 \registers_reg[375][1]  ( .D(n8706), .E(n673), .CK(clk), .Q(
        \registers[375][1] ) );
  EDFFX1 \registers_reg[375][0]  ( .D(n8031), .E(n673), .CK(clk), .Q(
        \registers[375][0] ) );
  EDFFX1 \registers_reg[371][7]  ( .D(n8433), .E(n669), .CK(clk), .Q(
        \registers[371][7] ) );
  EDFFX1 \registers_reg[371][6]  ( .D(n8375), .E(n669), .CK(clk), .Q(
        \registers[371][6] ) );
  EDFFX1 \registers_reg[371][5]  ( .D(n8317), .E(n669), .CK(clk), .Q(
        \registers[371][5] ) );
  EDFFX1 \registers_reg[371][4]  ( .D(n8259), .E(n669), .CK(clk), .Q(
        \registers[371][4] ) );
  EDFFX1 \registers_reg[371][3]  ( .D(n8201), .E(n669), .CK(clk), .Q(
        \registers[371][3] ) );
  EDFFX1 \registers_reg[371][2]  ( .D(n8133), .E(n669), .CK(clk), .Q(
        \registers[371][2] ) );
  EDFFX1 \registers_reg[371][1]  ( .D(n8077), .E(n669), .CK(clk), .Q(
        \registers[371][1] ) );
  EDFFX1 \registers_reg[371][0]  ( .D(n8047), .E(n669), .CK(clk), .Q(
        \registers[371][0] ) );
  EDFFX1 \registers_reg[367][7]  ( .D(n8434), .E(n665), .CK(clk), .Q(
        \registers[367][7] ) );
  EDFFX1 \registers_reg[367][6]  ( .D(n8376), .E(n665), .CK(clk), .Q(
        \registers[367][6] ) );
  EDFFX1 \registers_reg[367][5]  ( .D(n8318), .E(n665), .CK(clk), .Q(
        \registers[367][5] ) );
  EDFFX1 \registers_reg[367][4]  ( .D(n8260), .E(n665), .CK(clk), .Q(
        \registers[367][4] ) );
  EDFFX1 \registers_reg[367][3]  ( .D(n8197), .E(n665), .CK(clk), .Q(
        \registers[367][3] ) );
  EDFFX1 \registers_reg[367][2]  ( .D(n8725), .E(n665), .CK(clk), .Q(
        \registers[367][2] ) );
  EDFFX1 \registers_reg[367][1]  ( .D(n8697), .E(n665), .CK(clk), .Q(
        \registers[367][1] ) );
  EDFFX1 \registers_reg[367][0]  ( .D(n8046), .E(n665), .CK(clk), .Q(
        \registers[367][0] ) );
  EDFFX1 \registers_reg[363][7]  ( .D(n8433), .E(n661), .CK(clk), .Q(
        \registers[363][7] ) );
  EDFFX1 \registers_reg[363][6]  ( .D(n8375), .E(n661), .CK(clk), .Q(
        \registers[363][6] ) );
  EDFFX1 \registers_reg[363][5]  ( .D(n8317), .E(n661), .CK(clk), .Q(
        \registers[363][5] ) );
  EDFFX1 \registers_reg[363][4]  ( .D(n8259), .E(n661), .CK(clk), .Q(
        \registers[363][4] ) );
  EDFFX1 \registers_reg[363][3]  ( .D(n8198), .E(n661), .CK(clk), .Q(
        \registers[363][3] ) );
  EDFFX1 \registers_reg[363][2]  ( .D(n8130), .E(n661), .CK(clk), .Q(
        \registers[363][2] ) );
  EDFFX1 \registers_reg[363][1]  ( .D(n8074), .E(n661), .CK(clk), .Q(
        \registers[363][1] ) );
  EDFFX1 \registers_reg[363][0]  ( .D(n8047), .E(n661), .CK(clk), .Q(
        \registers[363][0] ) );
  EDFFX1 \registers_reg[359][7]  ( .D(n8433), .E(n994), .CK(clk), .Q(
        \registers[359][7] ) );
  EDFFX1 \registers_reg[359][6]  ( .D(n8375), .E(n994), .CK(clk), .Q(
        \registers[359][6] ) );
  EDFFX1 \registers_reg[359][5]  ( .D(n8317), .E(n994), .CK(clk), .Q(
        \registers[359][5] ) );
  EDFFX1 \registers_reg[359][4]  ( .D(n8259), .E(n994), .CK(clk), .Q(
        \registers[359][4] ) );
  EDFFX1 \registers_reg[359][3]  ( .D(n8199), .E(n994), .CK(clk), .Q(
        \registers[359][3] ) );
  EDFFX1 \registers_reg[359][2]  ( .D(n8134), .E(n994), .CK(clk), .Q(
        \registers[359][2] ) );
  EDFFX1 \registers_reg[359][1]  ( .D(n8078), .E(n994), .CK(clk), .Q(
        \registers[359][1] ) );
  EDFFX1 \registers_reg[359][0]  ( .D(n8048), .E(n994), .CK(clk), .Q(
        \registers[359][0] ) );
  EDFFX1 \registers_reg[355][7]  ( .D(n8434), .E(n990), .CK(clk), .Q(
        \registers[355][7] ) );
  EDFFX1 \registers_reg[355][6]  ( .D(n8376), .E(n990), .CK(clk), .Q(
        \registers[355][6] ) );
  EDFFX1 \registers_reg[355][5]  ( .D(n8318), .E(n990), .CK(clk), .Q(
        \registers[355][5] ) );
  EDFFX1 \registers_reg[355][4]  ( .D(n8260), .E(n990), .CK(clk), .Q(
        \registers[355][4] ) );
  EDFFX1 \registers_reg[355][3]  ( .D(n8167), .E(n990), .CK(clk), .Q(
        \registers[355][3] ) );
  EDFFX1 \registers_reg[355][2]  ( .D(n8738), .E(n990), .CK(clk), .Q(
        \registers[355][2] ) );
  EDFFX1 \registers_reg[355][1]  ( .D(n8710), .E(n990), .CK(clk), .Q(
        \registers[355][1] ) );
  EDFFX1 \registers_reg[355][0]  ( .D(n8046), .E(n990), .CK(clk), .Q(
        \registers[355][0] ) );
  EDFFX1 \registers_reg[351][7]  ( .D(n8430), .E(n657), .CK(clk), .Q(
        \registers[351][7] ) );
  EDFFX1 \registers_reg[351][6]  ( .D(n8372), .E(n657), .CK(clk), .Q(
        \registers[351][6] ) );
  EDFFX1 \registers_reg[351][5]  ( .D(n8314), .E(n657), .CK(clk), .Q(
        \registers[351][5] ) );
  EDFFX1 \registers_reg[351][4]  ( .D(n8256), .E(n657), .CK(clk), .Q(
        \registers[351][4] ) );
  EDFFX1 \registers_reg[351][3]  ( .D(n8184), .E(n657), .CK(clk), .Q(
        \registers[351][3] ) );
  EDFFX1 \registers_reg[351][2]  ( .D(n8131), .E(n657), .CK(clk), .Q(
        \registers[351][2] ) );
  EDFFX1 \registers_reg[351][1]  ( .D(n8075), .E(n657), .CK(clk), .Q(
        \registers[351][1] ) );
  EDFFX1 \registers_reg[351][0]  ( .D(n8047), .E(n657), .CK(clk), .Q(
        \registers[351][0] ) );
  EDFFX1 \registers_reg[347][7]  ( .D(n8431), .E(n653), .CK(clk), .Q(
        \registers[347][7] ) );
  EDFFX1 \registers_reg[347][6]  ( .D(n8373), .E(n653), .CK(clk), .Q(
        \registers[347][6] ) );
  EDFFX1 \registers_reg[347][5]  ( .D(n8315), .E(n653), .CK(clk), .Q(
        \registers[347][5] ) );
  EDFFX1 \registers_reg[347][4]  ( .D(n8257), .E(n653), .CK(clk), .Q(
        \registers[347][4] ) );
  EDFFX1 \registers_reg[347][3]  ( .D(n8196), .E(n653), .CK(clk), .Q(
        \registers[347][3] ) );
  EDFFX1 \registers_reg[347][2]  ( .D(n8143), .E(n653), .CK(clk), .Q(
        \registers[347][2] ) );
  EDFFX1 \registers_reg[347][1]  ( .D(n8087), .E(n653), .CK(clk), .Q(
        \registers[347][1] ) );
  EDFFX1 \registers_reg[347][0]  ( .D(n8048), .E(n653), .CK(clk), .Q(
        \registers[347][0] ) );
  EDFFX1 \registers_reg[343][7]  ( .D(n8432), .E(n649), .CK(clk), .Q(
        \registers[343][7] ) );
  EDFFX1 \registers_reg[343][6]  ( .D(n8374), .E(n649), .CK(clk), .Q(
        \registers[343][6] ) );
  EDFFX1 \registers_reg[343][5]  ( .D(n8316), .E(n649), .CK(clk), .Q(
        \registers[343][5] ) );
  EDFFX1 \registers_reg[343][4]  ( .D(n8258), .E(n649), .CK(clk), .Q(
        \registers[343][4] ) );
  EDFFX1 \registers_reg[343][3]  ( .D(n8168), .E(n649), .CK(clk), .Q(
        \registers[343][3] ) );
  EDFFX1 \registers_reg[343][2]  ( .D(n8737), .E(n649), .CK(clk), .Q(
        \registers[343][2] ) );
  EDFFX1 \registers_reg[343][1]  ( .D(n8709), .E(n649), .CK(clk), .Q(
        \registers[343][1] ) );
  EDFFX1 \registers_reg[343][0]  ( .D(n8046), .E(n649), .CK(clk), .Q(
        \registers[343][0] ) );
  EDFFX1 \registers_reg[339][7]  ( .D(n8430), .E(n645), .CK(clk), .Q(
        \registers[339][7] ) );
  EDFFX1 \registers_reg[339][6]  ( .D(n8372), .E(n645), .CK(clk), .Q(
        \registers[339][6] ) );
  EDFFX1 \registers_reg[339][5]  ( .D(n8314), .E(n645), .CK(clk), .Q(
        \registers[339][5] ) );
  EDFFX1 \registers_reg[339][4]  ( .D(n8256), .E(n645), .CK(clk), .Q(
        \registers[339][4] ) );
  EDFFX1 \registers_reg[339][3]  ( .D(n8182), .E(n645), .CK(clk), .Q(
        \registers[339][3] ) );
  EDFFX1 \registers_reg[339][2]  ( .D(n8123), .E(n645), .CK(clk), .Q(
        \registers[339][2] ) );
  EDFFX1 \registers_reg[339][1]  ( .D(n8067), .E(n645), .CK(clk), .Q(
        \registers[339][1] ) );
  EDFFX1 \registers_reg[339][0]  ( .D(n8047), .E(n645), .CK(clk), .Q(
        \registers[339][0] ) );
  EDFFX1 \registers_reg[335][7]  ( .D(n8431), .E(n641), .CK(clk), .Q(
        \registers[335][7] ) );
  EDFFX1 \registers_reg[335][6]  ( .D(n8373), .E(n641), .CK(clk), .Q(
        \registers[335][6] ) );
  EDFFX1 \registers_reg[335][5]  ( .D(n8315), .E(n641), .CK(clk), .Q(
        \registers[335][5] ) );
  EDFFX1 \registers_reg[335][4]  ( .D(n8257), .E(n641), .CK(clk), .Q(
        \registers[335][4] ) );
  EDFFX1 \registers_reg[335][3]  ( .D(n8191), .E(n641), .CK(clk), .Q(
        \registers[335][3] ) );
  EDFFX1 \registers_reg[335][2]  ( .D(n8141), .E(n641), .CK(clk), .Q(
        \registers[335][2] ) );
  EDFFX1 \registers_reg[335][1]  ( .D(n8085), .E(n641), .CK(clk), .Q(
        \registers[335][1] ) );
  EDFFX1 \registers_reg[335][0]  ( .D(n8048), .E(n641), .CK(clk), .Q(
        \registers[335][0] ) );
  EDFFX1 \registers_reg[331][7]  ( .D(n8432), .E(n637), .CK(clk), .Q(
        \registers[331][7] ) );
  EDFFX1 \registers_reg[331][6]  ( .D(n8374), .E(n637), .CK(clk), .Q(
        \registers[331][6] ) );
  EDFFX1 \registers_reg[331][5]  ( .D(n8316), .E(n637), .CK(clk), .Q(
        \registers[331][5] ) );
  EDFFX1 \registers_reg[331][4]  ( .D(n8258), .E(n637), .CK(clk), .Q(
        \registers[331][4] ) );
  EDFFX1 \registers_reg[331][3]  ( .D(n8169), .E(n637), .CK(clk), .Q(
        \registers[331][3] ) );
  EDFFX1 \registers_reg[331][2]  ( .D(n8156), .E(n637), .CK(clk), .Q(
        \registers[331][2] ) );
  EDFFX1 \registers_reg[331][1]  ( .D(n8100), .E(n637), .CK(clk), .Q(
        \registers[331][1] ) );
  EDFFX1 \registers_reg[331][0]  ( .D(n8046), .E(n637), .CK(clk), .Q(
        \registers[331][0] ) );
  EDFFX1 \registers_reg[327][7]  ( .D(n8430), .E(n987), .CK(clk), .Q(
        \registers[327][7] ) );
  EDFFX1 \registers_reg[327][6]  ( .D(n8372), .E(n987), .CK(clk), .Q(
        \registers[327][6] ) );
  EDFFX1 \registers_reg[327][5]  ( .D(n8314), .E(n987), .CK(clk), .Q(
        \registers[327][5] ) );
  EDFFX1 \registers_reg[327][4]  ( .D(n8256), .E(n987), .CK(clk), .Q(
        \registers[327][4] ) );
  EDFFX1 \registers_reg[327][3]  ( .D(n8183), .E(n987), .CK(clk), .Q(
        \registers[327][3] ) );
  EDFFX1 \registers_reg[327][2]  ( .D(n8124), .E(n987), .CK(clk), .Q(
        \registers[327][2] ) );
  EDFFX1 \registers_reg[327][1]  ( .D(n8068), .E(n987), .CK(clk), .Q(
        \registers[327][1] ) );
  EDFFX1 \registers_reg[327][0]  ( .D(n8047), .E(n987), .CK(clk), .Q(
        \registers[327][0] ) );
  EDFFX1 \registers_reg[323][7]  ( .D(n8431), .E(n983), .CK(clk), .Q(
        \registers[323][7] ) );
  EDFFX1 \registers_reg[323][6]  ( .D(n8373), .E(n983), .CK(clk), .Q(
        \registers[323][6] ) );
  EDFFX1 \registers_reg[323][5]  ( .D(n8315), .E(n983), .CK(clk), .Q(
        \registers[323][5] ) );
  EDFFX1 \registers_reg[323][4]  ( .D(n8257), .E(n983), .CK(clk), .Q(
        \registers[323][4] ) );
  EDFFX1 \registers_reg[323][3]  ( .D(n8192), .E(n983), .CK(clk), .Q(
        \registers[323][3] ) );
  EDFFX1 \registers_reg[323][2]  ( .D(n8142), .E(n983), .CK(clk), .Q(
        \registers[323][2] ) );
  EDFFX1 \registers_reg[323][1]  ( .D(n8086), .E(n983), .CK(clk), .Q(
        \registers[323][1] ) );
  EDFFX1 \registers_reg[323][0]  ( .D(n8048), .E(n983), .CK(clk), .Q(
        \registers[323][0] ) );
  EDFFX1 \registers_reg[319][7]  ( .D(n8430), .E(n633), .CK(clk), .Q(
        \registers[319][7] ) );
  EDFFX1 \registers_reg[319][6]  ( .D(n8372), .E(n633), .CK(clk), .Q(
        \registers[319][6] ) );
  EDFFX1 \registers_reg[319][5]  ( .D(n8314), .E(n633), .CK(clk), .Q(
        \registers[319][5] ) );
  EDFFX1 \registers_reg[319][4]  ( .D(n8256), .E(n633), .CK(clk), .Q(
        \registers[319][4] ) );
  EDFFX1 \registers_reg[319][3]  ( .D(n8179), .E(n633), .CK(clk), .Q(
        \registers[319][3] ) );
  EDFFX1 \registers_reg[319][2]  ( .D(n8160), .E(n633), .CK(clk), .Q(
        \registers[319][2] ) );
  EDFFX1 \registers_reg[319][1]  ( .D(n8104), .E(n633), .CK(clk), .Q(
        \registers[319][1] ) );
  EDFFX1 \registers_reg[319][0]  ( .D(n8044), .E(n633), .CK(clk), .Q(
        \registers[319][0] ) );
  EDFFX1 \registers_reg[315][7]  ( .D(n8431), .E(n629), .CK(clk), .Q(
        \registers[315][7] ) );
  EDFFX1 \registers_reg[315][6]  ( .D(n8373), .E(n629), .CK(clk), .Q(
        \registers[315][6] ) );
  EDFFX1 \registers_reg[315][5]  ( .D(n8315), .E(n629), .CK(clk), .Q(
        \registers[315][5] ) );
  EDFFX1 \registers_reg[315][4]  ( .D(n8257), .E(n629), .CK(clk), .Q(
        \registers[315][4] ) );
  EDFFX1 \registers_reg[315][3]  ( .D(n8193), .E(n629), .CK(clk), .Q(
        \registers[315][3] ) );
  EDFFX1 \registers_reg[315][2]  ( .D(n8158), .E(n629), .CK(clk), .Q(
        \registers[315][2] ) );
  EDFFX1 \registers_reg[315][1]  ( .D(n8102), .E(n629), .CK(clk), .Q(
        \registers[315][1] ) );
  EDFFX1 \registers_reg[315][0]  ( .D(n8045), .E(n629), .CK(clk), .Q(
        \registers[315][0] ) );
  EDFFX1 \registers_reg[311][7]  ( .D(n8432), .E(n625), .CK(clk), .Q(
        \registers[311][7] ) );
  EDFFX1 \registers_reg[311][6]  ( .D(n8374), .E(n625), .CK(clk), .Q(
        \registers[311][6] ) );
  EDFFX1 \registers_reg[311][5]  ( .D(n8316), .E(n625), .CK(clk), .Q(
        \registers[311][5] ) );
  EDFFX1 \registers_reg[311][4]  ( .D(n8258), .E(n625), .CK(clk), .Q(
        \registers[311][4] ) );
  EDFFX1 \registers_reg[311][3]  ( .D(n8166), .E(n625), .CK(clk), .Q(
        \registers[311][3] ) );
  EDFFX1 \registers_reg[311][2]  ( .D(n8159), .E(n625), .CK(clk), .Q(
        \registers[311][2] ) );
  EDFFX1 \registers_reg[311][1]  ( .D(n8103), .E(n625), .CK(clk), .Q(
        \registers[311][1] ) );
  EDFFX1 \registers_reg[311][0]  ( .D(n8043), .E(n625), .CK(clk), .Q(
        \registers[311][0] ) );
  EDFFX1 \registers_reg[307][7]  ( .D(n8430), .E(n621), .CK(clk), .Q(
        \registers[307][7] ) );
  EDFFX1 \registers_reg[307][6]  ( .D(n8372), .E(n621), .CK(clk), .Q(
        \registers[307][6] ) );
  EDFFX1 \registers_reg[307][5]  ( .D(n8314), .E(n621), .CK(clk), .Q(
        \registers[307][5] ) );
  EDFFX1 \registers_reg[307][4]  ( .D(n8256), .E(n621), .CK(clk), .Q(
        \registers[307][4] ) );
  EDFFX1 \registers_reg[307][3]  ( .D(n8180), .E(n621), .CK(clk), .Q(
        \registers[307][3] ) );
  EDFFX1 \registers_reg[307][2]  ( .D(n8160), .E(n621), .CK(clk), .Q(
        \registers[307][2] ) );
  EDFFX1 \registers_reg[307][1]  ( .D(n8104), .E(n621), .CK(clk), .Q(
        \registers[307][1] ) );
  EDFFX1 \registers_reg[307][0]  ( .D(n8044), .E(n621), .CK(clk), .Q(
        \registers[307][0] ) );
  EDFFX1 \registers_reg[303][7]  ( .D(n8431), .E(n617), .CK(clk), .Q(
        \registers[303][7] ) );
  EDFFX1 \registers_reg[303][6]  ( .D(n8373), .E(n617), .CK(clk), .Q(
        \registers[303][6] ) );
  EDFFX1 \registers_reg[303][5]  ( .D(n8315), .E(n617), .CK(clk), .Q(
        \registers[303][5] ) );
  EDFFX1 \registers_reg[303][4]  ( .D(n8257), .E(n617), .CK(clk), .Q(
        \registers[303][4] ) );
  EDFFX1 \registers_reg[303][3]  ( .D(n8202), .E(n617), .CK(clk), .Q(
        \registers[303][3] ) );
  EDFFX1 \registers_reg[303][2]  ( .D(n8158), .E(n617), .CK(clk), .Q(
        \registers[303][2] ) );
  EDFFX1 \registers_reg[303][1]  ( .D(n8102), .E(n617), .CK(clk), .Q(
        \registers[303][1] ) );
  EDFFX1 \registers_reg[303][0]  ( .D(n8045), .E(n617), .CK(clk), .Q(
        \registers[303][0] ) );
  EDFFX1 \registers_reg[299][7]  ( .D(n8428), .E(n613), .CK(clk), .Q(
        \registers[299][7] ) );
  EDFFX1 \registers_reg[299][6]  ( .D(n8370), .E(n613), .CK(clk), .Q(
        \registers[299][6] ) );
  EDFFX1 \registers_reg[299][5]  ( .D(n8312), .E(n613), .CK(clk), .Q(
        \registers[299][5] ) );
  EDFFX1 \registers_reg[299][4]  ( .D(n8254), .E(n613), .CK(clk), .Q(
        \registers[299][4] ) );
  EDFFX1 \registers_reg[299][3]  ( .D(n8164), .E(n613), .CK(clk), .Q(
        \registers[299][3] ) );
  EDFFX1 \registers_reg[299][2]  ( .D(n8159), .E(n613), .CK(clk), .Q(
        \registers[299][2] ) );
  EDFFX1 \registers_reg[299][1]  ( .D(n8103), .E(n613), .CK(clk), .Q(
        \registers[299][1] ) );
  EDFFX1 \registers_reg[299][0]  ( .D(n8043), .E(n613), .CK(clk), .Q(
        \registers[299][0] ) );
  EDFFX1 \registers_reg[295][7]  ( .D(n8429), .E(n980), .CK(clk), .Q(
        \registers[295][7] ) );
  EDFFX1 \registers_reg[295][6]  ( .D(n8371), .E(n980), .CK(clk), .Q(
        \registers[295][6] ) );
  EDFFX1 \registers_reg[295][5]  ( .D(n8313), .E(n980), .CK(clk), .Q(
        \registers[295][5] ) );
  EDFFX1 \registers_reg[295][4]  ( .D(n8255), .E(n980), .CK(clk), .Q(
        \registers[295][4] ) );
  EDFFX1 \registers_reg[295][3]  ( .D(n8200), .E(n980), .CK(clk), .Q(
        \registers[295][3] ) );
  EDFFX1 \registers_reg[295][2]  ( .D(n8160), .E(n980), .CK(clk), .Q(
        \registers[295][2] ) );
  EDFFX1 \registers_reg[295][1]  ( .D(n8104), .E(n980), .CK(clk), .Q(
        \registers[295][1] ) );
  EDFFX1 \registers_reg[295][0]  ( .D(n8044), .E(n980), .CK(clk), .Q(
        \registers[295][0] ) );
  EDFFX1 \registers_reg[291][7]  ( .D(n8411), .E(n976), .CK(clk), .Q(
        \registers[291][7] ) );
  EDFFX1 \registers_reg[291][6]  ( .D(n8353), .E(n976), .CK(clk), .Q(
        \registers[291][6] ) );
  EDFFX1 \registers_reg[291][5]  ( .D(n8295), .E(n976), .CK(clk), .Q(
        \registers[291][5] ) );
  EDFFX1 \registers_reg[291][4]  ( .D(n8237), .E(n976), .CK(clk), .Q(
        \registers[291][4] ) );
  EDFFX1 \registers_reg[291][3]  ( .D(n8201), .E(n976), .CK(clk), .Q(
        \registers[291][3] ) );
  EDFFX1 \registers_reg[291][2]  ( .D(n8158), .E(n976), .CK(clk), .Q(
        \registers[291][2] ) );
  EDFFX1 \registers_reg[291][1]  ( .D(n8102), .E(n976), .CK(clk), .Q(
        \registers[291][1] ) );
  EDFFX1 \registers_reg[291][0]  ( .D(n8045), .E(n976), .CK(clk), .Q(
        \registers[291][0] ) );
  EDFFX1 \registers_reg[287][7]  ( .D(n8428), .E(n609), .CK(clk), .Q(
        \registers[287][7] ) );
  EDFFX1 \registers_reg[287][6]  ( .D(n8370), .E(n609), .CK(clk), .Q(
        \registers[287][6] ) );
  EDFFX1 \registers_reg[287][5]  ( .D(n8312), .E(n609), .CK(clk), .Q(
        \registers[287][5] ) );
  EDFFX1 \registers_reg[287][4]  ( .D(n8254), .E(n609), .CK(clk), .Q(
        \registers[287][4] ) );
  EDFFX1 \registers_reg[287][3]  ( .D(n8202), .E(n609), .CK(clk), .Q(
        \registers[287][3] ) );
  EDFFX1 \registers_reg[287][2]  ( .D(n8159), .E(n609), .CK(clk), .Q(
        \registers[287][2] ) );
  EDFFX1 \registers_reg[287][1]  ( .D(n8103), .E(n609), .CK(clk), .Q(
        \registers[287][1] ) );
  EDFFX1 \registers_reg[287][0]  ( .D(n8043), .E(n609), .CK(clk), .Q(
        \registers[287][0] ) );
  EDFFX1 \registers_reg[283][7]  ( .D(n8429), .E(n605), .CK(clk), .Q(
        \registers[283][7] ) );
  EDFFX1 \registers_reg[283][6]  ( .D(n8371), .E(n605), .CK(clk), .Q(
        \registers[283][6] ) );
  EDFFX1 \registers_reg[283][5]  ( .D(n8313), .E(n605), .CK(clk), .Q(
        \registers[283][5] ) );
  EDFFX1 \registers_reg[283][4]  ( .D(n8255), .E(n605), .CK(clk), .Q(
        \registers[283][4] ) );
  EDFFX1 \registers_reg[283][3]  ( .D(n8200), .E(n605), .CK(clk), .Q(
        \registers[283][3] ) );
  EDFFX1 \registers_reg[283][2]  ( .D(n8160), .E(n605), .CK(clk), .Q(
        \registers[283][2] ) );
  EDFFX1 \registers_reg[283][1]  ( .D(n8104), .E(n605), .CK(clk), .Q(
        \registers[283][1] ) );
  EDFFX1 \registers_reg[283][0]  ( .D(n8044), .E(n605), .CK(clk), .Q(
        \registers[283][0] ) );
  EDFFX1 \registers_reg[279][7]  ( .D(n8410), .E(n601), .CK(clk), .Q(
        \registers[279][7] ) );
  EDFFX1 \registers_reg[279][6]  ( .D(n8352), .E(n601), .CK(clk), .Q(
        \registers[279][6] ) );
  EDFFX1 \registers_reg[279][5]  ( .D(n8294), .E(n601), .CK(clk), .Q(
        \registers[279][5] ) );
  EDFFX1 \registers_reg[279][4]  ( .D(n8236), .E(n601), .CK(clk), .Q(
        \registers[279][4] ) );
  EDFFX1 \registers_reg[279][3]  ( .D(n8201), .E(n601), .CK(clk), .Q(
        \registers[279][3] ) );
  EDFFX1 \registers_reg[279][2]  ( .D(n8158), .E(n601), .CK(clk), .Q(
        \registers[279][2] ) );
  EDFFX1 \registers_reg[279][1]  ( .D(n8102), .E(n601), .CK(clk), .Q(
        \registers[279][1] ) );
  EDFFX1 \registers_reg[279][0]  ( .D(n8045), .E(n601), .CK(clk), .Q(
        \registers[279][0] ) );
  EDFFX1 \registers_reg[275][7]  ( .D(n8428), .E(n597), .CK(clk), .Q(
        \registers[275][7] ) );
  EDFFX1 \registers_reg[275][6]  ( .D(n8370), .E(n597), .CK(clk), .Q(
        \registers[275][6] ) );
  EDFFX1 \registers_reg[275][5]  ( .D(n8312), .E(n597), .CK(clk), .Q(
        \registers[275][5] ) );
  EDFFX1 \registers_reg[275][4]  ( .D(n8254), .E(n597), .CK(clk), .Q(
        \registers[275][4] ) );
  EDFFX1 \registers_reg[275][3]  ( .D(n8202), .E(n597), .CK(clk), .Q(
        \registers[275][3] ) );
  EDFFX1 \registers_reg[275][2]  ( .D(n8159), .E(n597), .CK(clk), .Q(
        \registers[275][2] ) );
  EDFFX1 \registers_reg[275][1]  ( .D(n8103), .E(n597), .CK(clk), .Q(
        \registers[275][1] ) );
  EDFFX1 \registers_reg[275][0]  ( .D(n8043), .E(n597), .CK(clk), .Q(
        \registers[275][0] ) );
  EDFFX1 \registers_reg[271][7]  ( .D(n8429), .E(n593), .CK(clk), .Q(
        \registers[271][7] ) );
  EDFFX1 \registers_reg[271][6]  ( .D(n8371), .E(n593), .CK(clk), .Q(
        \registers[271][6] ) );
  EDFFX1 \registers_reg[271][5]  ( .D(n8313), .E(n593), .CK(clk), .Q(
        \registers[271][5] ) );
  EDFFX1 \registers_reg[271][4]  ( .D(n8255), .E(n593), .CK(clk), .Q(
        \registers[271][4] ) );
  EDFFX1 \registers_reg[271][3]  ( .D(n8200), .E(n593), .CK(clk), .Q(
        \registers[271][3] ) );
  EDFFX1 \registers_reg[271][2]  ( .D(n8160), .E(n593), .CK(clk), .Q(
        \registers[271][2] ) );
  EDFFX1 \registers_reg[271][1]  ( .D(n8104), .E(n593), .CK(clk), .Q(
        \registers[271][1] ) );
  EDFFX1 \registers_reg[271][0]  ( .D(n8044), .E(n593), .CK(clk), .Q(
        \registers[271][0] ) );
  EDFFX1 \registers_reg[267][7]  ( .D(n8433), .E(n589), .CK(clk), .Q(
        \registers[267][7] ) );
  EDFFX1 \registers_reg[267][6]  ( .D(n8375), .E(n589), .CK(clk), .Q(
        \registers[267][6] ) );
  EDFFX1 \registers_reg[267][5]  ( .D(n8317), .E(n589), .CK(clk), .Q(
        \registers[267][5] ) );
  EDFFX1 \registers_reg[267][4]  ( .D(n8259), .E(n589), .CK(clk), .Q(
        \registers[267][4] ) );
  EDFFX1 \registers_reg[267][3]  ( .D(n8201), .E(n589), .CK(clk), .Q(
        \registers[267][3] ) );
  EDFFX1 \registers_reg[267][2]  ( .D(n8155), .E(n589), .CK(clk), .Q(
        \registers[267][2] ) );
  EDFFX1 \registers_reg[267][1]  ( .D(n8099), .E(n589), .CK(clk), .Q(
        \registers[267][1] ) );
  EDFFX1 \registers_reg[267][0]  ( .D(n8042), .E(n589), .CK(clk), .Q(
        \registers[267][0] ) );
  EDFFX1 \registers_reg[263][7]  ( .D(n8428), .E(n973), .CK(clk), .Q(
        \registers[263][7] ) );
  EDFFX1 \registers_reg[263][6]  ( .D(n8370), .E(n973), .CK(clk), .Q(
        \registers[263][6] ) );
  EDFFX1 \registers_reg[263][5]  ( .D(n8312), .E(n973), .CK(clk), .Q(
        \registers[263][5] ) );
  EDFFX1 \registers_reg[263][4]  ( .D(n8254), .E(n973), .CK(clk), .Q(
        \registers[263][4] ) );
  EDFFX1 \registers_reg[263][3]  ( .D(n8202), .E(n973), .CK(clk), .Q(
        \registers[263][3] ) );
  EDFFX1 \registers_reg[263][2]  ( .D(n8156), .E(n973), .CK(clk), .Q(
        \registers[263][2] ) );
  EDFFX1 \registers_reg[263][1]  ( .D(n8100), .E(n973), .CK(clk), .Q(
        \registers[263][1] ) );
  EDFFX1 \registers_reg[263][0]  ( .D(n8040), .E(n973), .CK(clk), .Q(
        \registers[263][0] ) );
  EDFFX1 \registers_reg[259][7]  ( .D(n8429), .E(n969), .CK(clk), .Q(
        \registers[259][7] ) );
  EDFFX1 \registers_reg[259][6]  ( .D(n8371), .E(n969), .CK(clk), .Q(
        \registers[259][6] ) );
  EDFFX1 \registers_reg[259][5]  ( .D(n8313), .E(n969), .CK(clk), .Q(
        \registers[259][5] ) );
  EDFFX1 \registers_reg[259][4]  ( .D(n8255), .E(n969), .CK(clk), .Q(
        \registers[259][4] ) );
  EDFFX1 \registers_reg[259][3]  ( .D(n8200), .E(n969), .CK(clk), .Q(
        \registers[259][3] ) );
  EDFFX1 \registers_reg[259][2]  ( .D(n8157), .E(n969), .CK(clk), .Q(
        \registers[259][2] ) );
  EDFFX1 \registers_reg[259][1]  ( .D(n8101), .E(n969), .CK(clk), .Q(
        \registers[259][1] ) );
  EDFFX1 \registers_reg[259][0]  ( .D(n8041), .E(n969), .CK(clk), .Q(
        \registers[259][0] ) );
  EDFFX1 \registers_reg[255][7]  ( .D(n8412), .E(n585), .CK(clk), .Q(
        \registers[255][7] ) );
  EDFFX1 \registers_reg[255][6]  ( .D(n8354), .E(n585), .CK(clk), .Q(
        \registers[255][6] ) );
  EDFFX1 \registers_reg[255][5]  ( .D(n8296), .E(n585), .CK(clk), .Q(
        \registers[255][5] ) );
  EDFFX1 \registers_reg[255][4]  ( .D(n8238), .E(n585), .CK(clk), .Q(
        \registers[255][4] ) );
  EDFFX1 \registers_reg[255][3]  ( .D(n8189), .E(n585), .CK(clk), .Q(
        \registers[255][3] ) );
  EDFFX1 \registers_reg[255][2]  ( .D(n8141), .E(n585), .CK(clk), .Q(
        \registers[255][2] ) );
  EDFFX1 \registers_reg[255][1]  ( .D(n8085), .E(n585), .CK(clk), .Q(
        \registers[255][1] ) );
  EDFFX1 \registers_reg[255][0]  ( .D(n8027), .E(n585), .CK(clk), .Q(
        \registers[255][0] ) );
  EDFFX1 \registers_reg[251][7]  ( .D(n8410), .E(n581), .CK(clk), .Q(
        \registers[251][7] ) );
  EDFFX1 \registers_reg[251][6]  ( .D(n8352), .E(n581), .CK(clk), .Q(
        \registers[251][6] ) );
  EDFFX1 \registers_reg[251][5]  ( .D(n8294), .E(n581), .CK(clk), .Q(
        \registers[251][5] ) );
  EDFFX1 \registers_reg[251][4]  ( .D(n8236), .E(n581), .CK(clk), .Q(
        \registers[251][4] ) );
  EDFFX1 \registers_reg[251][3]  ( .D(n8190), .E(n581), .CK(clk), .Q(
        \registers[251][3] ) );
  EDFFX1 \registers_reg[251][2]  ( .D(n8142), .E(n581), .CK(clk), .Q(
        \registers[251][2] ) );
  EDFFX1 \registers_reg[251][1]  ( .D(n8086), .E(n581), .CK(clk), .Q(
        \registers[251][1] ) );
  EDFFX1 \registers_reg[251][0]  ( .D(n8025), .E(n581), .CK(clk), .Q(
        \registers[251][0] ) );
  EDFFX1 \registers_reg[247][7]  ( .D(n8411), .E(n577), .CK(clk), .Q(
        \registers[247][7] ) );
  EDFFX1 \registers_reg[247][6]  ( .D(n8353), .E(n577), .CK(clk), .Q(
        \registers[247][6] ) );
  EDFFX1 \registers_reg[247][5]  ( .D(n8295), .E(n577), .CK(clk), .Q(
        \registers[247][5] ) );
  EDFFX1 \registers_reg[247][4]  ( .D(n8237), .E(n577), .CK(clk), .Q(
        \registers[247][4] ) );
  EDFFX1 \registers_reg[247][3]  ( .D(n8188), .E(n577), .CK(clk), .Q(
        \registers[247][3] ) );
  EDFFX1 \registers_reg[247][2]  ( .D(n8143), .E(n577), .CK(clk), .Q(
        \registers[247][2] ) );
  EDFFX1 \registers_reg[247][1]  ( .D(n8087), .E(n577), .CK(clk), .Q(
        \registers[247][1] ) );
  EDFFX1 \registers_reg[247][0]  ( .D(n8026), .E(n577), .CK(clk), .Q(
        \registers[247][0] ) );
  EDFFX1 \registers_reg[243][7]  ( .D(n8412), .E(n573), .CK(clk), .Q(
        \registers[243][7] ) );
  EDFFX1 \registers_reg[243][6]  ( .D(n8354), .E(n573), .CK(clk), .Q(
        \registers[243][6] ) );
  EDFFX1 \registers_reg[243][5]  ( .D(n8296), .E(n573), .CK(clk), .Q(
        \registers[243][5] ) );
  EDFFX1 \registers_reg[243][4]  ( .D(n8238), .E(n573), .CK(clk), .Q(
        \registers[243][4] ) );
  EDFFX1 \registers_reg[243][3]  ( .D(n8189), .E(n573), .CK(clk), .Q(
        \registers[243][3] ) );
  EDFFX1 \registers_reg[243][2]  ( .D(n8141), .E(n573), .CK(clk), .Q(
        \registers[243][2] ) );
  EDFFX1 \registers_reg[243][1]  ( .D(n8085), .E(n573), .CK(clk), .Q(
        \registers[243][1] ) );
  EDFFX1 \registers_reg[243][0]  ( .D(n8027), .E(n573), .CK(clk), .Q(
        \registers[243][0] ) );
  EDFFX1 \registers_reg[239][7]  ( .D(n8410), .E(n569), .CK(clk), .Q(
        \registers[239][7] ) );
  EDFFX1 \registers_reg[239][6]  ( .D(n8352), .E(n569), .CK(clk), .Q(
        \registers[239][6] ) );
  EDFFX1 \registers_reg[239][5]  ( .D(n8294), .E(n569), .CK(clk), .Q(
        \registers[239][5] ) );
  EDFFX1 \registers_reg[239][4]  ( .D(n8236), .E(n569), .CK(clk), .Q(
        \registers[239][4] ) );
  EDFFX1 \registers_reg[239][3]  ( .D(n8190), .E(n569), .CK(clk), .Q(
        \registers[239][3] ) );
  EDFFX1 \registers_reg[239][2]  ( .D(n8142), .E(n569), .CK(clk), .Q(
        \registers[239][2] ) );
  EDFFX1 \registers_reg[239][1]  ( .D(n8086), .E(n569), .CK(clk), .Q(
        \registers[239][1] ) );
  EDFFX1 \registers_reg[239][0]  ( .D(n8025), .E(n569), .CK(clk), .Q(
        \registers[239][0] ) );
  EDFFX1 \registers_reg[235][7]  ( .D(n8411), .E(n565), .CK(clk), .Q(
        \registers[235][7] ) );
  EDFFX1 \registers_reg[235][6]  ( .D(n8353), .E(n565), .CK(clk), .Q(
        \registers[235][6] ) );
  EDFFX1 \registers_reg[235][5]  ( .D(n8295), .E(n565), .CK(clk), .Q(
        \registers[235][5] ) );
  EDFFX1 \registers_reg[235][4]  ( .D(n8237), .E(n565), .CK(clk), .Q(
        \registers[235][4] ) );
  EDFFX1 \registers_reg[235][3]  ( .D(n8185), .E(n565), .CK(clk), .Q(
        \registers[235][3] ) );
  EDFFX1 \registers_reg[235][2]  ( .D(n8143), .E(n565), .CK(clk), .Q(
        \registers[235][2] ) );
  EDFFX1 \registers_reg[235][1]  ( .D(n8087), .E(n565), .CK(clk), .Q(
        \registers[235][1] ) );
  EDFFX1 \registers_reg[235][0]  ( .D(n8026), .E(n565), .CK(clk), .Q(
        \registers[235][0] ) );
  EDFFX1 \registers_reg[231][7]  ( .D(n8412), .E(n1033), .CK(clk), .Q(
        \registers[231][7] ) );
  EDFFX1 \registers_reg[231][6]  ( .D(n8354), .E(n1033), .CK(clk), .Q(
        \registers[231][6] ) );
  EDFFX1 \registers_reg[231][5]  ( .D(n8296), .E(n1033), .CK(clk), .Q(
        \registers[231][5] ) );
  EDFFX1 \registers_reg[231][4]  ( .D(n8238), .E(n1033), .CK(clk), .Q(
        \registers[231][4] ) );
  EDFFX1 \registers_reg[231][3]  ( .D(n8186), .E(n1033), .CK(clk), .Q(
        \registers[231][3] ) );
  EDFFX1 \registers_reg[231][2]  ( .D(n8141), .E(n1033), .CK(clk), .Q(
        \registers[231][2] ) );
  EDFFX1 \registers_reg[231][1]  ( .D(n8085), .E(n1033), .CK(clk), .Q(
        \registers[231][1] ) );
  EDFFX1 \registers_reg[231][0]  ( .D(n8027), .E(n1033), .CK(clk), .Q(
        \registers[231][0] ) );
  EDFFX1 \registers_reg[227][7]  ( .D(n8410), .E(n966), .CK(clk), .Q(
        \registers[227][7] ) );
  EDFFX1 \registers_reg[227][6]  ( .D(n8352), .E(n966), .CK(clk), .Q(
        \registers[227][6] ) );
  EDFFX1 \registers_reg[227][5]  ( .D(n8294), .E(n966), .CK(clk), .Q(
        \registers[227][5] ) );
  EDFFX1 \registers_reg[227][4]  ( .D(n8236), .E(n966), .CK(clk), .Q(
        \registers[227][4] ) );
  EDFFX1 \registers_reg[227][3]  ( .D(n8187), .E(n966), .CK(clk), .Q(
        \registers[227][3] ) );
  EDFFX1 \registers_reg[227][2]  ( .D(n8142), .E(n966), .CK(clk), .Q(
        \registers[227][2] ) );
  EDFFX1 \registers_reg[227][1]  ( .D(n8086), .E(n966), .CK(clk), .Q(
        \registers[227][1] ) );
  EDFFX1 \registers_reg[227][0]  ( .D(n8025), .E(n966), .CK(clk), .Q(
        \registers[227][0] ) );
  EDFFX1 \registers_reg[223][7]  ( .D(n8411), .E(n561), .CK(clk), .Q(
        \registers[223][7] ) );
  EDFFX1 \registers_reg[223][6]  ( .D(n8353), .E(n561), .CK(clk), .Q(
        \registers[223][6] ) );
  EDFFX1 \registers_reg[223][5]  ( .D(n8295), .E(n561), .CK(clk), .Q(
        \registers[223][5] ) );
  EDFFX1 \registers_reg[223][4]  ( .D(n8237), .E(n561), .CK(clk), .Q(
        \registers[223][4] ) );
  EDFFX1 \registers_reg[223][3]  ( .D(n8185), .E(n561), .CK(clk), .Q(
        \registers[223][3] ) );
  EDFFX1 \registers_reg[223][2]  ( .D(n8143), .E(n561), .CK(clk), .Q(
        \registers[223][2] ) );
  EDFFX1 \registers_reg[223][1]  ( .D(n8087), .E(n561), .CK(clk), .Q(
        \registers[223][1] ) );
  EDFFX1 \registers_reg[223][0]  ( .D(n8026), .E(n561), .CK(clk), .Q(
        \registers[223][0] ) );
  EDFFX1 \registers_reg[219][7]  ( .D(n8412), .E(n557), .CK(clk), .Q(
        \registers[219][7] ) );
  EDFFX1 \registers_reg[219][6]  ( .D(n8354), .E(n557), .CK(clk), .Q(
        \registers[219][6] ) );
  EDFFX1 \registers_reg[219][5]  ( .D(n8296), .E(n557), .CK(clk), .Q(
        \registers[219][5] ) );
  EDFFX1 \registers_reg[219][4]  ( .D(n8238), .E(n557), .CK(clk), .Q(
        \registers[219][4] ) );
  EDFFX1 \registers_reg[219][3]  ( .D(n8186), .E(n557), .CK(clk), .Q(
        \registers[219][3] ) );
  EDFFX1 \registers_reg[219][2]  ( .D(n8138), .E(n557), .CK(clk), .Q(
        \registers[219][2] ) );
  EDFFX1 \registers_reg[219][1]  ( .D(n8082), .E(n557), .CK(clk), .Q(
        \registers[219][1] ) );
  EDFFX1 \registers_reg[219][0]  ( .D(n8027), .E(n557), .CK(clk), .Q(
        \registers[219][0] ) );
  EDFFX1 \registers_reg[215][7]  ( .D(n8410), .E(n553), .CK(clk), .Q(
        \registers[215][7] ) );
  EDFFX1 \registers_reg[215][6]  ( .D(n8352), .E(n553), .CK(clk), .Q(
        \registers[215][6] ) );
  EDFFX1 \registers_reg[215][5]  ( .D(n8294), .E(n553), .CK(clk), .Q(
        \registers[215][5] ) );
  EDFFX1 \registers_reg[215][4]  ( .D(n8236), .E(n553), .CK(clk), .Q(
        \registers[215][4] ) );
  EDFFX1 \registers_reg[215][3]  ( .D(n8187), .E(n553), .CK(clk), .Q(
        \registers[215][3] ) );
  EDFFX1 \registers_reg[215][2]  ( .D(n8139), .E(n553), .CK(clk), .Q(
        \registers[215][2] ) );
  EDFFX1 \registers_reg[215][1]  ( .D(n8083), .E(n553), .CK(clk), .Q(
        \registers[215][1] ) );
  EDFFX1 \registers_reg[215][0]  ( .D(n8022), .E(n553), .CK(clk), .Q(
        \registers[215][0] ) );
  EDFFX1 \registers_reg[211][7]  ( .D(n8411), .E(n549), .CK(clk), .Q(
        \registers[211][7] ) );
  EDFFX1 \registers_reg[211][6]  ( .D(n8353), .E(n549), .CK(clk), .Q(
        \registers[211][6] ) );
  EDFFX1 \registers_reg[211][5]  ( .D(n8295), .E(n549), .CK(clk), .Q(
        \registers[211][5] ) );
  EDFFX1 \registers_reg[211][4]  ( .D(n8237), .E(n549), .CK(clk), .Q(
        \registers[211][4] ) );
  EDFFX1 \registers_reg[211][3]  ( .D(n8185), .E(n549), .CK(clk), .Q(
        \registers[211][3] ) );
  EDFFX1 \registers_reg[211][2]  ( .D(n8140), .E(n549), .CK(clk), .Q(
        \registers[211][2] ) );
  EDFFX1 \registers_reg[211][1]  ( .D(n8084), .E(n549), .CK(clk), .Q(
        \registers[211][1] ) );
  EDFFX1 \registers_reg[211][0]  ( .D(n8023), .E(n549), .CK(clk), .Q(
        \registers[211][0] ) );
  EDFFX1 \registers_reg[207][7]  ( .D(n8407), .E(n545), .CK(clk), .Q(
        \registers[207][7] ) );
  EDFFX1 \registers_reg[207][6]  ( .D(n8349), .E(n545), .CK(clk), .Q(
        \registers[207][6] ) );
  EDFFX1 \registers_reg[207][5]  ( .D(n8291), .E(n545), .CK(clk), .Q(
        \registers[207][5] ) );
  EDFFX1 \registers_reg[207][4]  ( .D(n8233), .E(n545), .CK(clk), .Q(
        \registers[207][4] ) );
  EDFFX1 \registers_reg[207][3]  ( .D(n8186), .E(n545), .CK(clk), .Q(
        \registers[207][3] ) );
  EDFFX1 \registers_reg[207][2]  ( .D(n8138), .E(n545), .CK(clk), .Q(
        \registers[207][2] ) );
  EDFFX1 \registers_reg[207][1]  ( .D(n8082), .E(n545), .CK(clk), .Q(
        \registers[207][1] ) );
  EDFFX1 \registers_reg[207][0]  ( .D(n8024), .E(n545), .CK(clk), .Q(
        \registers[207][0] ) );
  EDFFX1 \registers_reg[203][7]  ( .D(n8408), .E(n541), .CK(clk), .Q(
        \registers[203][7] ) );
  EDFFX1 \registers_reg[203][6]  ( .D(n8350), .E(n541), .CK(clk), .Q(
        \registers[203][6] ) );
  EDFFX1 \registers_reg[203][5]  ( .D(n8292), .E(n541), .CK(clk), .Q(
        \registers[203][5] ) );
  EDFFX1 \registers_reg[203][4]  ( .D(n8234), .E(n541), .CK(clk), .Q(
        \registers[203][4] ) );
  EDFFX1 \registers_reg[203][3]  ( .D(n8187), .E(n541), .CK(clk), .Q(
        \registers[203][3] ) );
  EDFFX1 \registers_reg[203][2]  ( .D(n8139), .E(n541), .CK(clk), .Q(
        \registers[203][2] ) );
  EDFFX1 \registers_reg[203][1]  ( .D(n8083), .E(n541), .CK(clk), .Q(
        \registers[203][1] ) );
  EDFFX1 \registers_reg[203][0]  ( .D(n8022), .E(n541), .CK(clk), .Q(
        \registers[203][0] ) );
  EDFFX1 \registers_reg[199][7]  ( .D(n8409), .E(n1029), .CK(clk), .Q(
        \registers[199][7] ) );
  EDFFX1 \registers_reg[199][6]  ( .D(n8351), .E(n1029), .CK(clk), .Q(
        \registers[199][6] ) );
  EDFFX1 \registers_reg[199][5]  ( .D(n8293), .E(n1029), .CK(clk), .Q(
        \registers[199][5] ) );
  EDFFX1 \registers_reg[199][4]  ( .D(n8235), .E(n1029), .CK(clk), .Q(
        \registers[199][4] ) );
  EDFFX1 \registers_reg[199][3]  ( .D(n8185), .E(n1029), .CK(clk), .Q(
        \registers[199][3] ) );
  EDFFX1 \registers_reg[199][2]  ( .D(n8140), .E(n1029), .CK(clk), .Q(
        \registers[199][2] ) );
  EDFFX1 \registers_reg[199][1]  ( .D(n8084), .E(n1029), .CK(clk), .Q(
        \registers[199][1] ) );
  EDFFX1 \registers_reg[199][0]  ( .D(n8023), .E(n1029), .CK(clk), .Q(
        \registers[199][0] ) );
  EDFFX1 \registers_reg[195][7]  ( .D(n8407), .E(n963), .CK(clk), .Q(
        \registers[195][7] ) );
  EDFFX1 \registers_reg[195][6]  ( .D(n8349), .E(n963), .CK(clk), .Q(
        \registers[195][6] ) );
  EDFFX1 \registers_reg[195][5]  ( .D(n8291), .E(n963), .CK(clk), .Q(
        \registers[195][5] ) );
  EDFFX1 \registers_reg[195][4]  ( .D(n8233), .E(n963), .CK(clk), .Q(
        \registers[195][4] ) );
  EDFFX1 \registers_reg[195][3]  ( .D(n8186), .E(n963), .CK(clk), .Q(
        \registers[195][3] ) );
  EDFFX1 \registers_reg[195][2]  ( .D(n8138), .E(n963), .CK(clk), .Q(
        \registers[195][2] ) );
  EDFFX1 \registers_reg[195][1]  ( .D(n8082), .E(n963), .CK(clk), .Q(
        \registers[195][1] ) );
  EDFFX1 \registers_reg[195][0]  ( .D(n8024), .E(n963), .CK(clk), .Q(
        \registers[195][0] ) );
  EDFFX1 \registers_reg[191][7]  ( .D(n8409), .E(n537), .CK(clk), .Q(
        \registers[191][7] ) );
  EDFFX1 \registers_reg[191][6]  ( .D(n8351), .E(n537), .CK(clk), .Q(
        \registers[191][6] ) );
  EDFFX1 \registers_reg[191][5]  ( .D(n8293), .E(n537), .CK(clk), .Q(
        \registers[191][5] ) );
  EDFFX1 \registers_reg[191][4]  ( .D(n8235), .E(n537), .CK(clk), .Q(
        \registers[191][4] ) );
  EDFFX1 \registers_reg[191][3]  ( .D(n8185), .E(n537), .CK(clk), .Q(
        \registers[191][3] ) );
  EDFFX1 \registers_reg[191][2]  ( .D(n8140), .E(n537), .CK(clk), .Q(
        \registers[191][2] ) );
  EDFFX1 \registers_reg[191][1]  ( .D(n8084), .E(n537), .CK(clk), .Q(
        \registers[191][1] ) );
  EDFFX1 \registers_reg[191][0]  ( .D(n8023), .E(n537), .CK(clk), .Q(
        \registers[191][0] ) );
  EDFFX1 \registers_reg[187][7]  ( .D(n8407), .E(n533), .CK(clk), .Q(
        \registers[187][7] ) );
  EDFFX1 \registers_reg[187][6]  ( .D(n8349), .E(n533), .CK(clk), .Q(
        \registers[187][6] ) );
  EDFFX1 \registers_reg[187][5]  ( .D(n8291), .E(n533), .CK(clk), .Q(
        \registers[187][5] ) );
  EDFFX1 \registers_reg[187][4]  ( .D(n8233), .E(n533), .CK(clk), .Q(
        \registers[187][4] ) );
  EDFFX1 \registers_reg[187][3]  ( .D(n8186), .E(n533), .CK(clk), .Q(
        \registers[187][3] ) );
  EDFFX1 \registers_reg[187][2]  ( .D(n8138), .E(n533), .CK(clk), .Q(
        \registers[187][2] ) );
  EDFFX1 \registers_reg[187][1]  ( .D(n8082), .E(n533), .CK(clk), .Q(
        \registers[187][1] ) );
  EDFFX1 \registers_reg[187][0]  ( .D(n8024), .E(n533), .CK(clk), .Q(
        \registers[187][0] ) );
  EDFFX1 \registers_reg[183][7]  ( .D(n8408), .E(n529), .CK(clk), .Q(
        \registers[183][7] ) );
  EDFFX1 \registers_reg[183][6]  ( .D(n8350), .E(n529), .CK(clk), .Q(
        \registers[183][6] ) );
  EDFFX1 \registers_reg[183][5]  ( .D(n8292), .E(n529), .CK(clk), .Q(
        \registers[183][5] ) );
  EDFFX1 \registers_reg[183][4]  ( .D(n8234), .E(n529), .CK(clk), .Q(
        \registers[183][4] ) );
  EDFFX1 \registers_reg[183][3]  ( .D(n8187), .E(n529), .CK(clk), .Q(
        \registers[183][3] ) );
  EDFFX1 \registers_reg[183][2]  ( .D(n8139), .E(n529), .CK(clk), .Q(
        \registers[183][2] ) );
  EDFFX1 \registers_reg[183][1]  ( .D(n8083), .E(n529), .CK(clk), .Q(
        \registers[183][1] ) );
  EDFFX1 \registers_reg[183][0]  ( .D(n8022), .E(n529), .CK(clk), .Q(
        \registers[183][0] ) );
  EDFFX1 \registers_reg[179][7]  ( .D(n8409), .E(n525), .CK(clk), .Q(
        \registers[179][7] ) );
  EDFFX1 \registers_reg[179][6]  ( .D(n8351), .E(n525), .CK(clk), .Q(
        \registers[179][6] ) );
  EDFFX1 \registers_reg[179][5]  ( .D(n8293), .E(n525), .CK(clk), .Q(
        \registers[179][5] ) );
  EDFFX1 \registers_reg[179][4]  ( .D(n8235), .E(n525), .CK(clk), .Q(
        \registers[179][4] ) );
  EDFFX1 \registers_reg[179][3]  ( .D(n8185), .E(n525), .CK(clk), .Q(
        \registers[179][3] ) );
  EDFFX1 \registers_reg[179][2]  ( .D(n8140), .E(n525), .CK(clk), .Q(
        \registers[179][2] ) );
  EDFFX1 \registers_reg[179][1]  ( .D(n8084), .E(n525), .CK(clk), .Q(
        \registers[179][1] ) );
  EDFFX1 \registers_reg[179][0]  ( .D(n8023), .E(n525), .CK(clk), .Q(
        \registers[179][0] ) );
  EDFFX1 \registers_reg[175][7]  ( .D(n8407), .E(n521), .CK(clk), .Q(
        \registers[175][7] ) );
  EDFFX1 \registers_reg[175][6]  ( .D(n8349), .E(n521), .CK(clk), .Q(
        \registers[175][6] ) );
  EDFFX1 \registers_reg[175][5]  ( .D(n8291), .E(n521), .CK(clk), .Q(
        \registers[175][5] ) );
  EDFFX1 \registers_reg[175][4]  ( .D(n8233), .E(n521), .CK(clk), .Q(
        \registers[175][4] ) );
  EDFFX1 \registers_reg[175][3]  ( .D(n8186), .E(n521), .CK(clk), .Q(
        \registers[175][3] ) );
  EDFFX1 \registers_reg[175][2]  ( .D(n8138), .E(n521), .CK(clk), .Q(
        \registers[175][2] ) );
  EDFFX1 \registers_reg[175][1]  ( .D(n8082), .E(n521), .CK(clk), .Q(
        \registers[175][1] ) );
  EDFFX1 \registers_reg[175][0]  ( .D(n8024), .E(n521), .CK(clk), .Q(
        \registers[175][0] ) );
  EDFFX1 \registers_reg[171][7]  ( .D(n8408), .E(n517), .CK(clk), .Q(
        \registers[171][7] ) );
  EDFFX1 \registers_reg[171][6]  ( .D(n8350), .E(n517), .CK(clk), .Q(
        \registers[171][6] ) );
  EDFFX1 \registers_reg[171][5]  ( .D(n8292), .E(n517), .CK(clk), .Q(
        \registers[171][5] ) );
  EDFFX1 \registers_reg[171][4]  ( .D(n8234), .E(n517), .CK(clk), .Q(
        \registers[171][4] ) );
  EDFFX1 \registers_reg[171][3]  ( .D(n8184), .E(n517), .CK(clk), .Q(
        \registers[171][3] ) );
  EDFFX1 \registers_reg[171][2]  ( .D(n8139), .E(n517), .CK(clk), .Q(
        \registers[171][2] ) );
  EDFFX1 \registers_reg[171][1]  ( .D(n8083), .E(n517), .CK(clk), .Q(
        \registers[171][1] ) );
  EDFFX1 \registers_reg[171][0]  ( .D(n8022), .E(n517), .CK(clk), .Q(
        \registers[171][0] ) );
  EDFFX1 \registers_reg[167][7]  ( .D(n8409), .E(n1025), .CK(clk), .Q(
        \registers[167][7] ) );
  EDFFX1 \registers_reg[167][6]  ( .D(n8351), .E(n1025), .CK(clk), .Q(
        \registers[167][6] ) );
  EDFFX1 \registers_reg[167][5]  ( .D(n8293), .E(n1025), .CK(clk), .Q(
        \registers[167][5] ) );
  EDFFX1 \registers_reg[167][4]  ( .D(n8235), .E(n1025), .CK(clk), .Q(
        \registers[167][4] ) );
  EDFFX1 \registers_reg[167][3]  ( .D(n8182), .E(n1025), .CK(clk), .Q(
        \registers[167][3] ) );
  EDFFX1 \registers_reg[167][2]  ( .D(n8137), .E(n1025), .CK(clk), .Q(
        \registers[167][2] ) );
  EDFFX1 \registers_reg[167][1]  ( .D(n8081), .E(n1025), .CK(clk), .Q(
        \registers[167][1] ) );
  EDFFX1 \registers_reg[167][0]  ( .D(n8020), .E(n1025), .CK(clk), .Q(
        \registers[167][0] ) );
  EDFFX1 \registers_reg[163][7]  ( .D(n8407), .E(n960), .CK(clk), .Q(
        \registers[163][7] ) );
  EDFFX1 \registers_reg[163][6]  ( .D(n8349), .E(n960), .CK(clk), .Q(
        \registers[163][6] ) );
  EDFFX1 \registers_reg[163][5]  ( .D(n8291), .E(n960), .CK(clk), .Q(
        \registers[163][5] ) );
  EDFFX1 \registers_reg[163][4]  ( .D(n8233), .E(n960), .CK(clk), .Q(
        \registers[163][4] ) );
  EDFFX1 \registers_reg[163][3]  ( .D(n8183), .E(n960), .CK(clk), .Q(
        \registers[163][3] ) );
  EDFFX1 \registers_reg[163][2]  ( .D(n8135), .E(n960), .CK(clk), .Q(
        \registers[163][2] ) );
  EDFFX1 \registers_reg[163][1]  ( .D(n8079), .E(n960), .CK(clk), .Q(
        \registers[163][1] ) );
  EDFFX1 \registers_reg[163][0]  ( .D(n8021), .E(n960), .CK(clk), .Q(
        \registers[163][0] ) );
  EDFFX1 \registers_reg[159][7]  ( .D(n8408), .E(n513), .CK(clk), .Q(
        \registers[159][7] ) );
  EDFFX1 \registers_reg[159][6]  ( .D(n8350), .E(n513), .CK(clk), .Q(
        \registers[159][6] ) );
  EDFFX1 \registers_reg[159][5]  ( .D(n8292), .E(n513), .CK(clk), .Q(
        \registers[159][5] ) );
  EDFFX1 \registers_reg[159][4]  ( .D(n8234), .E(n513), .CK(clk), .Q(
        \registers[159][4] ) );
  EDFFX1 \registers_reg[159][3]  ( .D(n8184), .E(n513), .CK(clk), .Q(
        \registers[159][3] ) );
  EDFFX1 \registers_reg[159][2]  ( .D(n8136), .E(n513), .CK(clk), .Q(
        \registers[159][2] ) );
  EDFFX1 \registers_reg[159][1]  ( .D(n8080), .E(n513), .CK(clk), .Q(
        \registers[159][1] ) );
  EDFFX1 \registers_reg[159][0]  ( .D(n8019), .E(n513), .CK(clk), .Q(
        \registers[159][0] ) );
  EDFFX1 \registers_reg[155][7]  ( .D(n8404), .E(n509), .CK(clk), .Q(
        \registers[155][7] ) );
  EDFFX1 \registers_reg[155][6]  ( .D(n8346), .E(n509), .CK(clk), .Q(
        \registers[155][6] ) );
  EDFFX1 \registers_reg[155][5]  ( .D(n8288), .E(n509), .CK(clk), .Q(
        \registers[155][5] ) );
  EDFFX1 \registers_reg[155][4]  ( .D(n8230), .E(n509), .CK(clk), .Q(
        \registers[155][4] ) );
  EDFFX1 \registers_reg[155][3]  ( .D(n8182), .E(n509), .CK(clk), .Q(
        \registers[155][3] ) );
  EDFFX1 \registers_reg[155][2]  ( .D(n8137), .E(n509), .CK(clk), .Q(
        \registers[155][2] ) );
  EDFFX1 \registers_reg[155][1]  ( .D(n8081), .E(n509), .CK(clk), .Q(
        \registers[155][1] ) );
  EDFFX1 \registers_reg[155][0]  ( .D(n8020), .E(n509), .CK(clk), .Q(
        \registers[155][0] ) );
  EDFFX1 \registers_reg[151][7]  ( .D(n8405), .E(n505), .CK(clk), .Q(
        \registers[151][7] ) );
  EDFFX1 \registers_reg[151][6]  ( .D(n8347), .E(n505), .CK(clk), .Q(
        \registers[151][6] ) );
  EDFFX1 \registers_reg[151][5]  ( .D(n8289), .E(n505), .CK(clk), .Q(
        \registers[151][5] ) );
  EDFFX1 \registers_reg[151][4]  ( .D(n8231), .E(n505), .CK(clk), .Q(
        \registers[151][4] ) );
  EDFFX1 \registers_reg[151][3]  ( .D(n8183), .E(n505), .CK(clk), .Q(
        \registers[151][3] ) );
  EDFFX1 \registers_reg[151][2]  ( .D(n8135), .E(n505), .CK(clk), .Q(
        \registers[151][2] ) );
  EDFFX1 \registers_reg[151][1]  ( .D(n8079), .E(n505), .CK(clk), .Q(
        \registers[151][1] ) );
  EDFFX1 \registers_reg[151][0]  ( .D(n8021), .E(n505), .CK(clk), .Q(
        \registers[151][0] ) );
  EDFFX1 \registers_reg[147][7]  ( .D(n8406), .E(n501), .CK(clk), .Q(
        \registers[147][7] ) );
  EDFFX1 \registers_reg[147][6]  ( .D(n8348), .E(n501), .CK(clk), .Q(
        \registers[147][6] ) );
  EDFFX1 \registers_reg[147][5]  ( .D(n8290), .E(n501), .CK(clk), .Q(
        \registers[147][5] ) );
  EDFFX1 \registers_reg[147][4]  ( .D(n8232), .E(n501), .CK(clk), .Q(
        \registers[147][4] ) );
  EDFFX1 \registers_reg[147][3]  ( .D(n8184), .E(n501), .CK(clk), .Q(
        \registers[147][3] ) );
  EDFFX1 \registers_reg[147][2]  ( .D(n8136), .E(n501), .CK(clk), .Q(
        \registers[147][2] ) );
  EDFFX1 \registers_reg[147][1]  ( .D(n8080), .E(n501), .CK(clk), .Q(
        \registers[147][1] ) );
  EDFFX1 \registers_reg[147][0]  ( .D(n8019), .E(n501), .CK(clk), .Q(
        \registers[147][0] ) );
  EDFFX1 \registers_reg[143][7]  ( .D(n8404), .E(n497), .CK(clk), .Q(
        \registers[143][7] ) );
  EDFFX1 \registers_reg[143][6]  ( .D(n8346), .E(n497), .CK(clk), .Q(
        \registers[143][6] ) );
  EDFFX1 \registers_reg[143][5]  ( .D(n8288), .E(n497), .CK(clk), .Q(
        \registers[143][5] ) );
  EDFFX1 \registers_reg[143][4]  ( .D(n8230), .E(n497), .CK(clk), .Q(
        \registers[143][4] ) );
  EDFFX1 \registers_reg[143][3]  ( .D(n8182), .E(n497), .CK(clk), .Q(
        \registers[143][3] ) );
  EDFFX1 \registers_reg[143][2]  ( .D(n8137), .E(n497), .CK(clk), .Q(
        \registers[143][2] ) );
  EDFFX1 \registers_reg[143][1]  ( .D(n8081), .E(n497), .CK(clk), .Q(
        \registers[143][1] ) );
  EDFFX1 \registers_reg[143][0]  ( .D(n8020), .E(n497), .CK(clk), .Q(
        \registers[143][0] ) );
  EDFFX1 \registers_reg[139][7]  ( .D(n8405), .E(n493), .CK(clk), .Q(
        \registers[139][7] ) );
  EDFFX1 \registers_reg[139][6]  ( .D(n8347), .E(n493), .CK(clk), .Q(
        \registers[139][6] ) );
  EDFFX1 \registers_reg[139][5]  ( .D(n8289), .E(n493), .CK(clk), .Q(
        \registers[139][5] ) );
  EDFFX1 \registers_reg[139][4]  ( .D(n8231), .E(n493), .CK(clk), .Q(
        \registers[139][4] ) );
  EDFFX1 \registers_reg[139][3]  ( .D(n8183), .E(n493), .CK(clk), .Q(
        \registers[139][3] ) );
  EDFFX1 \registers_reg[139][2]  ( .D(n8135), .E(n493), .CK(clk), .Q(
        \registers[139][2] ) );
  EDFFX1 \registers_reg[139][1]  ( .D(n8079), .E(n493), .CK(clk), .Q(
        \registers[139][1] ) );
  EDFFX1 \registers_reg[139][0]  ( .D(n8021), .E(n493), .CK(clk), .Q(
        \registers[139][0] ) );
  EDFFX1 \registers_reg[135][7]  ( .D(n8406), .E(n1021), .CK(clk), .Q(
        \registers[135][7] ) );
  EDFFX1 \registers_reg[135][6]  ( .D(n8348), .E(n1021), .CK(clk), .Q(
        \registers[135][6] ) );
  EDFFX1 \registers_reg[135][5]  ( .D(n8290), .E(n1021), .CK(clk), .Q(
        \registers[135][5] ) );
  EDFFX1 \registers_reg[135][4]  ( .D(n8232), .E(n1021), .CK(clk), .Q(
        \registers[135][4] ) );
  EDFFX1 \registers_reg[135][3]  ( .D(n8184), .E(n1021), .CK(clk), .Q(
        \registers[135][3] ) );
  EDFFX1 \registers_reg[135][2]  ( .D(n8136), .E(n1021), .CK(clk), .Q(
        \registers[135][2] ) );
  EDFFX1 \registers_reg[135][1]  ( .D(n8080), .E(n1021), .CK(clk), .Q(
        \registers[135][1] ) );
  EDFFX1 \registers_reg[135][0]  ( .D(n8019), .E(n1021), .CK(clk), .Q(
        \registers[135][0] ) );
  EDFFX1 \registers_reg[131][7]  ( .D(n8404), .E(n957), .CK(clk), .Q(
        \registers[131][7] ) );
  EDFFX1 \registers_reg[131][6]  ( .D(n8346), .E(n957), .CK(clk), .Q(
        \registers[131][6] ) );
  EDFFX1 \registers_reg[131][5]  ( .D(n8288), .E(n957), .CK(clk), .Q(
        \registers[131][5] ) );
  EDFFX1 \registers_reg[131][4]  ( .D(n8230), .E(n957), .CK(clk), .Q(
        \registers[131][4] ) );
  EDFFX1 \registers_reg[131][3]  ( .D(n8182), .E(n957), .CK(clk), .Q(
        \registers[131][3] ) );
  EDFFX1 \registers_reg[131][2]  ( .D(n8137), .E(n957), .CK(clk), .Q(
        \registers[131][2] ) );
  EDFFX1 \registers_reg[131][1]  ( .D(n8081), .E(n957), .CK(clk), .Q(
        \registers[131][1] ) );
  EDFFX1 \registers_reg[131][0]  ( .D(n8020), .E(n957), .CK(clk), .Q(
        \registers[131][0] ) );
  EDFFX1 \registers_reg[127][7]  ( .D(n8419), .E(n489), .CK(clk), .Q(
        \registers[127][7] ) );
  EDFFX1 \registers_reg[127][6]  ( .D(n8361), .E(n489), .CK(clk), .Q(
        \registers[127][6] ) );
  EDFFX1 \registers_reg[127][5]  ( .D(n8303), .E(n489), .CK(clk), .Q(
        \registers[127][5] ) );
  EDFFX1 \registers_reg[127][4]  ( .D(n8245), .E(n489), .CK(clk), .Q(
        \registers[127][4] ) );
  EDFFX1 \registers_reg[127][3]  ( .D(n8196), .E(n489), .CK(clk), .Q(
        \registers[127][3] ) );
  EDFFX1 \registers_reg[127][2]  ( .D(n8151), .E(n489), .CK(clk), .Q(
        \registers[127][2] ) );
  EDFFX1 \registers_reg[127][1]  ( .D(n8095), .E(n489), .CK(clk), .Q(
        \registers[127][1] ) );
  EDFFX1 \registers_reg[127][0]  ( .D(n8034), .E(n489), .CK(clk), .Q(
        \registers[127][0] ) );
  EDFFX1 \registers_reg[123][7]  ( .D(n8420), .E(n485), .CK(clk), .Q(
        \registers[123][7] ) );
  EDFFX1 \registers_reg[123][6]  ( .D(n8362), .E(n485), .CK(clk), .Q(
        \registers[123][6] ) );
  EDFFX1 \registers_reg[123][5]  ( .D(n8304), .E(n485), .CK(clk), .Q(
        \registers[123][5] ) );
  EDFFX1 \registers_reg[123][4]  ( .D(n8246), .E(n485), .CK(clk), .Q(
        \registers[123][4] ) );
  EDFFX1 \registers_reg[123][3]  ( .D(n8194), .E(n485), .CK(clk), .Q(
        \registers[123][3] ) );
  EDFFX1 \registers_reg[123][2]  ( .D(n8727), .E(n485), .CK(clk), .Q(
        \registers[123][2] ) );
  EDFFX1 \registers_reg[123][1]  ( .D(n8699), .E(n485), .CK(clk), .Q(
        \registers[123][1] ) );
  EDFFX1 \registers_reg[123][0]  ( .D(n8036), .E(n485), .CK(clk), .Q(
        \registers[123][0] ) );
  EDFFX1 \registers_reg[119][7]  ( .D(n8421), .E(n481), .CK(clk), .Q(
        \registers[119][7] ) );
  EDFFX1 \registers_reg[119][6]  ( .D(n8363), .E(n481), .CK(clk), .Q(
        \registers[119][6] ) );
  EDFFX1 \registers_reg[119][5]  ( .D(n8305), .E(n481), .CK(clk), .Q(
        \registers[119][5] ) );
  EDFFX1 \registers_reg[119][4]  ( .D(n8247), .E(n481), .CK(clk), .Q(
        \registers[119][4] ) );
  EDFFX1 \registers_reg[119][3]  ( .D(n8195), .E(n481), .CK(clk), .Q(
        \registers[119][3] ) );
  EDFFX1 \registers_reg[119][2]  ( .D(n8150), .E(n481), .CK(clk), .Q(
        \registers[119][2] ) );
  EDFFX1 \registers_reg[119][1]  ( .D(n8094), .E(n481), .CK(clk), .Q(
        \registers[119][1] ) );
  EDFFX1 \registers_reg[119][0]  ( .D(n8034), .E(n481), .CK(clk), .Q(
        \registers[119][0] ) );
  EDFFX1 \registers_reg[115][7]  ( .D(n8419), .E(n477), .CK(clk), .Q(
        \registers[115][7] ) );
  EDFFX1 \registers_reg[115][6]  ( .D(n8361), .E(n477), .CK(clk), .Q(
        \registers[115][6] ) );
  EDFFX1 \registers_reg[115][5]  ( .D(n8303), .E(n477), .CK(clk), .Q(
        \registers[115][5] ) );
  EDFFX1 \registers_reg[115][4]  ( .D(n8245), .E(n477), .CK(clk), .Q(
        \registers[115][4] ) );
  EDFFX1 \registers_reg[115][3]  ( .D(n8196), .E(n477), .CK(clk), .Q(
        \registers[115][3] ) );
  EDFFX1 \registers_reg[115][2]  ( .D(n8148), .E(n477), .CK(clk), .Q(
        \registers[115][2] ) );
  EDFFX1 \registers_reg[115][1]  ( .D(n8092), .E(n477), .CK(clk), .Q(
        \registers[115][1] ) );
  EDFFX1 \registers_reg[115][0]  ( .D(n8032), .E(n477), .CK(clk), .Q(
        \registers[115][0] ) );
  EDFFX1 \registers_reg[111][7]  ( .D(n8420), .E(n473), .CK(clk), .Q(
        \registers[111][7] ) );
  EDFFX1 \registers_reg[111][6]  ( .D(n8362), .E(n473), .CK(clk), .Q(
        \registers[111][6] ) );
  EDFFX1 \registers_reg[111][5]  ( .D(n8304), .E(n473), .CK(clk), .Q(
        \registers[111][5] ) );
  EDFFX1 \registers_reg[111][4]  ( .D(n8246), .E(n473), .CK(clk), .Q(
        \registers[111][4] ) );
  EDFFX1 \registers_reg[111][3]  ( .D(n8194), .E(n473), .CK(clk), .Q(
        \registers[111][3] ) );
  EDFFX1 \registers_reg[111][2]  ( .D(n8149), .E(n473), .CK(clk), .Q(
        \registers[111][2] ) );
  EDFFX1 \registers_reg[111][1]  ( .D(n8093), .E(n473), .CK(clk), .Q(
        \registers[111][1] ) );
  EDFFX1 \registers_reg[111][0]  ( .D(n8033), .E(n473), .CK(clk), .Q(
        \registers[111][0] ) );
  EDFFX1 \registers_reg[107][7]  ( .D(n8421), .E(n469), .CK(clk), .Q(
        \registers[107][7] ) );
  EDFFX1 \registers_reg[107][6]  ( .D(n8363), .E(n469), .CK(clk), .Q(
        \registers[107][6] ) );
  EDFFX1 \registers_reg[107][5]  ( .D(n8305), .E(n469), .CK(clk), .Q(
        \registers[107][5] ) );
  EDFFX1 \registers_reg[107][4]  ( .D(n8247), .E(n469), .CK(clk), .Q(
        \registers[107][4] ) );
  EDFFX1 \registers_reg[107][3]  ( .D(n8195), .E(n469), .CK(clk), .Q(
        \registers[107][3] ) );
  EDFFX1 \registers_reg[107][2]  ( .D(n8147), .E(n469), .CK(clk), .Q(
        \registers[107][2] ) );
  EDFFX1 \registers_reg[107][1]  ( .D(n8091), .E(n469), .CK(clk), .Q(
        \registers[107][1] ) );
  EDFFX1 \registers_reg[107][0]  ( .D(n8031), .E(n469), .CK(clk), .Q(
        \registers[107][0] ) );
  EDFFX1 \registers_reg[103][7]  ( .D(n8419), .E(n954), .CK(clk), .Q(
        \registers[103][7] ) );
  EDFFX1 \registers_reg[103][6]  ( .D(n8361), .E(n954), .CK(clk), .Q(
        \registers[103][6] ) );
  EDFFX1 \registers_reg[103][5]  ( .D(n8303), .E(n954), .CK(clk), .Q(
        \registers[103][5] ) );
  EDFFX1 \registers_reg[103][4]  ( .D(n8245), .E(n954), .CK(clk), .Q(
        \registers[103][4] ) );
  EDFFX1 \registers_reg[103][3]  ( .D(n8193), .E(n954), .CK(clk), .Q(
        \registers[103][3] ) );
  EDFFX1 \registers_reg[103][2]  ( .D(n8148), .E(n954), .CK(clk), .Q(
        \registers[103][2] ) );
  EDFFX1 \registers_reg[103][1]  ( .D(n8092), .E(n954), .CK(clk), .Q(
        \registers[103][1] ) );
  EDFFX1 \registers_reg[103][0]  ( .D(n8032), .E(n954), .CK(clk), .Q(
        \registers[103][0] ) );
  EDFFX1 \registers_reg[99][7]  ( .D(n8418), .E(n950), .CK(clk), .Q(
        \registers[99][7] ) );
  EDFFX1 \registers_reg[99][6]  ( .D(n8360), .E(n950), .CK(clk), .Q(
        \registers[99][6] ) );
  EDFFX1 \registers_reg[99][5]  ( .D(n8302), .E(n950), .CK(clk), .Q(
        \registers[99][5] ) );
  EDFFX1 \registers_reg[99][4]  ( .D(n8244), .E(n950), .CK(clk), .Q(
        \registers[99][4] ) );
  EDFFX1 \registers_reg[99][3]  ( .D(n8191), .E(n950), .CK(clk), .Q(
        \registers[99][3] ) );
  EDFFX1 \registers_reg[99][2]  ( .D(n8149), .E(n950), .CK(clk), .Q(
        \registers[99][2] ) );
  EDFFX1 \registers_reg[99][1]  ( .D(n8093), .E(n950), .CK(clk), .Q(
        \registers[99][1] ) );
  EDFFX1 \registers_reg[99][0]  ( .D(n8033), .E(n950), .CK(clk), .Q(
        \registers[99][0] ) );
  EDFFX1 \registers_reg[95][7]  ( .D(n8416), .E(n465), .CK(clk), .Q(
        \registers[95][7] ) );
  EDFFX1 \registers_reg[95][6]  ( .D(n8358), .E(n465), .CK(clk), .Q(
        \registers[95][6] ) );
  EDFFX1 \registers_reg[95][5]  ( .D(n8300), .E(n465), .CK(clk), .Q(
        \registers[95][5] ) );
  EDFFX1 \registers_reg[95][4]  ( .D(n8242), .E(n465), .CK(clk), .Q(
        \registers[95][4] ) );
  EDFFX1 \registers_reg[95][3]  ( .D(n8192), .E(n465), .CK(clk), .Q(
        \registers[95][3] ) );
  EDFFX1 \registers_reg[95][2]  ( .D(n8147), .E(n465), .CK(clk), .Q(
        \registers[95][2] ) );
  EDFFX1 \registers_reg[95][1]  ( .D(n8091), .E(n465), .CK(clk), .Q(
        \registers[95][1] ) );
  EDFFX1 \registers_reg[95][0]  ( .D(n8031), .E(n465), .CK(clk), .Q(
        \registers[95][0] ) );
  EDFFX1 \registers_reg[91][7]  ( .D(n8417), .E(n461), .CK(clk), .Q(
        \registers[91][7] ) );
  EDFFX1 \registers_reg[91][6]  ( .D(n8359), .E(n461), .CK(clk), .Q(
        \registers[91][6] ) );
  EDFFX1 \registers_reg[91][5]  ( .D(n8301), .E(n461), .CK(clk), .Q(
        \registers[91][5] ) );
  EDFFX1 \registers_reg[91][4]  ( .D(n8243), .E(n461), .CK(clk), .Q(
        \registers[91][4] ) );
  EDFFX1 \registers_reg[91][3]  ( .D(n8193), .E(n461), .CK(clk), .Q(
        \registers[91][3] ) );
  EDFFX1 \registers_reg[91][2]  ( .D(n8148), .E(n461), .CK(clk), .Q(
        \registers[91][2] ) );
  EDFFX1 \registers_reg[91][1]  ( .D(n8092), .E(n461), .CK(clk), .Q(
        \registers[91][1] ) );
  EDFFX1 \registers_reg[91][0]  ( .D(n8032), .E(n461), .CK(clk), .Q(
        \registers[91][0] ) );
  EDFFX1 \registers_reg[87][7]  ( .D(n8418), .E(n457), .CK(clk), .Q(
        \registers[87][7] ) );
  EDFFX1 \registers_reg[87][6]  ( .D(n8360), .E(n457), .CK(clk), .Q(
        \registers[87][6] ) );
  EDFFX1 \registers_reg[87][5]  ( .D(n8302), .E(n457), .CK(clk), .Q(
        \registers[87][5] ) );
  EDFFX1 \registers_reg[87][4]  ( .D(n8244), .E(n457), .CK(clk), .Q(
        \registers[87][4] ) );
  EDFFX1 \registers_reg[87][3]  ( .D(n8191), .E(n457), .CK(clk), .Q(
        \registers[87][3] ) );
  EDFFX1 \registers_reg[87][2]  ( .D(n8149), .E(n457), .CK(clk), .Q(
        \registers[87][2] ) );
  EDFFX1 \registers_reg[87][1]  ( .D(n8093), .E(n457), .CK(clk), .Q(
        \registers[87][1] ) );
  EDFFX1 \registers_reg[87][0]  ( .D(n8033), .E(n457), .CK(clk), .Q(
        \registers[87][0] ) );
  EDFFX1 \registers_reg[83][7]  ( .D(n8416), .E(n453), .CK(clk), .Q(
        \registers[83][7] ) );
  EDFFX1 \registers_reg[83][6]  ( .D(n8358), .E(n453), .CK(clk), .Q(
        \registers[83][6] ) );
  EDFFX1 \registers_reg[83][5]  ( .D(n8300), .E(n453), .CK(clk), .Q(
        \registers[83][5] ) );
  EDFFX1 \registers_reg[83][4]  ( .D(n8242), .E(n453), .CK(clk), .Q(
        \registers[83][4] ) );
  EDFFX1 \registers_reg[83][3]  ( .D(n8192), .E(n453), .CK(clk), .Q(
        \registers[83][3] ) );
  EDFFX1 \registers_reg[83][2]  ( .D(n8147), .E(n453), .CK(clk), .Q(
        \registers[83][2] ) );
  EDFFX1 \registers_reg[83][1]  ( .D(n8091), .E(n453), .CK(clk), .Q(
        \registers[83][1] ) );
  EDFFX1 \registers_reg[83][0]  ( .D(n8031), .E(n453), .CK(clk), .Q(
        \registers[83][0] ) );
  EDFFX1 \registers_reg[79][7]  ( .D(n8417), .E(n449), .CK(clk), .Q(
        \registers[79][7] ) );
  EDFFX1 \registers_reg[79][6]  ( .D(n8359), .E(n449), .CK(clk), .Q(
        \registers[79][6] ) );
  EDFFX1 \registers_reg[79][5]  ( .D(n8301), .E(n449), .CK(clk), .Q(
        \registers[79][5] ) );
  EDFFX1 \registers_reg[79][4]  ( .D(n8243), .E(n449), .CK(clk), .Q(
        \registers[79][4] ) );
  EDFFX1 \registers_reg[79][3]  ( .D(n8193), .E(n449), .CK(clk), .Q(
        \registers[79][3] ) );
  EDFFX1 \registers_reg[79][2]  ( .D(n8148), .E(n449), .CK(clk), .Q(
        \registers[79][2] ) );
  EDFFX1 \registers_reg[79][1]  ( .D(n8092), .E(n449), .CK(clk), .Q(
        \registers[79][1] ) );
  EDFFX1 \registers_reg[79][0]  ( .D(n8032), .E(n449), .CK(clk), .Q(
        \registers[79][0] ) );
  EDFFX1 \registers_reg[75][7]  ( .D(n8418), .E(n445), .CK(clk), .Q(
        \registers[75][7] ) );
  EDFFX1 \registers_reg[75][6]  ( .D(n8360), .E(n445), .CK(clk), .Q(
        \registers[75][6] ) );
  EDFFX1 \registers_reg[75][5]  ( .D(n8302), .E(n445), .CK(clk), .Q(
        \registers[75][5] ) );
  EDFFX1 \registers_reg[75][4]  ( .D(n8244), .E(n445), .CK(clk), .Q(
        \registers[75][4] ) );
  EDFFX1 \registers_reg[75][3]  ( .D(n8191), .E(n445), .CK(clk), .Q(
        \registers[75][3] ) );
  EDFFX1 \registers_reg[75][2]  ( .D(n8149), .E(n445), .CK(clk), .Q(
        \registers[75][2] ) );
  EDFFX1 \registers_reg[75][1]  ( .D(n8093), .E(n445), .CK(clk), .Q(
        \registers[75][1] ) );
  EDFFX1 \registers_reg[75][0]  ( .D(n8033), .E(n445), .CK(clk), .Q(
        \registers[75][0] ) );
  EDFFX1 \registers_reg[71][7]  ( .D(n8416), .E(n947), .CK(clk), .Q(
        \registers[71][7] ) );
  EDFFX1 \registers_reg[71][6]  ( .D(n8358), .E(n947), .CK(clk), .Q(
        \registers[71][6] ) );
  EDFFX1 \registers_reg[71][5]  ( .D(n8300), .E(n947), .CK(clk), .Q(
        \registers[71][5] ) );
  EDFFX1 \registers_reg[71][4]  ( .D(n8242), .E(n947), .CK(clk), .Q(
        \registers[71][4] ) );
  EDFFX1 \registers_reg[71][3]  ( .D(n8192), .E(n947), .CK(clk), .Q(
        \registers[71][3] ) );
  EDFFX1 \registers_reg[71][2]  ( .D(n8147), .E(n947), .CK(clk), .Q(
        \registers[71][2] ) );
  EDFFX1 \registers_reg[71][1]  ( .D(n8091), .E(n947), .CK(clk), .Q(
        \registers[71][1] ) );
  EDFFX1 \registers_reg[71][0]  ( .D(n8031), .E(n947), .CK(clk), .Q(
        \registers[71][0] ) );
  EDFFX1 \registers_reg[67][7]  ( .D(n8417), .E(n943), .CK(clk), .Q(
        \registers[67][7] ) );
  EDFFX1 \registers_reg[67][6]  ( .D(n8359), .E(n943), .CK(clk), .Q(
        \registers[67][6] ) );
  EDFFX1 \registers_reg[67][5]  ( .D(n8301), .E(n943), .CK(clk), .Q(
        \registers[67][5] ) );
  EDFFX1 \registers_reg[67][4]  ( .D(n8243), .E(n943), .CK(clk), .Q(
        \registers[67][4] ) );
  EDFFX1 \registers_reg[67][3]  ( .D(n8193), .E(n943), .CK(clk), .Q(
        \registers[67][3] ) );
  EDFFX1 \registers_reg[67][2]  ( .D(n8148), .E(n943), .CK(clk), .Q(
        \registers[67][2] ) );
  EDFFX1 \registers_reg[67][1]  ( .D(n8092), .E(n943), .CK(clk), .Q(
        \registers[67][1] ) );
  EDFFX1 \registers_reg[67][0]  ( .D(n8032), .E(n943), .CK(clk), .Q(
        \registers[67][0] ) );
  EDFFX1 \registers_reg[63][7]  ( .D(n8416), .E(n441), .CK(clk), .Q(
        \registers[63][7] ) );
  EDFFX1 \registers_reg[63][6]  ( .D(n8358), .E(n441), .CK(clk), .Q(
        \registers[63][6] ) );
  EDFFX1 \registers_reg[63][5]  ( .D(n8300), .E(n441), .CK(clk), .Q(
        \registers[63][5] ) );
  EDFFX1 \registers_reg[63][4]  ( .D(n8242), .E(n441), .CK(clk), .Q(
        \registers[63][4] ) );
  EDFFX1 \registers_reg[63][3]  ( .D(n8192), .E(n441), .CK(clk), .Q(
        \registers[63][3] ) );
  EDFFX1 \registers_reg[63][2]  ( .D(n8144), .E(n441), .CK(clk), .Q(
        \registers[63][2] ) );
  EDFFX1 \registers_reg[63][1]  ( .D(n8088), .E(n441), .CK(clk), .Q(
        \registers[63][1] ) );
  EDFFX1 \registers_reg[63][0]  ( .D(n8028), .E(n441), .CK(clk), .Q(
        \registers[63][0] ) );
  EDFFX1 \registers_reg[59][7]  ( .D(n8417), .E(n437), .CK(clk), .Q(
        \registers[59][7] ) );
  EDFFX1 \registers_reg[59][6]  ( .D(n8359), .E(n437), .CK(clk), .Q(
        \registers[59][6] ) );
  EDFFX1 \registers_reg[59][5]  ( .D(n8301), .E(n437), .CK(clk), .Q(
        \registers[59][5] ) );
  EDFFX1 \registers_reg[59][4]  ( .D(n8243), .E(n437), .CK(clk), .Q(
        \registers[59][4] ) );
  EDFFX1 \registers_reg[59][3]  ( .D(n8193), .E(n437), .CK(clk), .Q(
        \registers[59][3] ) );
  EDFFX1 \registers_reg[59][2]  ( .D(n8145), .E(n437), .CK(clk), .Q(
        \registers[59][2] ) );
  EDFFX1 \registers_reg[59][1]  ( .D(n8089), .E(n437), .CK(clk), .Q(
        \registers[59][1] ) );
  EDFFX1 \registers_reg[59][0]  ( .D(n8029), .E(n437), .CK(clk), .Q(
        \registers[59][0] ) );
  EDFFX1 \registers_reg[55][7]  ( .D(n8418), .E(n433), .CK(clk), .Q(
        \registers[55][7] ) );
  EDFFX1 \registers_reg[55][6]  ( .D(n8360), .E(n433), .CK(clk), .Q(
        \registers[55][6] ) );
  EDFFX1 \registers_reg[55][5]  ( .D(n8302), .E(n433), .CK(clk), .Q(
        \registers[55][5] ) );
  EDFFX1 \registers_reg[55][4]  ( .D(n8244), .E(n433), .CK(clk), .Q(
        \registers[55][4] ) );
  EDFFX1 \registers_reg[55][3]  ( .D(n8191), .E(n433), .CK(clk), .Q(
        \registers[55][3] ) );
  EDFFX1 \registers_reg[55][2]  ( .D(n8146), .E(n433), .CK(clk), .Q(
        \registers[55][2] ) );
  EDFFX1 \registers_reg[55][1]  ( .D(n8090), .E(n433), .CK(clk), .Q(
        \registers[55][1] ) );
  EDFFX1 \registers_reg[55][0]  ( .D(n8030), .E(n433), .CK(clk), .Q(
        \registers[55][0] ) );
  EDFFX1 \registers_reg[51][7]  ( .D(n8414), .E(n429), .CK(clk), .Q(
        \registers[51][7] ) );
  EDFFX1 \registers_reg[51][6]  ( .D(n8356), .E(n429), .CK(clk), .Q(
        \registers[51][6] ) );
  EDFFX1 \registers_reg[51][5]  ( .D(n8298), .E(n429), .CK(clk), .Q(
        \registers[51][5] ) );
  EDFFX1 \registers_reg[51][4]  ( .D(n8240), .E(n429), .CK(clk), .Q(
        \registers[51][4] ) );
  EDFFX1 \registers_reg[51][3]  ( .D(n8192), .E(n429), .CK(clk), .Q(
        \registers[51][3] ) );
  EDFFX1 \registers_reg[51][2]  ( .D(n8144), .E(n429), .CK(clk), .Q(
        \registers[51][2] ) );
  EDFFX1 \registers_reg[51][1]  ( .D(n8088), .E(n429), .CK(clk), .Q(
        \registers[51][1] ) );
  EDFFX1 \registers_reg[51][0]  ( .D(n8028), .E(n429), .CK(clk), .Q(
        \registers[51][0] ) );
  EDFFX1 \registers_reg[47][7]  ( .D(n8415), .E(n425), .CK(clk), .Q(
        \registers[47][7] ) );
  EDFFX1 \registers_reg[47][6]  ( .D(n8357), .E(n425), .CK(clk), .Q(
        \registers[47][6] ) );
  EDFFX1 \registers_reg[47][5]  ( .D(n8299), .E(n425), .CK(clk), .Q(
        \registers[47][5] ) );
  EDFFX1 \registers_reg[47][4]  ( .D(n8241), .E(n425), .CK(clk), .Q(
        \registers[47][4] ) );
  EDFFX1 \registers_reg[47][3]  ( .D(n8193), .E(n425), .CK(clk), .Q(
        \registers[47][3] ) );
  EDFFX1 \registers_reg[47][2]  ( .D(n8145), .E(n425), .CK(clk), .Q(
        \registers[47][2] ) );
  EDFFX1 \registers_reg[47][1]  ( .D(n8089), .E(n425), .CK(clk), .Q(
        \registers[47][1] ) );
  EDFFX1 \registers_reg[47][0]  ( .D(n8029), .E(n425), .CK(clk), .Q(
        \registers[47][0] ) );
  EDFFX1 \registers_reg[43][7]  ( .D(n8413), .E(n421), .CK(clk), .Q(
        \registers[43][7] ) );
  EDFFX1 \registers_reg[43][6]  ( .D(n8355), .E(n421), .CK(clk), .Q(
        \registers[43][6] ) );
  EDFFX1 \registers_reg[43][5]  ( .D(n8297), .E(n421), .CK(clk), .Q(
        \registers[43][5] ) );
  EDFFX1 \registers_reg[43][4]  ( .D(n8239), .E(n421), .CK(clk), .Q(
        \registers[43][4] ) );
  EDFFX1 \registers_reg[43][3]  ( .D(n8188), .E(n421), .CK(clk), .Q(
        \registers[43][3] ) );
  EDFFX1 \registers_reg[43][2]  ( .D(n8146), .E(n421), .CK(clk), .Q(
        \registers[43][2] ) );
  EDFFX1 \registers_reg[43][1]  ( .D(n8090), .E(n421), .CK(clk), .Q(
        \registers[43][1] ) );
  EDFFX1 \registers_reg[43][0]  ( .D(n8030), .E(n421), .CK(clk), .Q(
        \registers[43][0] ) );
  EDFFX1 \registers_reg[39][7]  ( .D(n8414), .E(n940), .CK(clk), .Q(
        \registers[39][7] ) );
  EDFFX1 \registers_reg[39][6]  ( .D(n8356), .E(n940), .CK(clk), .Q(
        \registers[39][6] ) );
  EDFFX1 \registers_reg[39][5]  ( .D(n8298), .E(n940), .CK(clk), .Q(
        \registers[39][5] ) );
  EDFFX1 \registers_reg[39][4]  ( .D(n8240), .E(n940), .CK(clk), .Q(
        \registers[39][4] ) );
  EDFFX1 \registers_reg[39][3]  ( .D(n8189), .E(n940), .CK(clk), .Q(
        \registers[39][3] ) );
  EDFFX1 \registers_reg[39][2]  ( .D(n8144), .E(n940), .CK(clk), .Q(
        \registers[39][2] ) );
  EDFFX1 \registers_reg[39][1]  ( .D(n8088), .E(n940), .CK(clk), .Q(
        \registers[39][1] ) );
  EDFFX1 \registers_reg[39][0]  ( .D(n8028), .E(n940), .CK(clk), .Q(
        \registers[39][0] ) );
  EDFFX1 \registers_reg[35][7]  ( .D(n8415), .E(n936), .CK(clk), .Q(
        \registers[35][7] ) );
  EDFFX1 \registers_reg[35][6]  ( .D(n8357), .E(n936), .CK(clk), .Q(
        \registers[35][6] ) );
  EDFFX1 \registers_reg[35][5]  ( .D(n8299), .E(n936), .CK(clk), .Q(
        \registers[35][5] ) );
  EDFFX1 \registers_reg[35][4]  ( .D(n8241), .E(n936), .CK(clk), .Q(
        \registers[35][4] ) );
  EDFFX1 \registers_reg[35][3]  ( .D(n8190), .E(n936), .CK(clk), .Q(
        \registers[35][3] ) );
  EDFFX1 \registers_reg[35][2]  ( .D(n8145), .E(n936), .CK(clk), .Q(
        \registers[35][2] ) );
  EDFFX1 \registers_reg[35][1]  ( .D(n8089), .E(n936), .CK(clk), .Q(
        \registers[35][1] ) );
  EDFFX1 \registers_reg[35][0]  ( .D(n8029), .E(n936), .CK(clk), .Q(
        \registers[35][0] ) );
  EDFFX1 \registers_reg[31][7]  ( .D(n8413), .E(n417), .CK(clk), .Q(
        \registers[31][7] ) );
  EDFFX1 \registers_reg[31][6]  ( .D(n8355), .E(n417), .CK(clk), .Q(
        \registers[31][6] ) );
  EDFFX1 \registers_reg[31][5]  ( .D(n8297), .E(n417), .CK(clk), .Q(
        \registers[31][5] ) );
  EDFFX1 \registers_reg[31][4]  ( .D(n8239), .E(n417), .CK(clk), .Q(
        \registers[31][4] ) );
  EDFFX1 \registers_reg[31][3]  ( .D(n8188), .E(n417), .CK(clk), .Q(
        \registers[31][3] ) );
  EDFFX1 \registers_reg[31][2]  ( .D(n8146), .E(n417), .CK(clk), .Q(
        \registers[31][2] ) );
  EDFFX1 \registers_reg[31][1]  ( .D(n8090), .E(n417), .CK(clk), .Q(
        \registers[31][1] ) );
  EDFFX1 \registers_reg[31][0]  ( .D(n8030), .E(n417), .CK(clk), .Q(
        \registers[31][0] ) );
  EDFFX1 \registers_reg[27][7]  ( .D(n8414), .E(n413), .CK(clk), .Q(
        \registers[27][7] ) );
  EDFFX1 \registers_reg[27][6]  ( .D(n8356), .E(n413), .CK(clk), .Q(
        \registers[27][6] ) );
  EDFFX1 \registers_reg[27][5]  ( .D(n8298), .E(n413), .CK(clk), .Q(
        \registers[27][5] ) );
  EDFFX1 \registers_reg[27][4]  ( .D(n8240), .E(n413), .CK(clk), .Q(
        \registers[27][4] ) );
  EDFFX1 \registers_reg[27][3]  ( .D(n8189), .E(n413), .CK(clk), .Q(
        \registers[27][3] ) );
  EDFFX1 \registers_reg[27][2]  ( .D(n8144), .E(n413), .CK(clk), .Q(
        \registers[27][2] ) );
  EDFFX1 \registers_reg[27][1]  ( .D(n8088), .E(n413), .CK(clk), .Q(
        \registers[27][1] ) );
  EDFFX1 \registers_reg[27][0]  ( .D(n8028), .E(n413), .CK(clk), .Q(
        \registers[27][0] ) );
  EDFFX1 \registers_reg[23][7]  ( .D(n8415), .E(n409), .CK(clk), .Q(
        \registers[23][7] ) );
  EDFFX1 \registers_reg[23][6]  ( .D(n8357), .E(n409), .CK(clk), .Q(
        \registers[23][6] ) );
  EDFFX1 \registers_reg[23][5]  ( .D(n8299), .E(n409), .CK(clk), .Q(
        \registers[23][5] ) );
  EDFFX1 \registers_reg[23][4]  ( .D(n8241), .E(n409), .CK(clk), .Q(
        \registers[23][4] ) );
  EDFFX1 \registers_reg[23][3]  ( .D(n8190), .E(n409), .CK(clk), .Q(
        \registers[23][3] ) );
  EDFFX1 \registers_reg[23][2]  ( .D(n8145), .E(n409), .CK(clk), .Q(
        \registers[23][2] ) );
  EDFFX1 \registers_reg[23][1]  ( .D(n8089), .E(n409), .CK(clk), .Q(
        \registers[23][1] ) );
  EDFFX1 \registers_reg[23][0]  ( .D(n8029), .E(n409), .CK(clk), .Q(
        \registers[23][0] ) );
  EDFFX1 \registers_reg[19][7]  ( .D(n8413), .E(n405), .CK(clk), .Q(
        \registers[19][7] ) );
  EDFFX1 \registers_reg[19][6]  ( .D(n8355), .E(n405), .CK(clk), .Q(
        \registers[19][6] ) );
  EDFFX1 \registers_reg[19][5]  ( .D(n8297), .E(n405), .CK(clk), .Q(
        \registers[19][5] ) );
  EDFFX1 \registers_reg[19][4]  ( .D(n8239), .E(n405), .CK(clk), .Q(
        \registers[19][4] ) );
  EDFFX1 \registers_reg[19][3]  ( .D(n8188), .E(n405), .CK(clk), .Q(
        \registers[19][3] ) );
  EDFFX1 \registers_reg[19][2]  ( .D(n8146), .E(n405), .CK(clk), .Q(
        \registers[19][2] ) );
  EDFFX1 \registers_reg[19][1]  ( .D(n8090), .E(n405), .CK(clk), .Q(
        \registers[19][1] ) );
  EDFFX1 \registers_reg[19][0]  ( .D(n8030), .E(n405), .CK(clk), .Q(
        \registers[19][0] ) );
  EDFFX1 \registers_reg[15][7]  ( .D(n8414), .E(n401), .CK(clk), .Q(
        \registers[15][7] ) );
  EDFFX1 \registers_reg[15][6]  ( .D(n8356), .E(n401), .CK(clk), .Q(
        \registers[15][6] ) );
  EDFFX1 \registers_reg[15][5]  ( .D(n8298), .E(n401), .CK(clk), .Q(
        \registers[15][5] ) );
  EDFFX1 \registers_reg[15][4]  ( .D(n8240), .E(n401), .CK(clk), .Q(
        \registers[15][4] ) );
  EDFFX1 \registers_reg[15][3]  ( .D(n8189), .E(n401), .CK(clk), .Q(
        \registers[15][3] ) );
  EDFFX1 \registers_reg[15][2]  ( .D(n8141), .E(n401), .CK(clk), .Q(
        \registers[15][2] ) );
  EDFFX1 \registers_reg[15][1]  ( .D(n8085), .E(n401), .CK(clk), .Q(
        \registers[15][1] ) );
  EDFFX1 \registers_reg[15][0]  ( .D(n8025), .E(n401), .CK(clk), .Q(
        \registers[15][0] ) );
  EDFFX1 \registers_reg[11][7]  ( .D(n8415), .E(n397), .CK(clk), .Q(
        \registers[11][7] ) );
  EDFFX1 \registers_reg[11][6]  ( .D(n8357), .E(n397), .CK(clk), .Q(
        \registers[11][6] ) );
  EDFFX1 \registers_reg[11][5]  ( .D(n8299), .E(n397), .CK(clk), .Q(
        \registers[11][5] ) );
  EDFFX1 \registers_reg[11][4]  ( .D(n8241), .E(n397), .CK(clk), .Q(
        \registers[11][4] ) );
  EDFFX1 \registers_reg[11][3]  ( .D(n8190), .E(n397), .CK(clk), .Q(
        \registers[11][3] ) );
  EDFFX1 \registers_reg[11][2]  ( .D(n8142), .E(n397), .CK(clk), .Q(
        \registers[11][2] ) );
  EDFFX1 \registers_reg[11][1]  ( .D(n8086), .E(n397), .CK(clk), .Q(
        \registers[11][1] ) );
  EDFFX1 \registers_reg[11][0]  ( .D(n8026), .E(n397), .CK(clk), .Q(
        \registers[11][0] ) );
  EDFFX1 \registers_reg[7][7]  ( .D(n8413), .E(n1017), .CK(clk), .Q(
        \registers[7][7] ) );
  EDFFX1 \registers_reg[7][6]  ( .D(n8355), .E(n1017), .CK(clk), .Q(
        \registers[7][6] ), .QN(n1120) );
  EDFFX1 \registers_reg[7][5]  ( .D(n8297), .E(n1017), .CK(clk), .Q(
        \registers[7][5] ), .QN(n1121) );
  EDFFX1 \registers_reg[7][4]  ( .D(n8239), .E(n1017), .CK(clk), .Q(
        \registers[7][4] ), .QN(n1122) );
  EDFFX1 \registers_reg[7][3]  ( .D(n8188), .E(n1017), .CK(clk), .Q(
        \registers[7][3] ), .QN(n1123) );
  EDFFX1 \registers_reg[7][2]  ( .D(n8143), .E(n1017), .CK(clk), .Q(
        \registers[7][2] ), .QN(n1124) );
  EDFFX1 \registers_reg[7][1]  ( .D(n8087), .E(n1017), .CK(clk), .Q(
        \registers[7][1] ), .QN(n1125) );
  EDFFX1 \registers_reg[7][0]  ( .D(n8027), .E(n1017), .CK(clk), .Q(
        \registers[7][0] ), .QN(n1126) );
  EDFFX1 \registers_reg[3][7]  ( .D(n8414), .E(n393), .CK(clk), .Q(
        \registers[3][7] ) );
  EDFFX1 \registers_reg[3][6]  ( .D(n8356), .E(n393), .CK(clk), .Q(
        \registers[3][6] ) );
  EDFFX1 \registers_reg[3][5]  ( .D(n8298), .E(n393), .CK(clk), .Q(
        \registers[3][5] ) );
  EDFFX1 \registers_reg[3][4]  ( .D(n8240), .E(n393), .CK(clk), .Q(
        \registers[3][4] ) );
  EDFFX1 \registers_reg[3][3]  ( .D(n8189), .E(n393), .CK(clk), .Q(
        \registers[3][3] ) );
  EDFFX1 \registers_reg[3][2]  ( .D(n8141), .E(n393), .CK(clk), .Q(
        \registers[3][2] ) );
  EDFFX1 \registers_reg[3][1]  ( .D(n8085), .E(n393), .CK(clk), .Q(
        \registers[3][1] ) );
  EDFFX1 \registers_reg[3][0]  ( .D(n8025), .E(n393), .CK(clk), .Q(
        \registers[3][0] ) );
  EDFFX1 \registers_reg[1020][7]  ( .D(n8397), .E(n930), .CK(clk), .Q(
        \registers[1020][7] ) );
  EDFFX1 \registers_reg[1020][6]  ( .D(n8339), .E(n930), .CK(clk), .Q(
        \registers[1020][6] ) );
  EDFFX1 \registers_reg[1020][5]  ( .D(n8281), .E(n930), .CK(clk), .Q(
        \registers[1020][5] ) );
  EDFFX1 \registers_reg[1020][4]  ( .D(n8223), .E(n930), .CK(clk), .Q(
        \registers[1020][4] ) );
  EDFFX1 \registers_reg[1020][3]  ( .D(n8178), .E(n930), .CK(clk), .Q(
        \registers[1020][3] ) );
  EDFFX1 \registers_reg[1020][2]  ( .D(n8127), .E(n930), .CK(clk), .Q(
        \registers[1020][2] ) );
  EDFFX1 \registers_reg[1020][1]  ( .D(n8071), .E(n930), .CK(clk), .Q(
        \registers[1020][1] ) );
  EDFFX1 \registers_reg[1020][0]  ( .D(n8010), .E(n930), .CK(clk), .Q(
        \registers[1020][0] ) );
  EDFFX1 \registers_reg[1016][7]  ( .D(n8395), .E(n926), .CK(clk), .Q(
        \registers[1016][7] ) );
  EDFFX1 \registers_reg[1016][6]  ( .D(n8337), .E(n926), .CK(clk), .Q(
        \registers[1016][6] ) );
  EDFFX1 \registers_reg[1016][5]  ( .D(n8279), .E(n926), .CK(clk), .Q(
        \registers[1016][5] ) );
  EDFFX1 \registers_reg[1016][4]  ( .D(n8221), .E(n926), .CK(clk), .Q(
        \registers[1016][4] ) );
  EDFFX1 \registers_reg[1016][3]  ( .D(n8176), .E(n926), .CK(clk), .Q(
        \registers[1016][3] ) );
  EDFFX1 \registers_reg[1016][2]  ( .D(n8128), .E(n926), .CK(clk), .Q(
        \registers[1016][2] ) );
  EDFFX1 \registers_reg[1016][1]  ( .D(n8072), .E(n926), .CK(clk), .Q(
        \registers[1016][1] ) );
  EDFFX1 \registers_reg[1016][0]  ( .D(n8011), .E(n926), .CK(clk), .Q(
        \registers[1016][0] ) );
  EDFFX1 \registers_reg[1012][7]  ( .D(n8396), .E(n922), .CK(clk), .Q(
        \registers[1012][7] ) );
  EDFFX1 \registers_reg[1012][6]  ( .D(n8338), .E(n922), .CK(clk), .Q(
        \registers[1012][6] ) );
  EDFFX1 \registers_reg[1012][5]  ( .D(n8280), .E(n922), .CK(clk), .Q(
        \registers[1012][5] ) );
  EDFFX1 \registers_reg[1012][4]  ( .D(n8222), .E(n922), .CK(clk), .Q(
        \registers[1012][4] ) );
  EDFFX1 \registers_reg[1012][3]  ( .D(n8177), .E(n922), .CK(clk), .Q(
        \registers[1012][3] ) );
  EDFFX1 \registers_reg[1012][2]  ( .D(n8126), .E(n922), .CK(clk), .Q(
        \registers[1012][2] ) );
  EDFFX1 \registers_reg[1012][1]  ( .D(n8070), .E(n922), .CK(clk), .Q(
        \registers[1012][1] ) );
  EDFFX1 \registers_reg[1012][0]  ( .D(n8012), .E(n922), .CK(clk), .Q(
        \registers[1012][0] ) );
  EDFFX1 \registers_reg[1008][7]  ( .D(n8397), .E(n235), .CK(clk), .Q(
        \registers[1008][7] ) );
  EDFFX1 \registers_reg[1008][6]  ( .D(n8339), .E(n235), .CK(clk), .Q(
        \registers[1008][6] ) );
  EDFFX1 \registers_reg[1008][5]  ( .D(n8281), .E(n235), .CK(clk), .Q(
        \registers[1008][5] ) );
  EDFFX1 \registers_reg[1008][4]  ( .D(n8223), .E(n235), .CK(clk), .Q(
        \registers[1008][4] ) );
  EDFFX1 \registers_reg[1008][3]  ( .D(n8178), .E(n235), .CK(clk), .Q(
        \registers[1008][3] ) );
  EDFFX1 \registers_reg[1008][2]  ( .D(n8127), .E(n235), .CK(clk), .Q(
        \registers[1008][2] ) );
  EDFFX1 \registers_reg[1008][1]  ( .D(n8071), .E(n235), .CK(clk), .Q(
        \registers[1008][1] ) );
  EDFFX1 \registers_reg[1008][0]  ( .D(n8010), .E(n235), .CK(clk), .Q(
        \registers[1008][0] ) );
  EDFFX1 \registers_reg[1004][7]  ( .D(n8395), .E(n231), .CK(clk), .Q(
        \registers[1004][7] ) );
  EDFFX1 \registers_reg[1004][6]  ( .D(n8337), .E(n231), .CK(clk), .Q(
        \registers[1004][6] ) );
  EDFFX1 \registers_reg[1004][5]  ( .D(n8279), .E(n231), .CK(clk), .Q(
        \registers[1004][5] ) );
  EDFFX1 \registers_reg[1004][4]  ( .D(n8221), .E(n231), .CK(clk), .Q(
        \registers[1004][4] ) );
  EDFFX1 \registers_reg[1004][3]  ( .D(n8173), .E(n231), .CK(clk), .Q(
        \registers[1004][3] ) );
  EDFFX1 \registers_reg[1004][2]  ( .D(n8128), .E(n231), .CK(clk), .Q(
        \registers[1004][2] ) );
  EDFFX1 \registers_reg[1004][1]  ( .D(n8072), .E(n231), .CK(clk), .Q(
        \registers[1004][1] ) );
  EDFFX1 \registers_reg[1004][0]  ( .D(n8011), .E(n231), .CK(clk), .Q(
        \registers[1004][0] ) );
  EDFFX1 \registers_reg[1000][7]  ( .D(n8396), .E(n227), .CK(clk), .Q(
        \registers[1000][7] ) );
  EDFFX1 \registers_reg[1000][6]  ( .D(n8338), .E(n227), .CK(clk), .Q(
        \registers[1000][6] ) );
  EDFFX1 \registers_reg[1000][5]  ( .D(n8280), .E(n227), .CK(clk), .Q(
        \registers[1000][5] ) );
  EDFFX1 \registers_reg[1000][4]  ( .D(n8222), .E(n227), .CK(clk), .Q(
        \registers[1000][4] ) );
  EDFFX1 \registers_reg[1000][3]  ( .D(n8174), .E(n227), .CK(clk), .Q(
        \registers[1000][3] ) );
  EDFFX1 \registers_reg[1000][2]  ( .D(n8126), .E(n227), .CK(clk), .Q(
        \registers[1000][2] ) );
  EDFFX1 \registers_reg[1000][1]  ( .D(n8070), .E(n227), .CK(clk), .Q(
        \registers[1000][1] ) );
  EDFFX1 \registers_reg[1000][0]  ( .D(n8012), .E(n227), .CK(clk), .Q(
        \registers[1000][0] ) );
  EDFFX1 \registers_reg[996][7]  ( .D(n8397), .E(n383), .CK(clk), .Q(
        \registers[996][7] ) );
  EDFFX1 \registers_reg[996][6]  ( .D(n8339), .E(n383), .CK(clk), .Q(
        \registers[996][6] ) );
  EDFFX1 \registers_reg[996][5]  ( .D(n8281), .E(n383), .CK(clk), .Q(
        \registers[996][5] ) );
  EDFFX1 \registers_reg[996][4]  ( .D(n8223), .E(n383), .CK(clk), .Q(
        \registers[996][4] ) );
  EDFFX1 \registers_reg[996][3]  ( .D(n8175), .E(n383), .CK(clk), .Q(
        \registers[996][3] ) );
  EDFFX1 \registers_reg[996][2]  ( .D(n8127), .E(n383), .CK(clk), .Q(
        \registers[996][2] ) );
  EDFFX1 \registers_reg[996][1]  ( .D(n8071), .E(n383), .CK(clk), .Q(
        \registers[996][1] ) );
  EDFFX1 \registers_reg[996][0]  ( .D(n8010), .E(n383), .CK(clk), .Q(
        \registers[996][0] ) );
  EDFFX1 \registers_reg[992][7]  ( .D(n8395), .E(n1013), .CK(clk), .Q(
        \registers[992][7] ) );
  EDFFX1 \registers_reg[992][6]  ( .D(n8337), .E(n1013), .CK(clk), .Q(
        \registers[992][6] ) );
  EDFFX1 \registers_reg[992][5]  ( .D(n8279), .E(n1013), .CK(clk), .Q(
        \registers[992][5] ) );
  EDFFX1 \registers_reg[992][4]  ( .D(n8221), .E(n1013), .CK(clk), .Q(
        \registers[992][4] ) );
  EDFFX1 \registers_reg[992][3]  ( .D(n8173), .E(n1013), .CK(clk), .Q(
        \registers[992][3] ) );
  EDFFX1 \registers_reg[992][2]  ( .D(n8128), .E(n1013), .CK(clk), .Q(
        \registers[992][2] ) );
  EDFFX1 \registers_reg[992][1]  ( .D(n8072), .E(n1013), .CK(clk), .Q(
        \registers[992][1] ) );
  EDFFX1 \registers_reg[992][0]  ( .D(n8011), .E(n1013), .CK(clk), .Q(
        \registers[992][0] ) );
  EDFFX1 \registers_reg[988][7]  ( .D(n8396), .E(n918), .CK(clk), .Q(
        \registers[988][7] ) );
  EDFFX1 \registers_reg[988][6]  ( .D(n8338), .E(n918), .CK(clk), .Q(
        \registers[988][6] ) );
  EDFFX1 \registers_reg[988][5]  ( .D(n8280), .E(n918), .CK(clk), .Q(
        \registers[988][5] ) );
  EDFFX1 \registers_reg[988][4]  ( .D(n8222), .E(n918), .CK(clk), .Q(
        \registers[988][4] ) );
  EDFFX1 \registers_reg[988][3]  ( .D(n8174), .E(n918), .CK(clk), .Q(
        \registers[988][3] ) );
  EDFFX1 \registers_reg[988][2]  ( .D(n8126), .E(n918), .CK(clk), .Q(
        \registers[988][2] ) );
  EDFFX1 \registers_reg[988][1]  ( .D(n8070), .E(n918), .CK(clk), .Q(
        \registers[988][1] ) );
  EDFFX1 \registers_reg[988][0]  ( .D(n8012), .E(n918), .CK(clk), .Q(
        \registers[988][0] ) );
  EDFFX1 \registers_reg[984][7]  ( .D(n8397), .E(n914), .CK(clk), .Q(
        \registers[984][7] ) );
  EDFFX1 \registers_reg[984][6]  ( .D(n8339), .E(n914), .CK(clk), .Q(
        \registers[984][6] ) );
  EDFFX1 \registers_reg[984][5]  ( .D(n8281), .E(n914), .CK(clk), .Q(
        \registers[984][5] ) );
  EDFFX1 \registers_reg[984][4]  ( .D(n8223), .E(n914), .CK(clk), .Q(
        \registers[984][4] ) );
  EDFFX1 \registers_reg[984][3]  ( .D(n8175), .E(n914), .CK(clk), .Q(
        \registers[984][3] ) );
  EDFFX1 \registers_reg[984][2]  ( .D(n8124), .E(n914), .CK(clk), .Q(
        \registers[984][2] ) );
  EDFFX1 \registers_reg[984][1]  ( .D(n8068), .E(n914), .CK(clk), .Q(
        \registers[984][1] ) );
  EDFFX1 \registers_reg[984][0]  ( .D(n8007), .E(n914), .CK(clk), .Q(
        \registers[984][0] ) );
  EDFFX1 \registers_reg[980][7]  ( .D(n8395), .E(n910), .CK(clk), .Q(
        \registers[980][7] ) );
  EDFFX1 \registers_reg[980][6]  ( .D(n8337), .E(n910), .CK(clk), .Q(
        \registers[980][6] ) );
  EDFFX1 \registers_reg[980][5]  ( .D(n8279), .E(n910), .CK(clk), .Q(
        \registers[980][5] ) );
  EDFFX1 \registers_reg[980][4]  ( .D(n8221), .E(n910), .CK(clk), .Q(
        \registers[980][4] ) );
  EDFFX1 \registers_reg[980][3]  ( .D(n8173), .E(n910), .CK(clk), .Q(
        \registers[980][3] ) );
  EDFFX1 \registers_reg[980][2]  ( .D(n8125), .E(n910), .CK(clk), .Q(
        \registers[980][2] ) );
  EDFFX1 \registers_reg[980][1]  ( .D(n8069), .E(n910), .CK(clk), .Q(
        \registers[980][1] ) );
  EDFFX1 \registers_reg[980][0]  ( .D(n8008), .E(n910), .CK(clk), .Q(
        \registers[980][0] ) );
  EDFFX1 \registers_reg[976][7]  ( .D(n8394), .E(n223), .CK(clk), .Q(
        \registers[976][7] ) );
  EDFFX1 \registers_reg[976][6]  ( .D(n8336), .E(n223), .CK(clk), .Q(
        \registers[976][6] ) );
  EDFFX1 \registers_reg[976][5]  ( .D(n8278), .E(n223), .CK(clk), .Q(
        \registers[976][5] ) );
  EDFFX1 \registers_reg[976][4]  ( .D(n8220), .E(n223), .CK(clk), .Q(
        \registers[976][4] ) );
  EDFFX1 \registers_reg[976][3]  ( .D(n8174), .E(n223), .CK(clk), .Q(
        \registers[976][3] ) );
  EDFFX1 \registers_reg[976][2]  ( .D(n8123), .E(n223), .CK(clk), .Q(
        \registers[976][2] ) );
  EDFFX1 \registers_reg[976][1]  ( .D(n8067), .E(n223), .CK(clk), .Q(
        \registers[976][1] ) );
  EDFFX1 \registers_reg[976][0]  ( .D(n8009), .E(n223), .CK(clk), .Q(
        \registers[976][0] ) );
  EDFFX1 \registers_reg[972][7]  ( .D(n8392), .E(n219), .CK(clk), .Q(
        \registers[972][7] ) );
  EDFFX1 \registers_reg[972][6]  ( .D(n8334), .E(n219), .CK(clk), .Q(
        \registers[972][6] ) );
  EDFFX1 \registers_reg[972][5]  ( .D(n8276), .E(n219), .CK(clk), .Q(
        \registers[972][5] ) );
  EDFFX1 \registers_reg[972][4]  ( .D(n8218), .E(n219), .CK(clk), .Q(
        \registers[972][4] ) );
  EDFFX1 \registers_reg[972][3]  ( .D(n8175), .E(n219), .CK(clk), .Q(
        \registers[972][3] ) );
  EDFFX1 \registers_reg[972][2]  ( .D(n8124), .E(n219), .CK(clk), .Q(
        \registers[972][2] ) );
  EDFFX1 \registers_reg[972][1]  ( .D(n8068), .E(n219), .CK(clk), .Q(
        \registers[972][1] ) );
  EDFFX1 \registers_reg[972][0]  ( .D(n8007), .E(n219), .CK(clk), .Q(
        \registers[972][0] ) );
  EDFFX1 \registers_reg[968][7]  ( .D(n8393), .E(n215), .CK(clk), .Q(
        \registers[968][7] ) );
  EDFFX1 \registers_reg[968][6]  ( .D(n8335), .E(n215), .CK(clk), .Q(
        \registers[968][6] ) );
  EDFFX1 \registers_reg[968][5]  ( .D(n8277), .E(n215), .CK(clk), .Q(
        \registers[968][5] ) );
  EDFFX1 \registers_reg[968][4]  ( .D(n8219), .E(n215), .CK(clk), .Q(
        \registers[968][4] ) );
  EDFFX1 \registers_reg[968][3]  ( .D(n8173), .E(n215), .CK(clk), .Q(
        \registers[968][3] ) );
  EDFFX1 \registers_reg[968][2]  ( .D(n8125), .E(n215), .CK(clk), .Q(
        \registers[968][2] ) );
  EDFFX1 \registers_reg[968][1]  ( .D(n8069), .E(n215), .CK(clk), .Q(
        \registers[968][1] ) );
  EDFFX1 \registers_reg[968][0]  ( .D(n8008), .E(n215), .CK(clk), .Q(
        \registers[968][0] ) );
  EDFFX1 \registers_reg[964][7]  ( .D(n8394), .E(n376), .CK(clk), .Q(
        \registers[964][7] ) );
  EDFFX1 \registers_reg[964][6]  ( .D(n8336), .E(n376), .CK(clk), .Q(
        \registers[964][6] ) );
  EDFFX1 \registers_reg[964][5]  ( .D(n8278), .E(n376), .CK(clk), .Q(
        \registers[964][5] ) );
  EDFFX1 \registers_reg[964][4]  ( .D(n8220), .E(n376), .CK(clk), .Q(
        \registers[964][4] ) );
  EDFFX1 \registers_reg[964][3]  ( .D(n8174), .E(n376), .CK(clk), .Q(
        \registers[964][3] ) );
  EDFFX1 \registers_reg[964][2]  ( .D(n8123), .E(n376), .CK(clk), .Q(
        \registers[964][2] ) );
  EDFFX1 \registers_reg[964][1]  ( .D(n8067), .E(n376), .CK(clk), .Q(
        \registers[964][1] ) );
  EDFFX1 \registers_reg[964][0]  ( .D(n8009), .E(n376), .CK(clk), .Q(
        \registers[964][0] ) );
  EDFFX1 \registers_reg[960][7]  ( .D(n8392), .E(n1012), .CK(clk), .Q(
        \registers[960][7] ) );
  EDFFX1 \registers_reg[960][6]  ( .D(n8334), .E(n1012), .CK(clk), .Q(
        \registers[960][6] ) );
  EDFFX1 \registers_reg[960][5]  ( .D(n8276), .E(n1012), .CK(clk), .Q(
        \registers[960][5] ) );
  EDFFX1 \registers_reg[960][4]  ( .D(n8218), .E(n1012), .CK(clk), .Q(
        \registers[960][4] ) );
  EDFFX1 \registers_reg[960][3]  ( .D(n8175), .E(n1012), .CK(clk), .Q(
        \registers[960][3] ) );
  EDFFX1 \registers_reg[960][2]  ( .D(n8124), .E(n1012), .CK(clk), .Q(
        \registers[960][2] ) );
  EDFFX1 \registers_reg[960][1]  ( .D(n8068), .E(n1012), .CK(clk), .Q(
        \registers[960][1] ) );
  EDFFX1 \registers_reg[960][0]  ( .D(n8007), .E(n1012), .CK(clk), .Q(
        \registers[960][0] ) );
  EDFFX1 \registers_reg[956][7]  ( .D(n8394), .E(n906), .CK(clk), .Q(
        \registers[956][7] ) );
  EDFFX1 \registers_reg[956][6]  ( .D(n8336), .E(n906), .CK(clk), .Q(
        \registers[956][6] ) );
  EDFFX1 \registers_reg[956][5]  ( .D(n8278), .E(n906), .CK(clk), .Q(
        \registers[956][5] ) );
  EDFFX1 \registers_reg[956][4]  ( .D(n8220), .E(n906), .CK(clk), .Q(
        \registers[956][4] ) );
  EDFFX1 \registers_reg[956][3]  ( .D(n8174), .E(n906), .CK(clk), .Q(
        \registers[956][3] ) );
  EDFFX1 \registers_reg[956][2]  ( .D(n8123), .E(n906), .CK(clk), .Q(
        \registers[956][2] ) );
  EDFFX1 \registers_reg[956][1]  ( .D(n8067), .E(n906), .CK(clk), .Q(
        \registers[956][1] ) );
  EDFFX1 \registers_reg[956][0]  ( .D(n8009), .E(n906), .CK(clk), .Q(
        \registers[956][0] ) );
  EDFFX1 \registers_reg[952][7]  ( .D(n8392), .E(n902), .CK(clk), .Q(
        \registers[952][7] ) );
  EDFFX1 \registers_reg[952][6]  ( .D(n8334), .E(n902), .CK(clk), .Q(
        \registers[952][6] ) );
  EDFFX1 \registers_reg[952][5]  ( .D(n8276), .E(n902), .CK(clk), .Q(
        \registers[952][5] ) );
  EDFFX1 \registers_reg[952][4]  ( .D(n8218), .E(n902), .CK(clk), .Q(
        \registers[952][4] ) );
  EDFFX1 \registers_reg[952][3]  ( .D(n8175), .E(n902), .CK(clk), .Q(
        \registers[952][3] ) );
  EDFFX1 \registers_reg[952][2]  ( .D(n8124), .E(n902), .CK(clk), .Q(
        \registers[952][2] ) );
  EDFFX1 \registers_reg[952][1]  ( .D(n8068), .E(n902), .CK(clk), .Q(
        \registers[952][1] ) );
  EDFFX1 \registers_reg[952][0]  ( .D(n8007), .E(n902), .CK(clk), .Q(
        \registers[952][0] ) );
  EDFFX1 \registers_reg[948][7]  ( .D(n8393), .E(n898), .CK(clk), .Q(
        \registers[948][7] ) );
  EDFFX1 \registers_reg[948][6]  ( .D(n8335), .E(n898), .CK(clk), .Q(
        \registers[948][6] ) );
  EDFFX1 \registers_reg[948][5]  ( .D(n8277), .E(n898), .CK(clk), .Q(
        \registers[948][5] ) );
  EDFFX1 \registers_reg[948][4]  ( .D(n8219), .E(n898), .CK(clk), .Q(
        \registers[948][4] ) );
  EDFFX1 \registers_reg[948][3]  ( .D(n8173), .E(n898), .CK(clk), .Q(
        \registers[948][3] ) );
  EDFFX1 \registers_reg[948][2]  ( .D(n8125), .E(n898), .CK(clk), .Q(
        \registers[948][2] ) );
  EDFFX1 \registers_reg[948][1]  ( .D(n8069), .E(n898), .CK(clk), .Q(
        \registers[948][1] ) );
  EDFFX1 \registers_reg[948][0]  ( .D(n8008), .E(n898), .CK(clk), .Q(
        \registers[948][0] ) );
  EDFFX1 \registers_reg[944][7]  ( .D(n8394), .E(n211), .CK(clk), .Q(
        \registers[944][7] ) );
  EDFFX1 \registers_reg[944][6]  ( .D(n8336), .E(n211), .CK(clk), .Q(
        \registers[944][6] ) );
  EDFFX1 \registers_reg[944][5]  ( .D(n8278), .E(n211), .CK(clk), .Q(
        \registers[944][5] ) );
  EDFFX1 \registers_reg[944][4]  ( .D(n8220), .E(n211), .CK(clk), .Q(
        \registers[944][4] ) );
  EDFFX1 \registers_reg[944][3]  ( .D(n8174), .E(n211), .CK(clk), .Q(
        \registers[944][3] ) );
  EDFFX1 \registers_reg[944][2]  ( .D(n8123), .E(n211), .CK(clk), .Q(
        \registers[944][2] ) );
  EDFFX1 \registers_reg[944][1]  ( .D(n8067), .E(n211), .CK(clk), .Q(
        \registers[944][1] ) );
  EDFFX1 \registers_reg[944][0]  ( .D(n8009), .E(n211), .CK(clk), .Q(
        \registers[944][0] ) );
  EDFFX1 \registers_reg[940][7]  ( .D(n8392), .E(n207), .CK(clk), .Q(
        \registers[940][7] ) );
  EDFFX1 \registers_reg[940][6]  ( .D(n8334), .E(n207), .CK(clk), .Q(
        \registers[940][6] ) );
  EDFFX1 \registers_reg[940][5]  ( .D(n8276), .E(n207), .CK(clk), .Q(
        \registers[940][5] ) );
  EDFFX1 \registers_reg[940][4]  ( .D(n8218), .E(n207), .CK(clk), .Q(
        \registers[940][4] ) );
  EDFFX1 \registers_reg[940][3]  ( .D(n8172), .E(n207), .CK(clk), .Q(
        \registers[940][3] ) );
  EDFFX1 \registers_reg[940][2]  ( .D(n8124), .E(n207), .CK(clk), .Q(
        \registers[940][2] ) );
  EDFFX1 \registers_reg[940][1]  ( .D(n8068), .E(n207), .CK(clk), .Q(
        \registers[940][1] ) );
  EDFFX1 \registers_reg[940][0]  ( .D(n8007), .E(n207), .CK(clk), .Q(
        \registers[940][0] ) );
  EDFFX1 \registers_reg[936][7]  ( .D(n8393), .E(n203), .CK(clk), .Q(
        \registers[936][7] ) );
  EDFFX1 \registers_reg[936][6]  ( .D(n8335), .E(n203), .CK(clk), .Q(
        \registers[936][6] ) );
  EDFFX1 \registers_reg[936][5]  ( .D(n8277), .E(n203), .CK(clk), .Q(
        \registers[936][5] ) );
  EDFFX1 \registers_reg[936][4]  ( .D(n8219), .E(n203), .CK(clk), .Q(
        \registers[936][4] ) );
  EDFFX1 \registers_reg[936][3]  ( .D(n8170), .E(n203), .CK(clk), .Q(
        \registers[936][3] ) );
  EDFFX1 \registers_reg[936][2]  ( .D(n8125), .E(n203), .CK(clk), .Q(
        \registers[936][2] ) );
  EDFFX1 \registers_reg[936][1]  ( .D(n8069), .E(n203), .CK(clk), .Q(
        \registers[936][1] ) );
  EDFFX1 \registers_reg[936][0]  ( .D(n8008), .E(n203), .CK(clk), .Q(
        \registers[936][0] ) );
  EDFFX1 \registers_reg[932][7]  ( .D(n8394), .E(n369), .CK(clk), .Q(
        \registers[932][7] ) );
  EDFFX1 \registers_reg[932][6]  ( .D(n8336), .E(n369), .CK(clk), .Q(
        \registers[932][6] ) );
  EDFFX1 \registers_reg[932][5]  ( .D(n8278), .E(n369), .CK(clk), .Q(
        \registers[932][5] ) );
  EDFFX1 \registers_reg[932][4]  ( .D(n8220), .E(n369), .CK(clk), .Q(
        \registers[932][4] ) );
  EDFFX1 \registers_reg[932][3]  ( .D(n8171), .E(n369), .CK(clk), .Q(
        \registers[932][3] ) );
  EDFFX1 \registers_reg[932][2]  ( .D(n8120), .E(n369), .CK(clk), .Q(
        \registers[932][2] ) );
  EDFFX1 \registers_reg[932][1]  ( .D(n8064), .E(n369), .CK(clk), .Q(
        \registers[932][1] ) );
  EDFFX1 \registers_reg[932][0]  ( .D(n8006), .E(n369), .CK(clk), .Q(
        \registers[932][0] ) );
  EDFFX1 \registers_reg[928][7]  ( .D(n8390), .E(n1011), .CK(clk), .Q(
        \registers[928][7] ) );
  EDFFX1 \registers_reg[928][6]  ( .D(n8332), .E(n1011), .CK(clk), .Q(
        \registers[928][6] ) );
  EDFFX1 \registers_reg[928][5]  ( .D(n8274), .E(n1011), .CK(clk), .Q(
        \registers[928][5] ) );
  EDFFX1 \registers_reg[928][4]  ( .D(n8216), .E(n1011), .CK(clk), .Q(
        \registers[928][4] ) );
  EDFFX1 \registers_reg[928][3]  ( .D(n8172), .E(n1011), .CK(clk), .Q(
        \registers[928][3] ) );
  EDFFX1 \registers_reg[928][2]  ( .D(n8121), .E(n1011), .CK(clk), .Q(
        \registers[928][2] ) );
  EDFFX1 \registers_reg[928][1]  ( .D(n8065), .E(n1011), .CK(clk), .Q(
        \registers[928][1] ) );
  EDFFX1 \registers_reg[928][0]  ( .D(n8004), .E(n1011), .CK(clk), .Q(
        \registers[928][0] ) );
  EDFFX1 \registers_reg[924][7]  ( .D(n8391), .E(n894), .CK(clk), .Q(
        \registers[924][7] ) );
  EDFFX1 \registers_reg[924][6]  ( .D(n8333), .E(n894), .CK(clk), .Q(
        \registers[924][6] ) );
  EDFFX1 \registers_reg[924][5]  ( .D(n8275), .E(n894), .CK(clk), .Q(
        \registers[924][5] ) );
  EDFFX1 \registers_reg[924][4]  ( .D(n8217), .E(n894), .CK(clk), .Q(
        \registers[924][4] ) );
  EDFFX1 \registers_reg[924][3]  ( .D(n8170), .E(n894), .CK(clk), .Q(
        \registers[924][3] ) );
  EDFFX1 \registers_reg[924][2]  ( .D(n8122), .E(n894), .CK(clk), .Q(
        \registers[924][2] ) );
  EDFFX1 \registers_reg[924][1]  ( .D(n8066), .E(n894), .CK(clk), .Q(
        \registers[924][1] ) );
  EDFFX1 \registers_reg[924][0]  ( .D(n8005), .E(n894), .CK(clk), .Q(
        \registers[924][0] ) );
  EDFFX1 \registers_reg[920][7]  ( .D(n8389), .E(n890), .CK(clk), .Q(
        \registers[920][7] ) );
  EDFFX1 \registers_reg[920][6]  ( .D(n8331), .E(n890), .CK(clk), .Q(
        \registers[920][6] ) );
  EDFFX1 \registers_reg[920][5]  ( .D(n8273), .E(n890), .CK(clk), .Q(
        \registers[920][5] ) );
  EDFFX1 \registers_reg[920][4]  ( .D(n8215), .E(n890), .CK(clk), .Q(
        \registers[920][4] ) );
  EDFFX1 \registers_reg[920][3]  ( .D(n8171), .E(n890), .CK(clk), .Q(
        \registers[920][3] ) );
  EDFFX1 \registers_reg[920][2]  ( .D(n8120), .E(n890), .CK(clk), .Q(
        \registers[920][2] ) );
  EDFFX1 \registers_reg[920][1]  ( .D(n8064), .E(n890), .CK(clk), .Q(
        \registers[920][1] ) );
  EDFFX1 \registers_reg[920][0]  ( .D(n8006), .E(n890), .CK(clk), .Q(
        \registers[920][0] ) );
  EDFFX1 \registers_reg[916][7]  ( .D(n8390), .E(n886), .CK(clk), .Q(
        \registers[916][7] ) );
  EDFFX1 \registers_reg[916][6]  ( .D(n8332), .E(n886), .CK(clk), .Q(
        \registers[916][6] ) );
  EDFFX1 \registers_reg[916][5]  ( .D(n8274), .E(n886), .CK(clk), .Q(
        \registers[916][5] ) );
  EDFFX1 \registers_reg[916][4]  ( .D(n8216), .E(n886), .CK(clk), .Q(
        \registers[916][4] ) );
  EDFFX1 \registers_reg[916][3]  ( .D(n8172), .E(n886), .CK(clk), .Q(
        \registers[916][3] ) );
  EDFFX1 \registers_reg[916][2]  ( .D(n8121), .E(n886), .CK(clk), .Q(
        \registers[916][2] ) );
  EDFFX1 \registers_reg[916][1]  ( .D(n8065), .E(n886), .CK(clk), .Q(
        \registers[916][1] ) );
  EDFFX1 \registers_reg[916][0]  ( .D(n8004), .E(n886), .CK(clk), .Q(
        \registers[916][0] ) );
  EDFFX1 \registers_reg[912][7]  ( .D(n8391), .E(n199), .CK(clk), .Q(
        \registers[912][7] ) );
  EDFFX1 \registers_reg[912][6]  ( .D(n8333), .E(n199), .CK(clk), .Q(
        \registers[912][6] ) );
  EDFFX1 \registers_reg[912][5]  ( .D(n8275), .E(n199), .CK(clk), .Q(
        \registers[912][5] ) );
  EDFFX1 \registers_reg[912][4]  ( .D(n8217), .E(n199), .CK(clk), .Q(
        \registers[912][4] ) );
  EDFFX1 \registers_reg[912][3]  ( .D(n8170), .E(n199), .CK(clk), .Q(
        \registers[912][3] ) );
  EDFFX1 \registers_reg[912][2]  ( .D(n8122), .E(n199), .CK(clk), .Q(
        \registers[912][2] ) );
  EDFFX1 \registers_reg[912][1]  ( .D(n8066), .E(n199), .CK(clk), .Q(
        \registers[912][1] ) );
  EDFFX1 \registers_reg[912][0]  ( .D(n8005), .E(n199), .CK(clk), .Q(
        \registers[912][0] ) );
  EDFFX1 \registers_reg[908][7]  ( .D(n8389), .E(n195), .CK(clk), .Q(
        \registers[908][7] ) );
  EDFFX1 \registers_reg[908][6]  ( .D(n8331), .E(n195), .CK(clk), .Q(
        \registers[908][6] ) );
  EDFFX1 \registers_reg[908][5]  ( .D(n8273), .E(n195), .CK(clk), .Q(
        \registers[908][5] ) );
  EDFFX1 \registers_reg[908][4]  ( .D(n8215), .E(n195), .CK(clk), .Q(
        \registers[908][4] ) );
  EDFFX1 \registers_reg[908][3]  ( .D(n8171), .E(n195), .CK(clk), .Q(
        \registers[908][3] ) );
  EDFFX1 \registers_reg[908][2]  ( .D(n8120), .E(n195), .CK(clk), .Q(
        \registers[908][2] ) );
  EDFFX1 \registers_reg[908][1]  ( .D(n8064), .E(n195), .CK(clk), .Q(
        \registers[908][1] ) );
  EDFFX1 \registers_reg[908][0]  ( .D(n8006), .E(n195), .CK(clk), .Q(
        \registers[908][0] ) );
  EDFFX1 \registers_reg[904][7]  ( .D(n8390), .E(n191), .CK(clk), .Q(
        \registers[904][7] ) );
  EDFFX1 \registers_reg[904][6]  ( .D(n8332), .E(n191), .CK(clk), .Q(
        \registers[904][6] ) );
  EDFFX1 \registers_reg[904][5]  ( .D(n8274), .E(n191), .CK(clk), .Q(
        \registers[904][5] ) );
  EDFFX1 \registers_reg[904][4]  ( .D(n8216), .E(n191), .CK(clk), .Q(
        \registers[904][4] ) );
  EDFFX1 \registers_reg[904][3]  ( .D(n8172), .E(n191), .CK(clk), .Q(
        \registers[904][3] ) );
  EDFFX1 \registers_reg[904][2]  ( .D(n8121), .E(n191), .CK(clk), .Q(
        \registers[904][2] ) );
  EDFFX1 \registers_reg[904][1]  ( .D(n8065), .E(n191), .CK(clk), .Q(
        \registers[904][1] ) );
  EDFFX1 \registers_reg[904][0]  ( .D(n8004), .E(n191), .CK(clk), .Q(
        \registers[904][0] ) );
  EDFFX1 \registers_reg[900][7]  ( .D(n8391), .E(n362), .CK(clk), .Q(
        \registers[900][7] ) );
  EDFFX1 \registers_reg[900][6]  ( .D(n8333), .E(n362), .CK(clk), .Q(
        \registers[900][6] ) );
  EDFFX1 \registers_reg[900][5]  ( .D(n8275), .E(n362), .CK(clk), .Q(
        \registers[900][5] ) );
  EDFFX1 \registers_reg[900][4]  ( .D(n8217), .E(n362), .CK(clk), .Q(
        \registers[900][4] ) );
  EDFFX1 \registers_reg[900][3]  ( .D(n8170), .E(n362), .CK(clk), .Q(
        \registers[900][3] ) );
  EDFFX1 \registers_reg[900][2]  ( .D(n8122), .E(n362), .CK(clk), .Q(
        \registers[900][2] ) );
  EDFFX1 \registers_reg[900][1]  ( .D(n8066), .E(n362), .CK(clk), .Q(
        \registers[900][1] ) );
  EDFFX1 \registers_reg[900][0]  ( .D(n8005), .E(n362), .CK(clk), .Q(
        \registers[900][0] ) );
  EDFFX1 \registers_reg[896][7]  ( .D(n8389), .E(n1010), .CK(clk), .Q(
        \registers[896][7] ) );
  EDFFX1 \registers_reg[896][6]  ( .D(n8331), .E(n1010), .CK(clk), .Q(
        \registers[896][6] ) );
  EDFFX1 \registers_reg[896][5]  ( .D(n8273), .E(n1010), .CK(clk), .Q(
        \registers[896][5] ) );
  EDFFX1 \registers_reg[896][4]  ( .D(n8215), .E(n1010), .CK(clk), .Q(
        \registers[896][4] ) );
  EDFFX1 \registers_reg[896][3]  ( .D(n8171), .E(n1010), .CK(clk), .Q(
        \registers[896][3] ) );
  EDFFX1 \registers_reg[896][2]  ( .D(n8120), .E(n1010), .CK(clk), .Q(
        \registers[896][2] ) );
  EDFFX1 \registers_reg[896][1]  ( .D(n8064), .E(n1010), .CK(clk), .Q(
        \registers[896][1] ) );
  EDFFX1 \registers_reg[896][0]  ( .D(n8006), .E(n1010), .CK(clk), .Q(
        \registers[896][0] ) );
  EDFFX1 \registers_reg[892][7]  ( .D(n8405), .E(n882), .CK(clk), .Q(
        \registers[892][7] ) );
  EDFFX1 \registers_reg[892][6]  ( .D(n8347), .E(n882), .CK(clk), .Q(
        \registers[892][6] ) );
  EDFFX1 \registers_reg[892][5]  ( .D(n8289), .E(n882), .CK(clk), .Q(
        \registers[892][5] ) );
  EDFFX1 \registers_reg[892][4]  ( .D(n8231), .E(n882), .CK(clk), .Q(
        \registers[892][4] ) );
  EDFFX1 \registers_reg[892][3]  ( .D(n8183), .E(n882), .CK(clk), .Q(
        \registers[892][3] ) );
  EDFFX1 \registers_reg[892][2]  ( .D(n8135), .E(n882), .CK(clk), .Q(
        \registers[892][2] ) );
  EDFFX1 \registers_reg[892][1]  ( .D(n8079), .E(n882), .CK(clk), .Q(
        \registers[892][1] ) );
  EDFFX1 \registers_reg[892][0]  ( .D(n8021), .E(n882), .CK(clk), .Q(
        \registers[892][0] ) );
  EDFFX1 \registers_reg[888][7]  ( .D(n8406), .E(n878), .CK(clk), .Q(
        \registers[888][7] ) );
  EDFFX1 \registers_reg[888][6]  ( .D(n8348), .E(n878), .CK(clk), .Q(
        \registers[888][6] ) );
  EDFFX1 \registers_reg[888][5]  ( .D(n8290), .E(n878), .CK(clk), .Q(
        \registers[888][5] ) );
  EDFFX1 \registers_reg[888][4]  ( .D(n8232), .E(n878), .CK(clk), .Q(
        \registers[888][4] ) );
  EDFFX1 \registers_reg[888][3]  ( .D(n8184), .E(n878), .CK(clk), .Q(
        \registers[888][3] ) );
  EDFFX1 \registers_reg[888][2]  ( .D(n8136), .E(n878), .CK(clk), .Q(
        \registers[888][2] ) );
  EDFFX1 \registers_reg[888][1]  ( .D(n8080), .E(n878), .CK(clk), .Q(
        \registers[888][1] ) );
  EDFFX1 \registers_reg[888][0]  ( .D(n8019), .E(n878), .CK(clk), .Q(
        \registers[888][0] ) );
  EDFFX1 \registers_reg[884][7]  ( .D(n8404), .E(n874), .CK(clk), .Q(
        \registers[884][7] ) );
  EDFFX1 \registers_reg[884][6]  ( .D(n8346), .E(n874), .CK(clk), .Q(
        \registers[884][6] ) );
  EDFFX1 \registers_reg[884][5]  ( .D(n8288), .E(n874), .CK(clk), .Q(
        \registers[884][5] ) );
  EDFFX1 \registers_reg[884][4]  ( .D(n8230), .E(n874), .CK(clk), .Q(
        \registers[884][4] ) );
  EDFFX1 \registers_reg[884][3]  ( .D(n8182), .E(n874), .CK(clk), .Q(
        \registers[884][3] ) );
  EDFFX1 \registers_reg[884][2]  ( .D(n8137), .E(n874), .CK(clk), .Q(
        \registers[884][2] ) );
  EDFFX1 \registers_reg[884][1]  ( .D(n8081), .E(n874), .CK(clk), .Q(
        \registers[884][1] ) );
  EDFFX1 \registers_reg[884][0]  ( .D(n8020), .E(n874), .CK(clk), .Q(
        \registers[884][0] ) );
  EDFFX1 \registers_reg[880][7]  ( .D(n8405), .E(n187), .CK(clk), .Q(
        \registers[880][7] ) );
  EDFFX1 \registers_reg[880][6]  ( .D(n8347), .E(n187), .CK(clk), .Q(
        \registers[880][6] ) );
  EDFFX1 \registers_reg[880][5]  ( .D(n8289), .E(n187), .CK(clk), .Q(
        \registers[880][5] ) );
  EDFFX1 \registers_reg[880][4]  ( .D(n8231), .E(n187), .CK(clk), .Q(
        \registers[880][4] ) );
  EDFFX1 \registers_reg[880][3]  ( .D(n8183), .E(n187), .CK(clk), .Q(
        \registers[880][3] ) );
  EDFFX1 \registers_reg[880][2]  ( .D(n8132), .E(n187), .CK(clk), .Q(
        \registers[880][2] ) );
  EDFFX1 \registers_reg[880][1]  ( .D(n8076), .E(n187), .CK(clk), .Q(
        \registers[880][1] ) );
  EDFFX1 \registers_reg[880][0]  ( .D(n8018), .E(n187), .CK(clk), .Q(
        \registers[880][0] ) );
  EDFFX1 \registers_reg[876][7]  ( .D(n8406), .E(n183), .CK(clk), .Q(
        \registers[876][7] ) );
  EDFFX1 \registers_reg[876][6]  ( .D(n8348), .E(n183), .CK(clk), .Q(
        \registers[876][6] ) );
  EDFFX1 \registers_reg[876][5]  ( .D(n8290), .E(n183), .CK(clk), .Q(
        \registers[876][5] ) );
  EDFFX1 \registers_reg[876][4]  ( .D(n8232), .E(n183), .CK(clk), .Q(
        \registers[876][4] ) );
  EDFFX1 \registers_reg[876][3]  ( .D(n8184), .E(n183), .CK(clk), .Q(
        \registers[876][3] ) );
  EDFFX1 \registers_reg[876][2]  ( .D(n8133), .E(n183), .CK(clk), .Q(
        \registers[876][2] ) );
  EDFFX1 \registers_reg[876][1]  ( .D(n8077), .E(n183), .CK(clk), .Q(
        \registers[876][1] ) );
  EDFFX1 \registers_reg[876][0]  ( .D(n8016), .E(n183), .CK(clk), .Q(
        \registers[876][0] ) );
  EDFFX1 \registers_reg[872][7]  ( .D(n8402), .E(n179), .CK(clk), .Q(
        \registers[872][7] ) );
  EDFFX1 \registers_reg[872][6]  ( .D(n8344), .E(n179), .CK(clk), .Q(
        \registers[872][6] ) );
  EDFFX1 \registers_reg[872][5]  ( .D(n8286), .E(n179), .CK(clk), .Q(
        \registers[872][5] ) );
  EDFFX1 \registers_reg[872][4]  ( .D(n8228), .E(n179), .CK(clk), .Q(
        \registers[872][4] ) );
  EDFFX1 \registers_reg[872][3]  ( .D(n8179), .E(n179), .CK(clk), .Q(
        \registers[872][3] ) );
  EDFFX1 \registers_reg[872][2]  ( .D(n8134), .E(n179), .CK(clk), .Q(
        \registers[872][2] ) );
  EDFFX1 \registers_reg[872][1]  ( .D(n8078), .E(n179), .CK(clk), .Q(
        \registers[872][1] ) );
  EDFFX1 \registers_reg[872][0]  ( .D(n8017), .E(n179), .CK(clk), .Q(
        \registers[872][0] ) );
  EDFFX1 \registers_reg[868][7]  ( .D(n8403), .E(n355), .CK(clk), .Q(
        \registers[868][7] ) );
  EDFFX1 \registers_reg[868][6]  ( .D(n8345), .E(n355), .CK(clk), .Q(
        \registers[868][6] ) );
  EDFFX1 \registers_reg[868][5]  ( .D(n8287), .E(n355), .CK(clk), .Q(
        \registers[868][5] ) );
  EDFFX1 \registers_reg[868][4]  ( .D(n8229), .E(n355), .CK(clk), .Q(
        \registers[868][4] ) );
  EDFFX1 \registers_reg[868][3]  ( .D(n8180), .E(n355), .CK(clk), .Q(
        \registers[868][3] ) );
  EDFFX1 \registers_reg[868][2]  ( .D(n8132), .E(n355), .CK(clk), .Q(
        \registers[868][2] ) );
  EDFFX1 \registers_reg[868][1]  ( .D(n8076), .E(n355), .CK(clk), .Q(
        \registers[868][1] ) );
  EDFFX1 \registers_reg[868][0]  ( .D(n8018), .E(n355), .CK(clk), .Q(
        \registers[868][0] ) );
  EDFFX1 \registers_reg[864][7]  ( .D(n8401), .E(n1009), .CK(clk), .Q(
        \registers[864][7] ) );
  EDFFX1 \registers_reg[864][6]  ( .D(n8343), .E(n1009), .CK(clk), .Q(
        \registers[864][6] ) );
  EDFFX1 \registers_reg[864][5]  ( .D(n8285), .E(n1009), .CK(clk), .Q(
        \registers[864][5] ) );
  EDFFX1 \registers_reg[864][4]  ( .D(n8227), .E(n1009), .CK(clk), .Q(
        \registers[864][4] ) );
  EDFFX1 \registers_reg[864][3]  ( .D(n8181), .E(n1009), .CK(clk), .Q(
        \registers[864][3] ) );
  EDFFX1 \registers_reg[864][2]  ( .D(n8133), .E(n1009), .CK(clk), .Q(
        \registers[864][2] ) );
  EDFFX1 \registers_reg[864][1]  ( .D(n8077), .E(n1009), .CK(clk), .Q(
        \registers[864][1] ) );
  EDFFX1 \registers_reg[864][0]  ( .D(n8016), .E(n1009), .CK(clk), .Q(
        \registers[864][0] ) );
  EDFFX1 \registers_reg[860][7]  ( .D(n8402), .E(n870), .CK(clk), .Q(
        \registers[860][7] ) );
  EDFFX1 \registers_reg[860][6]  ( .D(n8344), .E(n870), .CK(clk), .Q(
        \registers[860][6] ) );
  EDFFX1 \registers_reg[860][5]  ( .D(n8286), .E(n870), .CK(clk), .Q(
        \registers[860][5] ) );
  EDFFX1 \registers_reg[860][4]  ( .D(n8228), .E(n870), .CK(clk), .Q(
        \registers[860][4] ) );
  EDFFX1 \registers_reg[860][3]  ( .D(n8179), .E(n870), .CK(clk), .Q(
        \registers[860][3] ) );
  EDFFX1 \registers_reg[860][2]  ( .D(n8134), .E(n870), .CK(clk), .Q(
        \registers[860][2] ) );
  EDFFX1 \registers_reg[860][1]  ( .D(n8078), .E(n870), .CK(clk), .Q(
        \registers[860][1] ) );
  EDFFX1 \registers_reg[860][0]  ( .D(n8017), .E(n870), .CK(clk), .Q(
        \registers[860][0] ) );
  EDFFX1 \registers_reg[856][7]  ( .D(n8403), .E(n866), .CK(clk), .Q(
        \registers[856][7] ) );
  EDFFX1 \registers_reg[856][6]  ( .D(n8345), .E(n866), .CK(clk), .Q(
        \registers[856][6] ) );
  EDFFX1 \registers_reg[856][5]  ( .D(n8287), .E(n866), .CK(clk), .Q(
        \registers[856][5] ) );
  EDFFX1 \registers_reg[856][4]  ( .D(n8229), .E(n866), .CK(clk), .Q(
        \registers[856][4] ) );
  EDFFX1 \registers_reg[856][3]  ( .D(n8180), .E(n866), .CK(clk), .Q(
        \registers[856][3] ) );
  EDFFX1 \registers_reg[856][2]  ( .D(n8132), .E(n866), .CK(clk), .Q(
        \registers[856][2] ) );
  EDFFX1 \registers_reg[856][1]  ( .D(n8076), .E(n866), .CK(clk), .Q(
        \registers[856][1] ) );
  EDFFX1 \registers_reg[856][0]  ( .D(n8018), .E(n866), .CK(clk), .Q(
        \registers[856][0] ) );
  EDFFX1 \registers_reg[852][7]  ( .D(n8401), .E(n862), .CK(clk), .Q(
        \registers[852][7] ) );
  EDFFX1 \registers_reg[852][6]  ( .D(n8343), .E(n862), .CK(clk), .Q(
        \registers[852][6] ) );
  EDFFX1 \registers_reg[852][5]  ( .D(n8285), .E(n862), .CK(clk), .Q(
        \registers[852][5] ) );
  EDFFX1 \registers_reg[852][4]  ( .D(n8227), .E(n862), .CK(clk), .Q(
        \registers[852][4] ) );
  EDFFX1 \registers_reg[852][3]  ( .D(n8181), .E(n862), .CK(clk), .Q(
        \registers[852][3] ) );
  EDFFX1 \registers_reg[852][2]  ( .D(n8133), .E(n862), .CK(clk), .Q(
        \registers[852][2] ) );
  EDFFX1 \registers_reg[852][1]  ( .D(n8077), .E(n862), .CK(clk), .Q(
        \registers[852][1] ) );
  EDFFX1 \registers_reg[852][0]  ( .D(n8016), .E(n862), .CK(clk), .Q(
        \registers[852][0] ) );
  EDFFX1 \registers_reg[848][7]  ( .D(n8402), .E(n175), .CK(clk), .Q(
        \registers[848][7] ) );
  EDFFX1 \registers_reg[848][6]  ( .D(n8344), .E(n175), .CK(clk), .Q(
        \registers[848][6] ) );
  EDFFX1 \registers_reg[848][5]  ( .D(n8286), .E(n175), .CK(clk), .Q(
        \registers[848][5] ) );
  EDFFX1 \registers_reg[848][4]  ( .D(n8228), .E(n175), .CK(clk), .Q(
        \registers[848][4] ) );
  EDFFX1 \registers_reg[848][3]  ( .D(n8179), .E(n175), .CK(clk), .Q(
        \registers[848][3] ) );
  EDFFX1 \registers_reg[848][2]  ( .D(n8134), .E(n175), .CK(clk), .Q(
        \registers[848][2] ) );
  EDFFX1 \registers_reg[848][1]  ( .D(n8078), .E(n175), .CK(clk), .Q(
        \registers[848][1] ) );
  EDFFX1 \registers_reg[848][0]  ( .D(n8017), .E(n175), .CK(clk), .Q(
        \registers[848][0] ) );
  EDFFX1 \registers_reg[844][7]  ( .D(n8403), .E(n171), .CK(clk), .Q(
        \registers[844][7] ) );
  EDFFX1 \registers_reg[844][6]  ( .D(n8345), .E(n171), .CK(clk), .Q(
        \registers[844][6] ) );
  EDFFX1 \registers_reg[844][5]  ( .D(n8287), .E(n171), .CK(clk), .Q(
        \registers[844][5] ) );
  EDFFX1 \registers_reg[844][4]  ( .D(n8229), .E(n171), .CK(clk), .Q(
        \registers[844][4] ) );
  EDFFX1 \registers_reg[844][3]  ( .D(n8180), .E(n171), .CK(clk), .Q(
        \registers[844][3] ) );
  EDFFX1 \registers_reg[844][2]  ( .D(n8132), .E(n171), .CK(clk), .Q(
        \registers[844][2] ) );
  EDFFX1 \registers_reg[844][1]  ( .D(n8076), .E(n171), .CK(clk), .Q(
        \registers[844][1] ) );
  EDFFX1 \registers_reg[844][0]  ( .D(n8018), .E(n171), .CK(clk), .Q(
        \registers[844][0] ) );
  EDFFX1 \registers_reg[840][7]  ( .D(n8401), .E(n167), .CK(clk), .Q(
        \registers[840][7] ) );
  EDFFX1 \registers_reg[840][6]  ( .D(n8343), .E(n167), .CK(clk), .Q(
        \registers[840][6] ) );
  EDFFX1 \registers_reg[840][5]  ( .D(n8285), .E(n167), .CK(clk), .Q(
        \registers[840][5] ) );
  EDFFX1 \registers_reg[840][4]  ( .D(n8227), .E(n167), .CK(clk), .Q(
        \registers[840][4] ) );
  EDFFX1 \registers_reg[840][3]  ( .D(n8181), .E(n167), .CK(clk), .Q(
        \registers[840][3] ) );
  EDFFX1 \registers_reg[840][2]  ( .D(n8133), .E(n167), .CK(clk), .Q(
        \registers[840][2] ) );
  EDFFX1 \registers_reg[840][1]  ( .D(n8077), .E(n167), .CK(clk), .Q(
        \registers[840][1] ) );
  EDFFX1 \registers_reg[840][0]  ( .D(n8016), .E(n167), .CK(clk), .Q(
        \registers[840][0] ) );
  EDFFX1 \registers_reg[836][7]  ( .D(n8402), .E(n348), .CK(clk), .Q(
        \registers[836][7] ) );
  EDFFX1 \registers_reg[836][6]  ( .D(n8344), .E(n348), .CK(clk), .Q(
        \registers[836][6] ) );
  EDFFX1 \registers_reg[836][5]  ( .D(n8286), .E(n348), .CK(clk), .Q(
        \registers[836][5] ) );
  EDFFX1 \registers_reg[836][4]  ( .D(n8228), .E(n348), .CK(clk), .Q(
        \registers[836][4] ) );
  EDFFX1 \registers_reg[836][3]  ( .D(n8179), .E(n348), .CK(clk), .Q(
        \registers[836][3] ) );
  EDFFX1 \registers_reg[836][2]  ( .D(n8134), .E(n348), .CK(clk), .Q(
        \registers[836][2] ) );
  EDFFX1 \registers_reg[836][1]  ( .D(n8078), .E(n348), .CK(clk), .Q(
        \registers[836][1] ) );
  EDFFX1 \registers_reg[836][0]  ( .D(n8017), .E(n348), .CK(clk), .Q(
        \registers[836][0] ) );
  EDFFX1 \registers_reg[832][7]  ( .D(n8403), .E(n1008), .CK(clk), .Q(
        \registers[832][7] ) );
  EDFFX1 \registers_reg[832][6]  ( .D(n8345), .E(n1008), .CK(clk), .Q(
        \registers[832][6] ) );
  EDFFX1 \registers_reg[832][5]  ( .D(n8287), .E(n1008), .CK(clk), .Q(
        \registers[832][5] ) );
  EDFFX1 \registers_reg[832][4]  ( .D(n8229), .E(n1008), .CK(clk), .Q(
        \registers[832][4] ) );
  EDFFX1 \registers_reg[832][3]  ( .D(n8180), .E(n1008), .CK(clk), .Q(
        \registers[832][3] ) );
  EDFFX1 \registers_reg[832][2]  ( .D(n8129), .E(n1008), .CK(clk), .Q(
        \registers[832][2] ) );
  EDFFX1 \registers_reg[832][1]  ( .D(n8073), .E(n1008), .CK(clk), .Q(
        \registers[832][1] ) );
  EDFFX1 \registers_reg[832][0]  ( .D(n8018), .E(n1008), .CK(clk), .Q(
        \registers[832][0] ) );
  EDFFX1 \registers_reg[828][7]  ( .D(n8402), .E(n858), .CK(clk), .Q(
        \registers[828][7] ) );
  EDFFX1 \registers_reg[828][6]  ( .D(n8344), .E(n858), .CK(clk), .Q(
        \registers[828][6] ) );
  EDFFX1 \registers_reg[828][5]  ( .D(n8286), .E(n858), .CK(clk), .Q(
        \registers[828][5] ) );
  EDFFX1 \registers_reg[828][4]  ( .D(n8228), .E(n858), .CK(clk), .Q(
        \registers[828][4] ) );
  EDFFX1 \registers_reg[828][3]  ( .D(n8179), .E(n858), .CK(clk), .Q(
        \registers[828][3] ) );
  EDFFX1 \registers_reg[828][2]  ( .D(n8131), .E(n858), .CK(clk), .Q(
        \registers[828][2] ) );
  EDFFX1 \registers_reg[828][1]  ( .D(n8075), .E(n858), .CK(clk), .Q(
        \registers[828][1] ) );
  EDFFX1 \registers_reg[828][0]  ( .D(n8014), .E(n858), .CK(clk), .Q(
        \registers[828][0] ) );
  EDFFX1 \registers_reg[824][7]  ( .D(n8398), .E(n854), .CK(clk), .Q(
        \registers[824][7] ) );
  EDFFX1 \registers_reg[824][6]  ( .D(n8340), .E(n854), .CK(clk), .Q(
        \registers[824][6] ) );
  EDFFX1 \registers_reg[824][5]  ( .D(n8282), .E(n854), .CK(clk), .Q(
        \registers[824][5] ) );
  EDFFX1 \registers_reg[824][4]  ( .D(n8224), .E(n854), .CK(clk), .Q(
        \registers[824][4] ) );
  EDFFX1 \registers_reg[824][3]  ( .D(n8180), .E(n854), .CK(clk), .Q(
        \registers[824][3] ) );
  EDFFX1 \registers_reg[824][2]  ( .D(n8129), .E(n854), .CK(clk), .Q(
        \registers[824][2] ) );
  EDFFX1 \registers_reg[824][1]  ( .D(n8073), .E(n854), .CK(clk), .Q(
        \registers[824][1] ) );
  EDFFX1 \registers_reg[824][0]  ( .D(n8015), .E(n854), .CK(clk), .Q(
        \registers[824][0] ) );
  EDFFX1 \registers_reg[820][7]  ( .D(n8399), .E(n850), .CK(clk), .Q(
        \registers[820][7] ) );
  EDFFX1 \registers_reg[820][6]  ( .D(n8341), .E(n850), .CK(clk), .Q(
        \registers[820][6] ) );
  EDFFX1 \registers_reg[820][5]  ( .D(n8283), .E(n850), .CK(clk), .Q(
        \registers[820][5] ) );
  EDFFX1 \registers_reg[820][4]  ( .D(n8225), .E(n850), .CK(clk), .Q(
        \registers[820][4] ) );
  EDFFX1 \registers_reg[820][3]  ( .D(n8181), .E(n850), .CK(clk), .Q(
        \registers[820][3] ) );
  EDFFX1 \registers_reg[820][2]  ( .D(n8130), .E(n850), .CK(clk), .Q(
        \registers[820][2] ) );
  EDFFX1 \registers_reg[820][1]  ( .D(n8074), .E(n850), .CK(clk), .Q(
        \registers[820][1] ) );
  EDFFX1 \registers_reg[820][0]  ( .D(n8013), .E(n850), .CK(clk), .Q(
        \registers[820][0] ) );
  EDFFX1 \registers_reg[816][7]  ( .D(n8400), .E(n163), .CK(clk), .Q(
        \registers[816][7] ) );
  EDFFX1 \registers_reg[816][6]  ( .D(n8342), .E(n163), .CK(clk), .Q(
        \registers[816][6] ) );
  EDFFX1 \registers_reg[816][5]  ( .D(n8284), .E(n163), .CK(clk), .Q(
        \registers[816][5] ) );
  EDFFX1 \registers_reg[816][4]  ( .D(n8226), .E(n163), .CK(clk), .Q(
        \registers[816][4] ) );
  EDFFX1 \registers_reg[816][3]  ( .D(n8179), .E(n163), .CK(clk), .Q(
        \registers[816][3] ) );
  EDFFX1 \registers_reg[816][2]  ( .D(n8131), .E(n163), .CK(clk), .Q(
        \registers[816][2] ) );
  EDFFX1 \registers_reg[816][1]  ( .D(n8075), .E(n163), .CK(clk), .Q(
        \registers[816][1] ) );
  EDFFX1 \registers_reg[816][0]  ( .D(n8014), .E(n163), .CK(clk), .Q(
        \registers[816][0] ) );
  EDFFX1 \registers_reg[812][7]  ( .D(n8398), .E(n159), .CK(clk), .Q(
        \registers[812][7] ) );
  EDFFX1 \registers_reg[812][6]  ( .D(n8340), .E(n159), .CK(clk), .Q(
        \registers[812][6] ) );
  EDFFX1 \registers_reg[812][5]  ( .D(n8282), .E(n159), .CK(clk), .Q(
        \registers[812][5] ) );
  EDFFX1 \registers_reg[812][4]  ( .D(n8224), .E(n159), .CK(clk), .Q(
        \registers[812][4] ) );
  EDFFX1 \registers_reg[812][3]  ( .D(n8177), .E(n159), .CK(clk), .Q(
        \registers[812][3] ) );
  EDFFX1 \registers_reg[812][2]  ( .D(n8129), .E(n159), .CK(clk), .Q(
        \registers[812][2] ) );
  EDFFX1 \registers_reg[812][1]  ( .D(n8073), .E(n159), .CK(clk), .Q(
        \registers[812][1] ) );
  EDFFX1 \registers_reg[812][0]  ( .D(n8015), .E(n159), .CK(clk), .Q(
        \registers[812][0] ) );
  EDFFX1 \registers_reg[808][7]  ( .D(n8399), .E(n155), .CK(clk), .Q(
        \registers[808][7] ) );
  EDFFX1 \registers_reg[808][6]  ( .D(n8341), .E(n155), .CK(clk), .Q(
        \registers[808][6] ) );
  EDFFX1 \registers_reg[808][5]  ( .D(n8283), .E(n155), .CK(clk), .Q(
        \registers[808][5] ) );
  EDFFX1 \registers_reg[808][4]  ( .D(n8225), .E(n155), .CK(clk), .Q(
        \registers[808][4] ) );
  EDFFX1 \registers_reg[808][3]  ( .D(n8178), .E(n155), .CK(clk), .Q(
        \registers[808][3] ) );
  EDFFX1 \registers_reg[808][2]  ( .D(n8130), .E(n155), .CK(clk), .Q(
        \registers[808][2] ) );
  EDFFX1 \registers_reg[808][1]  ( .D(n8074), .E(n155), .CK(clk), .Q(
        \registers[808][1] ) );
  EDFFX1 \registers_reg[808][0]  ( .D(n8013), .E(n155), .CK(clk), .Q(
        \registers[808][0] ) );
  EDFFX1 \registers_reg[804][7]  ( .D(n8400), .E(n326), .CK(clk), .Q(
        \registers[804][7] ) );
  EDFFX1 \registers_reg[804][6]  ( .D(n8342), .E(n326), .CK(clk), .Q(
        \registers[804][6] ) );
  EDFFX1 \registers_reg[804][5]  ( .D(n8284), .E(n326), .CK(clk), .Q(
        \registers[804][5] ) );
  EDFFX1 \registers_reg[804][4]  ( .D(n8226), .E(n326), .CK(clk), .Q(
        \registers[804][4] ) );
  EDFFX1 \registers_reg[804][3]  ( .D(n8176), .E(n326), .CK(clk), .Q(
        \registers[804][3] ) );
  EDFFX1 \registers_reg[804][2]  ( .D(n8131), .E(n326), .CK(clk), .Q(
        \registers[804][2] ) );
  EDFFX1 \registers_reg[804][1]  ( .D(n8075), .E(n326), .CK(clk), .Q(
        \registers[804][1] ) );
  EDFFX1 \registers_reg[804][0]  ( .D(n8014), .E(n326), .CK(clk), .Q(
        \registers[804][0] ) );
  EDFFX1 \registers_reg[800][7]  ( .D(n8398), .E(n1007), .CK(clk), .Q(
        \registers[800][7] ) );
  EDFFX1 \registers_reg[800][6]  ( .D(n8340), .E(n1007), .CK(clk), .Q(
        \registers[800][6] ) );
  EDFFX1 \registers_reg[800][5]  ( .D(n8282), .E(n1007), .CK(clk), .Q(
        \registers[800][5] ) );
  EDFFX1 \registers_reg[800][4]  ( .D(n8224), .E(n1007), .CK(clk), .Q(
        \registers[800][4] ) );
  EDFFX1 \registers_reg[800][3]  ( .D(n8177), .E(n1007), .CK(clk), .Q(
        \registers[800][3] ) );
  EDFFX1 \registers_reg[800][2]  ( .D(n8129), .E(n1007), .CK(clk), .Q(
        \registers[800][2] ) );
  EDFFX1 \registers_reg[800][1]  ( .D(n8073), .E(n1007), .CK(clk), .Q(
        \registers[800][1] ) );
  EDFFX1 \registers_reg[800][0]  ( .D(n8015), .E(n1007), .CK(clk), .Q(
        \registers[800][0] ) );
  EDFFX1 \registers_reg[796][7]  ( .D(n8399), .E(n846), .CK(clk), .Q(
        \registers[796][7] ) );
  EDFFX1 \registers_reg[796][6]  ( .D(n8341), .E(n846), .CK(clk), .Q(
        \registers[796][6] ) );
  EDFFX1 \registers_reg[796][5]  ( .D(n8283), .E(n846), .CK(clk), .Q(
        \registers[796][5] ) );
  EDFFX1 \registers_reg[796][4]  ( .D(n8225), .E(n846), .CK(clk), .Q(
        \registers[796][4] ) );
  EDFFX1 \registers_reg[796][3]  ( .D(n8178), .E(n846), .CK(clk), .Q(
        \registers[796][3] ) );
  EDFFX1 \registers_reg[796][2]  ( .D(n8130), .E(n846), .CK(clk), .Q(
        \registers[796][2] ) );
  EDFFX1 \registers_reg[796][1]  ( .D(n8074), .E(n846), .CK(clk), .Q(
        \registers[796][1] ) );
  EDFFX1 \registers_reg[796][0]  ( .D(n8013), .E(n846), .CK(clk), .Q(
        \registers[796][0] ) );
  EDFFX1 \registers_reg[792][7]  ( .D(n8400), .E(n842), .CK(clk), .Q(
        \registers[792][7] ) );
  EDFFX1 \registers_reg[792][6]  ( .D(n8342), .E(n842), .CK(clk), .Q(
        \registers[792][6] ) );
  EDFFX1 \registers_reg[792][5]  ( .D(n8284), .E(n842), .CK(clk), .Q(
        \registers[792][5] ) );
  EDFFX1 \registers_reg[792][4]  ( .D(n8226), .E(n842), .CK(clk), .Q(
        \registers[792][4] ) );
  EDFFX1 \registers_reg[792][3]  ( .D(n8176), .E(n842), .CK(clk), .Q(
        \registers[792][3] ) );
  EDFFX1 \registers_reg[792][2]  ( .D(n8131), .E(n842), .CK(clk), .Q(
        \registers[792][2] ) );
  EDFFX1 \registers_reg[792][1]  ( .D(n8075), .E(n842), .CK(clk), .Q(
        \registers[792][1] ) );
  EDFFX1 \registers_reg[792][0]  ( .D(n8014), .E(n842), .CK(clk), .Q(
        \registers[792][0] ) );
  EDFFX1 \registers_reg[788][7]  ( .D(n8398), .E(n838), .CK(clk), .Q(
        \registers[788][7] ) );
  EDFFX1 \registers_reg[788][6]  ( .D(n8340), .E(n838), .CK(clk), .Q(
        \registers[788][6] ) );
  EDFFX1 \registers_reg[788][5]  ( .D(n8282), .E(n838), .CK(clk), .Q(
        \registers[788][5] ) );
  EDFFX1 \registers_reg[788][4]  ( .D(n8224), .E(n838), .CK(clk), .Q(
        \registers[788][4] ) );
  EDFFX1 \registers_reg[788][3]  ( .D(n8177), .E(n838), .CK(clk), .Q(
        \registers[788][3] ) );
  EDFFX1 \registers_reg[788][2]  ( .D(n8129), .E(n838), .CK(clk), .Q(
        \registers[788][2] ) );
  EDFFX1 \registers_reg[788][1]  ( .D(n8073), .E(n838), .CK(clk), .Q(
        \registers[788][1] ) );
  EDFFX1 \registers_reg[788][0]  ( .D(n8015), .E(n838), .CK(clk), .Q(
        \registers[788][0] ) );
  EDFFX1 \registers_reg[784][7]  ( .D(n8399), .E(n151), .CK(clk), .Q(
        \registers[784][7] ) );
  EDFFX1 \registers_reg[784][6]  ( .D(n8341), .E(n151), .CK(clk), .Q(
        \registers[784][6] ) );
  EDFFX1 \registers_reg[784][5]  ( .D(n8283), .E(n151), .CK(clk), .Q(
        \registers[784][5] ) );
  EDFFX1 \registers_reg[784][4]  ( .D(n8225), .E(n151), .CK(clk), .Q(
        \registers[784][4] ) );
  EDFFX1 \registers_reg[784][3]  ( .D(n8178), .E(n151), .CK(clk), .Q(
        \registers[784][3] ) );
  EDFFX1 \registers_reg[784][2]  ( .D(n8130), .E(n151), .CK(clk), .Q(
        \registers[784][2] ) );
  EDFFX1 \registers_reg[784][1]  ( .D(n8074), .E(n151), .CK(clk), .Q(
        \registers[784][1] ) );
  EDFFX1 \registers_reg[784][0]  ( .D(n8013), .E(n151), .CK(clk), .Q(
        \registers[784][0] ) );
  EDFFX1 \registers_reg[780][7]  ( .D(n8400), .E(n147), .CK(clk), .Q(
        \registers[780][7] ) );
  EDFFX1 \registers_reg[780][6]  ( .D(n8342), .E(n147), .CK(clk), .Q(
        \registers[780][6] ) );
  EDFFX1 \registers_reg[780][5]  ( .D(n8284), .E(n147), .CK(clk), .Q(
        \registers[780][5] ) );
  EDFFX1 \registers_reg[780][4]  ( .D(n8226), .E(n147), .CK(clk), .Q(
        \registers[780][4] ) );
  EDFFX1 \registers_reg[780][3]  ( .D(n8176), .E(n147), .CK(clk), .Q(
        \registers[780][3] ) );
  EDFFX1 \registers_reg[780][2]  ( .D(n8128), .E(n147), .CK(clk), .Q(
        \registers[780][2] ) );
  EDFFX1 \registers_reg[780][1]  ( .D(n8072), .E(n147), .CK(clk), .Q(
        \registers[780][1] ) );
  EDFFX1 \registers_reg[780][0]  ( .D(n8011), .E(n147), .CK(clk), .Q(
        \registers[780][0] ) );
  EDFFX1 \registers_reg[776][7]  ( .D(n8398), .E(n143), .CK(clk), .Q(
        \registers[776][7] ) );
  EDFFX1 \registers_reg[776][6]  ( .D(n8340), .E(n143), .CK(clk), .Q(
        \registers[776][6] ) );
  EDFFX1 \registers_reg[776][5]  ( .D(n8282), .E(n143), .CK(clk), .Q(
        \registers[776][5] ) );
  EDFFX1 \registers_reg[776][4]  ( .D(n8224), .E(n143), .CK(clk), .Q(
        \registers[776][4] ) );
  EDFFX1 \registers_reg[776][3]  ( .D(n8177), .E(n143), .CK(clk), .Q(
        \registers[776][3] ) );
  EDFFX1 \registers_reg[776][2]  ( .D(n8126), .E(n143), .CK(clk), .Q(
        \registers[776][2] ) );
  EDFFX1 \registers_reg[776][1]  ( .D(n8070), .E(n143), .CK(clk), .Q(
        \registers[776][1] ) );
  EDFFX1 \registers_reg[776][0]  ( .D(n8012), .E(n143), .CK(clk), .Q(
        \registers[776][0] ) );
  EDFFX1 \registers_reg[772][7]  ( .D(n8397), .E(n319), .CK(clk), .Q(
        \registers[772][7] ) );
  EDFFX1 \registers_reg[772][6]  ( .D(n8339), .E(n319), .CK(clk), .Q(
        \registers[772][6] ) );
  EDFFX1 \registers_reg[772][5]  ( .D(n8281), .E(n319), .CK(clk), .Q(
        \registers[772][5] ) );
  EDFFX1 \registers_reg[772][4]  ( .D(n8223), .E(n319), .CK(clk), .Q(
        \registers[772][4] ) );
  EDFFX1 \registers_reg[772][3]  ( .D(n8178), .E(n319), .CK(clk), .Q(
        \registers[772][3] ) );
  EDFFX1 \registers_reg[772][2]  ( .D(n8127), .E(n319), .CK(clk), .Q(
        \registers[772][2] ) );
  EDFFX1 \registers_reg[772][1]  ( .D(n8071), .E(n319), .CK(clk), .Q(
        \registers[772][1] ) );
  EDFFX1 \registers_reg[772][0]  ( .D(n8010), .E(n319), .CK(clk), .Q(
        \registers[772][0] ) );
  EDFFX1 \registers_reg[768][7]  ( .D(n8395), .E(n1006), .CK(clk), .Q(
        \registers[768][7] ) );
  EDFFX1 \registers_reg[768][6]  ( .D(n8337), .E(n1006), .CK(clk), .Q(
        \registers[768][6] ) );
  EDFFX1 \registers_reg[768][5]  ( .D(n8279), .E(n1006), .CK(clk), .Q(
        \registers[768][5] ) );
  EDFFX1 \registers_reg[768][4]  ( .D(n8221), .E(n1006), .CK(clk), .Q(
        \registers[768][4] ) );
  EDFFX1 \registers_reg[768][3]  ( .D(n8176), .E(n1006), .CK(clk), .Q(
        \registers[768][3] ) );
  EDFFX1 \registers_reg[768][2]  ( .D(n8128), .E(n1006), .CK(clk), .Q(
        \registers[768][2] ) );
  EDFFX1 \registers_reg[768][1]  ( .D(n8072), .E(n1006), .CK(clk), .Q(
        \registers[768][1] ) );
  EDFFX1 \registers_reg[768][0]  ( .D(n8011), .E(n1006), .CK(clk), .Q(
        \registers[768][0] ) );
  EDFFX1 \registers_reg[764][7]  ( .D(n8381), .E(n834), .CK(clk), .Q(
        \registers[764][7] ) );
  EDFFX1 \registers_reg[764][6]  ( .D(n8323), .E(n834), .CK(clk), .Q(
        \registers[764][6] ) );
  EDFFX1 \registers_reg[764][5]  ( .D(n8265), .E(n834), .CK(clk), .Q(
        \registers[764][5] ) );
  EDFFX1 \registers_reg[764][4]  ( .D(n8207), .E(n834), .CK(clk), .Q(
        \registers[764][4] ) );
  EDFFX1 \registers_reg[764][3]  ( .D(n8165), .E(n834), .CK(clk), .Q(
        \registers[764][3] ) );
  EDFFX1 \registers_reg[764][2]  ( .D(n8111), .E(n834), .CK(clk), .Q(
        \registers[764][2] ) );
  EDFFX1 \registers_reg[764][1]  ( .D(n8055), .E(n834), .CK(clk), .Q(
        \registers[764][1] ) );
  EDFFX1 \registers_reg[764][0]  ( .D(n8679), .E(n834), .CK(clk), .Q(
        \registers[764][0] ) );
  EDFFX1 \registers_reg[760][7]  ( .D(n8382), .E(n830), .CK(clk), .Q(
        \registers[760][7] ) );
  EDFFX1 \registers_reg[760][6]  ( .D(n8324), .E(n830), .CK(clk), .Q(
        \registers[760][6] ) );
  EDFFX1 \registers_reg[760][5]  ( .D(n8266), .E(n830), .CK(clk), .Q(
        \registers[760][5] ) );
  EDFFX1 \registers_reg[760][4]  ( .D(n8208), .E(n830), .CK(clk), .Q(
        \registers[760][4] ) );
  EDFFX1 \registers_reg[760][3]  ( .D(n8166), .E(n830), .CK(clk), .Q(
        \registers[760][3] ) );
  EDFFX1 \registers_reg[760][2]  ( .D(n8112), .E(n830), .CK(clk), .Q(
        \registers[760][2] ) );
  EDFFX1 \registers_reg[760][1]  ( .D(n8056), .E(n830), .CK(clk), .Q(
        \registers[760][1] ) );
  EDFFX1 \registers_reg[760][0]  ( .D(n7996), .E(n830), .CK(clk), .Q(
        \registers[760][0] ) );
  EDFFX1 \registers_reg[756][7]  ( .D(n8383), .E(n826), .CK(clk), .Q(
        \registers[756][7] ) );
  EDFFX1 \registers_reg[756][6]  ( .D(n8325), .E(n826), .CK(clk), .Q(
        \registers[756][6] ) );
  EDFFX1 \registers_reg[756][5]  ( .D(n8267), .E(n826), .CK(clk), .Q(
        \registers[756][5] ) );
  EDFFX1 \registers_reg[756][4]  ( .D(n8209), .E(n826), .CK(clk), .Q(
        \registers[756][4] ) );
  EDFFX1 \registers_reg[756][3]  ( .D(n8164), .E(n826), .CK(clk), .Q(
        \registers[756][3] ) );
  EDFFX1 \registers_reg[756][2]  ( .D(n8113), .E(n826), .CK(clk), .Q(
        \registers[756][2] ) );
  EDFFX1 \registers_reg[756][1]  ( .D(n8057), .E(n826), .CK(clk), .Q(
        \registers[756][1] ) );
  EDFFX1 \registers_reg[756][0]  ( .D(n7997), .E(n826), .CK(clk), .Q(
        \registers[756][0] ) );
  EDFFX1 \registers_reg[752][7]  ( .D(n8381), .E(n139), .CK(clk), .Q(
        \registers[752][7] ) );
  EDFFX1 \registers_reg[752][6]  ( .D(n8323), .E(n139), .CK(clk), .Q(
        \registers[752][6] ) );
  EDFFX1 \registers_reg[752][5]  ( .D(n8265), .E(n139), .CK(clk), .Q(
        \registers[752][5] ) );
  EDFFX1 \registers_reg[752][4]  ( .D(n8207), .E(n139), .CK(clk), .Q(
        \registers[752][4] ) );
  EDFFX1 \registers_reg[752][3]  ( .D(n8162), .E(n139), .CK(clk), .Q(
        \registers[752][3] ) );
  EDFFX1 \registers_reg[752][2]  ( .D(n8111), .E(n139), .CK(clk), .Q(
        \registers[752][2] ) );
  EDFFX1 \registers_reg[752][1]  ( .D(n8055), .E(n139), .CK(clk), .Q(
        \registers[752][1] ) );
  EDFFX1 \registers_reg[752][0]  ( .D(n8680), .E(n139), .CK(clk), .Q(
        \registers[752][0] ) );
  EDFFX1 \registers_reg[748][7]  ( .D(n8382), .E(n135), .CK(clk), .Q(
        \registers[748][7] ) );
  EDFFX1 \registers_reg[748][6]  ( .D(n8324), .E(n135), .CK(clk), .Q(
        \registers[748][6] ) );
  EDFFX1 \registers_reg[748][5]  ( .D(n8266), .E(n135), .CK(clk), .Q(
        \registers[748][5] ) );
  EDFFX1 \registers_reg[748][4]  ( .D(n8208), .E(n135), .CK(clk), .Q(
        \registers[748][4] ) );
  EDFFX1 \registers_reg[748][3]  ( .D(n8163), .E(n135), .CK(clk), .Q(
        \registers[748][3] ) );
  EDFFX1 \registers_reg[748][2]  ( .D(n8112), .E(n135), .CK(clk), .Q(
        \registers[748][2] ) );
  EDFFX1 \registers_reg[748][1]  ( .D(n8056), .E(n135), .CK(clk), .Q(
        \registers[748][1] ) );
  EDFFX1 \registers_reg[748][0]  ( .D(n7996), .E(n135), .CK(clk), .Q(
        \registers[748][0] ) );
  EDFFX1 \registers_reg[744][7]  ( .D(n8383), .E(n131), .CK(clk), .Q(
        \registers[744][7] ) );
  EDFFX1 \registers_reg[744][6]  ( .D(n8325), .E(n131), .CK(clk), .Q(
        \registers[744][6] ) );
  EDFFX1 \registers_reg[744][5]  ( .D(n8267), .E(n131), .CK(clk), .Q(
        \registers[744][5] ) );
  EDFFX1 \registers_reg[744][4]  ( .D(n8209), .E(n131), .CK(clk), .Q(
        \registers[744][4] ) );
  EDFFX1 \registers_reg[744][3]  ( .D(n8755), .E(n131), .CK(clk), .Q(
        \registers[744][3] ) );
  EDFFX1 \registers_reg[744][2]  ( .D(n8113), .E(n131), .CK(clk), .Q(
        \registers[744][2] ) );
  EDFFX1 \registers_reg[744][1]  ( .D(n8057), .E(n131), .CK(clk), .Q(
        \registers[744][1] ) );
  EDFFX1 \registers_reg[744][0]  ( .D(n7997), .E(n131), .CK(clk), .Q(
        \registers[744][0] ) );
  EDFFX1 \registers_reg[740][7]  ( .D(n8381), .E(n312), .CK(clk), .Q(
        \registers[740][7] ) );
  EDFFX1 \registers_reg[740][6]  ( .D(n8323), .E(n312), .CK(clk), .Q(
        \registers[740][6] ) );
  EDFFX1 \registers_reg[740][5]  ( .D(n8265), .E(n312), .CK(clk), .Q(
        \registers[740][5] ) );
  EDFFX1 \registers_reg[740][4]  ( .D(n8207), .E(n312), .CK(clk), .Q(
        \registers[740][4] ) );
  EDFFX1 \registers_reg[740][3]  ( .D(n8162), .E(n312), .CK(clk), .Q(
        \registers[740][3] ) );
  EDFFX1 \registers_reg[740][2]  ( .D(n8111), .E(n312), .CK(clk), .Q(
        \registers[740][2] ) );
  EDFFX1 \registers_reg[740][1]  ( .D(n8055), .E(n312), .CK(clk), .Q(
        \registers[740][1] ) );
  EDFFX1 \registers_reg[740][0]  ( .D(n8674), .E(n312), .CK(clk), .Q(
        \registers[740][0] ) );
  EDFFX1 \registers_reg[736][7]  ( .D(n8382), .E(n1005), .CK(clk), .Q(
        \registers[736][7] ) );
  EDFFX1 \registers_reg[736][6]  ( .D(n8324), .E(n1005), .CK(clk), .Q(
        \registers[736][6] ) );
  EDFFX1 \registers_reg[736][5]  ( .D(n8266), .E(n1005), .CK(clk), .Q(
        \registers[736][5] ) );
  EDFFX1 \registers_reg[736][4]  ( .D(n8208), .E(n1005), .CK(clk), .Q(
        \registers[736][4] ) );
  EDFFX1 \registers_reg[736][3]  ( .D(n8163), .E(n1005), .CK(clk), .Q(
        \registers[736][3] ) );
  EDFFX1 \registers_reg[736][2]  ( .D(n8112), .E(n1005), .CK(clk), .Q(
        \registers[736][2] ) );
  EDFFX1 \registers_reg[736][1]  ( .D(n8056), .E(n1005), .CK(clk), .Q(
        \registers[736][1] ) );
  EDFFX1 \registers_reg[736][0]  ( .D(n7996), .E(n1005), .CK(clk), .Q(
        \registers[736][0] ) );
  EDFFX1 \registers_reg[732][7]  ( .D(n8383), .E(n822), .CK(clk), .Q(
        \registers[732][7] ) );
  EDFFX1 \registers_reg[732][6]  ( .D(n8325), .E(n822), .CK(clk), .Q(
        \registers[732][6] ) );
  EDFFX1 \registers_reg[732][5]  ( .D(n8267), .E(n822), .CK(clk), .Q(
        \registers[732][5] ) );
  EDFFX1 \registers_reg[732][4]  ( .D(n8209), .E(n822), .CK(clk), .Q(
        \registers[732][4] ) );
  EDFFX1 \registers_reg[732][3]  ( .D(n8768), .E(n822), .CK(clk), .Q(
        \registers[732][3] ) );
  EDFFX1 \registers_reg[732][2]  ( .D(n8113), .E(n822), .CK(clk), .Q(
        \registers[732][2] ) );
  EDFFX1 \registers_reg[732][1]  ( .D(n8057), .E(n822), .CK(clk), .Q(
        \registers[732][1] ) );
  EDFFX1 \registers_reg[732][0]  ( .D(n7997), .E(n822), .CK(clk), .Q(
        \registers[732][0] ) );
  EDFFX1 \registers_reg[728][7]  ( .D(n8379), .E(n818), .CK(clk), .Q(
        \registers[728][7] ) );
  EDFFX1 \registers_reg[728][6]  ( .D(n8321), .E(n818), .CK(clk), .Q(
        \registers[728][6] ) );
  EDFFX1 \registers_reg[728][5]  ( .D(n8263), .E(n818), .CK(clk), .Q(
        \registers[728][5] ) );
  EDFFX1 \registers_reg[728][4]  ( .D(n8205), .E(n818), .CK(clk), .Q(
        \registers[728][4] ) );
  EDFFX1 \registers_reg[728][3]  ( .D(n8162), .E(n818), .CK(clk), .Q(
        \registers[728][3] ) );
  EDFFX1 \registers_reg[728][2]  ( .D(n8108), .E(n818), .CK(clk), .Q(
        \registers[728][2] ) );
  EDFFX1 \registers_reg[728][1]  ( .D(n8052), .E(n818), .CK(clk), .Q(
        \registers[728][1] ) );
  EDFFX1 \registers_reg[728][0]  ( .D(n8040), .E(n818), .CK(clk), .Q(
        \registers[728][0] ) );
  EDFFX1 \registers_reg[724][7]  ( .D(n8380), .E(n814), .CK(clk), .Q(
        \registers[724][7] ) );
  EDFFX1 \registers_reg[724][6]  ( .D(n8322), .E(n814), .CK(clk), .Q(
        \registers[724][6] ) );
  EDFFX1 \registers_reg[724][5]  ( .D(n8264), .E(n814), .CK(clk), .Q(
        \registers[724][5] ) );
  EDFFX1 \registers_reg[724][4]  ( .D(n8206), .E(n814), .CK(clk), .Q(
        \registers[724][4] ) );
  EDFFX1 \registers_reg[724][3]  ( .D(n8163), .E(n814), .CK(clk), .Q(
        \registers[724][3] ) );
  EDFFX1 \registers_reg[724][2]  ( .D(n8109), .E(n814), .CK(clk), .Q(
        \registers[724][2] ) );
  EDFFX1 \registers_reg[724][1]  ( .D(n8053), .E(n814), .CK(clk), .Q(
        \registers[724][1] ) );
  EDFFX1 \registers_reg[724][0]  ( .D(n7995), .E(n814), .CK(clk), .Q(
        \registers[724][0] ) );
  EDFFX1 \registers_reg[720][7]  ( .D(n8378), .E(n127), .CK(clk), .Q(
        \registers[720][7] ) );
  EDFFX1 \registers_reg[720][6]  ( .D(n8320), .E(n127), .CK(clk), .Q(
        \registers[720][6] ) );
  EDFFX1 \registers_reg[720][5]  ( .D(n8262), .E(n127), .CK(clk), .Q(
        \registers[720][5] ) );
  EDFFX1 \registers_reg[720][4]  ( .D(n8204), .E(n127), .CK(clk), .Q(
        \registers[720][4] ) );
  EDFFX1 \registers_reg[720][3]  ( .D(n8751), .E(n127), .CK(clk), .Q(
        \registers[720][3] ) );
  EDFFX1 \registers_reg[720][2]  ( .D(n8110), .E(n127), .CK(clk), .Q(
        \registers[720][2] ) );
  EDFFX1 \registers_reg[720][1]  ( .D(n8054), .E(n127), .CK(clk), .Q(
        \registers[720][1] ) );
  EDFFX1 \registers_reg[720][0]  ( .D(n8017), .E(n127), .CK(clk), .Q(
        \registers[720][0] ) );
  EDFFX1 \registers_reg[716][7]  ( .D(n8379), .E(n123), .CK(clk), .Q(
        \registers[716][7] ) );
  EDFFX1 \registers_reg[716][6]  ( .D(n8321), .E(n123), .CK(clk), .Q(
        \registers[716][6] ) );
  EDFFX1 \registers_reg[716][5]  ( .D(n8263), .E(n123), .CK(clk), .Q(
        \registers[716][5] ) );
  EDFFX1 \registers_reg[716][4]  ( .D(n8205), .E(n123), .CK(clk), .Q(
        \registers[716][4] ) );
  EDFFX1 \registers_reg[716][3]  ( .D(n8162), .E(n123), .CK(clk), .Q(
        \registers[716][3] ) );
  EDFFX1 \registers_reg[716][2]  ( .D(n8108), .E(n123), .CK(clk), .Q(
        \registers[716][2] ) );
  EDFFX1 \registers_reg[716][1]  ( .D(n8052), .E(n123), .CK(clk), .Q(
        \registers[716][1] ) );
  EDFFX1 \registers_reg[716][0]  ( .D(n8044), .E(n123), .CK(clk), .Q(
        \registers[716][0] ) );
  EDFFX1 \registers_reg[712][7]  ( .D(n8380), .E(n119), .CK(clk), .Q(
        \registers[712][7] ) );
  EDFFX1 \registers_reg[712][6]  ( .D(n8322), .E(n119), .CK(clk), .Q(
        \registers[712][6] ) );
  EDFFX1 \registers_reg[712][5]  ( .D(n8264), .E(n119), .CK(clk), .Q(
        \registers[712][5] ) );
  EDFFX1 \registers_reg[712][4]  ( .D(n8206), .E(n119), .CK(clk), .Q(
        \registers[712][4] ) );
  EDFFX1 \registers_reg[712][3]  ( .D(n8163), .E(n119), .CK(clk), .Q(
        \registers[712][3] ) );
  EDFFX1 \registers_reg[712][2]  ( .D(n8109), .E(n119), .CK(clk), .Q(
        \registers[712][2] ) );
  EDFFX1 \registers_reg[712][1]  ( .D(n8053), .E(n119), .CK(clk), .Q(
        \registers[712][1] ) );
  EDFFX1 \registers_reg[712][0]  ( .D(n7995), .E(n119), .CK(clk), .Q(
        \registers[712][0] ) );
  EDFFX1 \registers_reg[708][7]  ( .D(n8378), .E(n305), .CK(clk), .Q(
        \registers[708][7] ) );
  EDFFX1 \registers_reg[708][6]  ( .D(n8320), .E(n305), .CK(clk), .Q(
        \registers[708][6] ) );
  EDFFX1 \registers_reg[708][5]  ( .D(n8262), .E(n305), .CK(clk), .Q(
        \registers[708][5] ) );
  EDFFX1 \registers_reg[708][4]  ( .D(n8204), .E(n305), .CK(clk), .Q(
        \registers[708][4] ) );
  EDFFX1 \registers_reg[708][3]  ( .D(n8759), .E(n305), .CK(clk), .Q(
        \registers[708][3] ) );
  EDFFX1 \registers_reg[708][2]  ( .D(n8110), .E(n305), .CK(clk), .Q(
        \registers[708][2] ) );
  EDFFX1 \registers_reg[708][1]  ( .D(n8054), .E(n305), .CK(clk), .Q(
        \registers[708][1] ) );
  EDFFX1 \registers_reg[708][0]  ( .D(n8018), .E(n305), .CK(clk), .Q(
        \registers[708][0] ) );
  EDFFX1 \registers_reg[704][7]  ( .D(n8379), .E(n1004), .CK(clk), .Q(
        \registers[704][7] ) );
  EDFFX1 \registers_reg[704][6]  ( .D(n8321), .E(n1004), .CK(clk), .Q(
        \registers[704][6] ) );
  EDFFX1 \registers_reg[704][5]  ( .D(n8263), .E(n1004), .CK(clk), .Q(
        \registers[704][5] ) );
  EDFFX1 \registers_reg[704][4]  ( .D(n8205), .E(n1004), .CK(clk), .Q(
        \registers[704][4] ) );
  EDFFX1 \registers_reg[704][3]  ( .D(n8162), .E(n1004), .CK(clk), .Q(
        \registers[704][3] ) );
  EDFFX1 \registers_reg[704][2]  ( .D(n8108), .E(n1004), .CK(clk), .Q(
        \registers[704][2] ) );
  EDFFX1 \registers_reg[704][1]  ( .D(n8052), .E(n1004), .CK(clk), .Q(
        \registers[704][1] ) );
  EDFFX1 \registers_reg[704][0]  ( .D(n8037), .E(n1004), .CK(clk), .Q(
        \registers[704][0] ) );
  EDFFX1 \registers_reg[700][7]  ( .D(n8378), .E(n810), .CK(clk), .Q(
        \registers[700][7] ) );
  EDFFX1 \registers_reg[700][6]  ( .D(n8320), .E(n810), .CK(clk), .Q(
        \registers[700][6] ) );
  EDFFX1 \registers_reg[700][5]  ( .D(n8262), .E(n810), .CK(clk), .Q(
        \registers[700][5] ) );
  EDFFX1 \registers_reg[700][4]  ( .D(n8204), .E(n810), .CK(clk), .Q(
        \registers[700][4] ) );
  EDFFX1 \registers_reg[700][3]  ( .D(n8758), .E(n810), .CK(clk), .Q(
        \registers[700][3] ) );
  EDFFX1 \registers_reg[700][2]  ( .D(n8110), .E(n810), .CK(clk), .Q(
        \registers[700][2] ) );
  EDFFX1 \registers_reg[700][1]  ( .D(n8054), .E(n810), .CK(clk), .Q(
        \registers[700][1] ) );
  EDFFX1 \registers_reg[700][0]  ( .D(n8027), .E(n810), .CK(clk), .Q(
        \registers[700][0] ) );
  EDFFX1 \registers_reg[696][7]  ( .D(n8379), .E(n806), .CK(clk), .Q(
        \registers[696][7] ) );
  EDFFX1 \registers_reg[696][6]  ( .D(n8321), .E(n806), .CK(clk), .Q(
        \registers[696][6] ) );
  EDFFX1 \registers_reg[696][5]  ( .D(n8263), .E(n806), .CK(clk), .Q(
        \registers[696][5] ) );
  EDFFX1 \registers_reg[696][4]  ( .D(n8205), .E(n806), .CK(clk), .Q(
        \registers[696][4] ) );
  EDFFX1 \registers_reg[696][3]  ( .D(n8162), .E(n806), .CK(clk), .Q(
        \registers[696][3] ) );
  EDFFX1 \registers_reg[696][2]  ( .D(n8108), .E(n806), .CK(clk), .Q(
        \registers[696][2] ) );
  EDFFX1 \registers_reg[696][1]  ( .D(n8052), .E(n806), .CK(clk), .Q(
        \registers[696][1] ) );
  EDFFX1 \registers_reg[696][0]  ( .D(n8038), .E(n806), .CK(clk), .Q(
        \registers[696][0] ) );
  EDFFX1 \registers_reg[692][7]  ( .D(n8380), .E(n802), .CK(clk), .Q(
        \registers[692][7] ) );
  EDFFX1 \registers_reg[692][6]  ( .D(n8322), .E(n802), .CK(clk), .Q(
        \registers[692][6] ) );
  EDFFX1 \registers_reg[692][5]  ( .D(n8264), .E(n802), .CK(clk), .Q(
        \registers[692][5] ) );
  EDFFX1 \registers_reg[692][4]  ( .D(n8206), .E(n802), .CK(clk), .Q(
        \registers[692][4] ) );
  EDFFX1 \registers_reg[692][3]  ( .D(n8163), .E(n802), .CK(clk), .Q(
        \registers[692][3] ) );
  EDFFX1 \registers_reg[692][2]  ( .D(n8109), .E(n802), .CK(clk), .Q(
        \registers[692][2] ) );
  EDFFX1 \registers_reg[692][1]  ( .D(n8053), .E(n802), .CK(clk), .Q(
        \registers[692][1] ) );
  EDFFX1 \registers_reg[692][0]  ( .D(n7995), .E(n802), .CK(clk), .Q(
        \registers[692][0] ) );
  EDFFX1 \registers_reg[688][7]  ( .D(n8378), .E(n115), .CK(clk), .Q(
        \registers[688][7] ) );
  EDFFX1 \registers_reg[688][6]  ( .D(n8320), .E(n115), .CK(clk), .Q(
        \registers[688][6] ) );
  EDFFX1 \registers_reg[688][5]  ( .D(n8262), .E(n115), .CK(clk), .Q(
        \registers[688][5] ) );
  EDFFX1 \registers_reg[688][4]  ( .D(n8204), .E(n115), .CK(clk), .Q(
        \registers[688][4] ) );
  EDFFX1 \registers_reg[688][3]  ( .D(n8161), .E(n115), .CK(clk), .Q(
        \registers[688][3] ) );
  EDFFX1 \registers_reg[688][2]  ( .D(n8110), .E(n115), .CK(clk), .Q(
        \registers[688][2] ) );
  EDFFX1 \registers_reg[688][1]  ( .D(n8054), .E(n115), .CK(clk), .Q(
        \registers[688][1] ) );
  EDFFX1 \registers_reg[688][0]  ( .D(n8025), .E(n115), .CK(clk), .Q(
        \registers[688][0] ) );
  EDFFX1 \registers_reg[684][7]  ( .D(n8379), .E(n111), .CK(clk), .Q(
        \registers[684][7] ) );
  EDFFX1 \registers_reg[684][6]  ( .D(n8321), .E(n111), .CK(clk), .Q(
        \registers[684][6] ) );
  EDFFX1 \registers_reg[684][5]  ( .D(n8263), .E(n111), .CK(clk), .Q(
        \registers[684][5] ) );
  EDFFX1 \registers_reg[684][4]  ( .D(n8205), .E(n111), .CK(clk), .Q(
        \registers[684][4] ) );
  EDFFX1 \registers_reg[684][3]  ( .D(n8161), .E(n111), .CK(clk), .Q(
        \registers[684][3] ) );
  EDFFX1 \registers_reg[684][2]  ( .D(n8108), .E(n111), .CK(clk), .Q(
        \registers[684][2] ) );
  EDFFX1 \registers_reg[684][1]  ( .D(n8052), .E(n111), .CK(clk), .Q(
        \registers[684][1] ) );
  EDFFX1 \registers_reg[684][0]  ( .D(n8039), .E(n111), .CK(clk), .Q(
        \registers[684][0] ) );
  EDFFX1 \registers_reg[680][7]  ( .D(n8377), .E(n107), .CK(clk), .Q(
        \registers[680][7] ) );
  EDFFX1 \registers_reg[680][6]  ( .D(n8319), .E(n107), .CK(clk), .Q(
        \registers[680][6] ) );
  EDFFX1 \registers_reg[680][5]  ( .D(n8261), .E(n107), .CK(clk), .Q(
        \registers[680][5] ) );
  EDFFX1 \registers_reg[680][4]  ( .D(n8203), .E(n107), .CK(clk), .Q(
        \registers[680][4] ) );
  EDFFX1 \registers_reg[680][3]  ( .D(n8161), .E(n107), .CK(clk), .Q(
        \registers[680][3] ) );
  EDFFX1 \registers_reg[680][2]  ( .D(n8106), .E(n107), .CK(clk), .Q(
        \registers[680][2] ) );
  EDFFX1 \registers_reg[680][1]  ( .D(n8050), .E(n107), .CK(clk), .Q(
        \registers[680][1] ) );
  EDFFX1 \registers_reg[680][0]  ( .D(n7994), .E(n107), .CK(clk), .Q(
        \registers[680][0] ) );
  EDFFX1 \registers_reg[676][7]  ( .D(n8377), .E(n298), .CK(clk), .Q(
        \registers[676][7] ) );
  EDFFX1 \registers_reg[676][6]  ( .D(n8319), .E(n298), .CK(clk), .Q(
        \registers[676][6] ) );
  EDFFX1 \registers_reg[676][5]  ( .D(n8261), .E(n298), .CK(clk), .Q(
        \registers[676][5] ) );
  EDFFX1 \registers_reg[676][4]  ( .D(n8203), .E(n298), .CK(clk), .Q(
        \registers[676][4] ) );
  EDFFX1 \registers_reg[676][3]  ( .D(n8753), .E(n298), .CK(clk), .Q(
        \registers[676][3] ) );
  EDFFX1 \registers_reg[676][2]  ( .D(n8107), .E(n298), .CK(clk), .Q(
        \registers[676][2] ) );
  EDFFX1 \registers_reg[676][1]  ( .D(n8051), .E(n298), .CK(clk), .Q(
        \registers[676][1] ) );
  EDFFX1 \registers_reg[676][0]  ( .D(n7994), .E(n298), .CK(clk), .Q(
        \registers[676][0] ) );
  EDFFX1 \registers_reg[672][7]  ( .D(n8377), .E(n1003), .CK(clk), .Q(
        \registers[672][7] ) );
  EDFFX1 \registers_reg[672][6]  ( .D(n8319), .E(n1003), .CK(clk), .Q(
        \registers[672][6] ) );
  EDFFX1 \registers_reg[672][5]  ( .D(n8261), .E(n1003), .CK(clk), .Q(
        \registers[672][5] ) );
  EDFFX1 \registers_reg[672][4]  ( .D(n8203), .E(n1003), .CK(clk), .Q(
        \registers[672][4] ) );
  EDFFX1 \registers_reg[672][3]  ( .D(n8752), .E(n1003), .CK(clk), .Q(
        \registers[672][3] ) );
  EDFFX1 \registers_reg[672][2]  ( .D(n8105), .E(n1003), .CK(clk), .Q(
        \registers[672][2] ) );
  EDFFX1 \registers_reg[672][1]  ( .D(n8049), .E(n1003), .CK(clk), .Q(
        \registers[672][1] ) );
  EDFFX1 \registers_reg[672][0]  ( .D(n7994), .E(n1003), .CK(clk), .Q(
        \registers[672][0] ) );
  EDFFX1 \registers_reg[668][7]  ( .D(n8381), .E(n798), .CK(clk), .Q(
        \registers[668][7] ) );
  EDFFX1 \registers_reg[668][6]  ( .D(n8323), .E(n798), .CK(clk), .Q(
        \registers[668][6] ) );
  EDFFX1 \registers_reg[668][5]  ( .D(n8265), .E(n798), .CK(clk), .Q(
        \registers[668][5] ) );
  EDFFX1 \registers_reg[668][4]  ( .D(n8207), .E(n798), .CK(clk), .Q(
        \registers[668][4] ) );
  EDFFX1 \registers_reg[668][3]  ( .D(n8761), .E(n798), .CK(clk), .Q(
        \registers[668][3] ) );
  EDFFX1 \registers_reg[668][2]  ( .D(n8106), .E(n798), .CK(clk), .Q(
        \registers[668][2] ) );
  EDFFX1 \registers_reg[668][1]  ( .D(n8050), .E(n798), .CK(clk), .Q(
        \registers[668][1] ) );
  EDFFX1 \registers_reg[668][0]  ( .D(n8045), .E(n798), .CK(clk), .Q(
        \registers[668][0] ) );
  EDFFX1 \registers_reg[664][7]  ( .D(n8380), .E(n794), .CK(clk), .Q(
        \registers[664][7] ) );
  EDFFX1 \registers_reg[664][6]  ( .D(n8322), .E(n794), .CK(clk), .Q(
        \registers[664][6] ) );
  EDFFX1 \registers_reg[664][5]  ( .D(n8264), .E(n794), .CK(clk), .Q(
        \registers[664][5] ) );
  EDFFX1 \registers_reg[664][4]  ( .D(n8206), .E(n794), .CK(clk), .Q(
        \registers[664][4] ) );
  EDFFX1 \registers_reg[664][3]  ( .D(n8760), .E(n794), .CK(clk), .Q(
        \registers[664][3] ) );
  EDFFX1 \registers_reg[664][2]  ( .D(n8107), .E(n794), .CK(clk), .Q(
        \registers[664][2] ) );
  EDFFX1 \registers_reg[664][1]  ( .D(n8051), .E(n794), .CK(clk), .Q(
        \registers[664][1] ) );
  EDFFX1 \registers_reg[664][0]  ( .D(n8043), .E(n794), .CK(clk), .Q(
        \registers[664][0] ) );
  EDFFX1 \registers_reg[660][7]  ( .D(n8378), .E(n790), .CK(clk), .Q(
        \registers[660][7] ) );
  EDFFX1 \registers_reg[660][6]  ( .D(n8320), .E(n790), .CK(clk), .Q(
        \registers[660][6] ) );
  EDFFX1 \registers_reg[660][5]  ( .D(n8262), .E(n790), .CK(clk), .Q(
        \registers[660][5] ) );
  EDFFX1 \registers_reg[660][4]  ( .D(n8204), .E(n790), .CK(clk), .Q(
        \registers[660][4] ) );
  EDFFX1 \registers_reg[660][3]  ( .D(n8166), .E(n790), .CK(clk), .Q(
        \registers[660][3] ) );
  EDFFX1 \registers_reg[660][2]  ( .D(n8105), .E(n790), .CK(clk), .Q(
        \registers[660][2] ) );
  EDFFX1 \registers_reg[660][1]  ( .D(n8049), .E(n790), .CK(clk), .Q(
        \registers[660][1] ) );
  EDFFX1 \registers_reg[660][0]  ( .D(data_in[0]), .E(n790), .CK(clk), .Q(
        \registers[660][0] ) );
  EDFFX1 \registers_reg[656][7]  ( .D(n8379), .E(n103), .CK(clk), .Q(
        \registers[656][7] ) );
  EDFFX1 \registers_reg[656][6]  ( .D(n8321), .E(n103), .CK(clk), .Q(
        \registers[656][6] ) );
  EDFFX1 \registers_reg[656][5]  ( .D(n8263), .E(n103), .CK(clk), .Q(
        \registers[656][5] ) );
  EDFFX1 \registers_reg[656][4]  ( .D(n8205), .E(n103), .CK(clk), .Q(
        \registers[656][4] ) );
  EDFFX1 \registers_reg[656][3]  ( .D(n8164), .E(n103), .CK(clk), .Q(
        \registers[656][3] ) );
  EDFFX1 \registers_reg[656][2]  ( .D(n8106), .E(n103), .CK(clk), .Q(
        \registers[656][2] ) );
  EDFFX1 \registers_reg[656][1]  ( .D(n8050), .E(n103), .CK(clk), .Q(
        \registers[656][1] ) );
  EDFFX1 \registers_reg[656][0]  ( .D(n8663), .E(n103), .CK(clk), .Q(
        \registers[656][0] ) );
  EDFFX1 \registers_reg[652][7]  ( .D(n8397), .E(n99), .CK(clk), .Q(
        \registers[652][7] ) );
  EDFFX1 \registers_reg[652][6]  ( .D(n8339), .E(n99), .CK(clk), .Q(
        \registers[652][6] ) );
  EDFFX1 \registers_reg[652][5]  ( .D(n8281), .E(n99), .CK(clk), .Q(
        \registers[652][5] ) );
  EDFFX1 \registers_reg[652][4]  ( .D(n8223), .E(n99), .CK(clk), .Q(
        \registers[652][4] ) );
  EDFFX1 \registers_reg[652][3]  ( .D(n8757), .E(n99), .CK(clk), .Q(
        \registers[652][3] ) );
  EDFFX1 \registers_reg[652][2]  ( .D(n8107), .E(n99), .CK(clk), .Q(
        \registers[652][2] ) );
  EDFFX1 \registers_reg[652][1]  ( .D(n8051), .E(n99), .CK(clk), .Q(
        \registers[652][1] ) );
  EDFFX1 \registers_reg[652][0]  ( .D(n8668), .E(n99), .CK(clk), .Q(
        \registers[652][0] ) );
  EDFFX1 \registers_reg[648][7]  ( .D(n8396), .E(n95), .CK(clk), .Q(
        \registers[648][7] ) );
  EDFFX1 \registers_reg[648][6]  ( .D(n8338), .E(n95), .CK(clk), .Q(
        \registers[648][6] ) );
  EDFFX1 \registers_reg[648][5]  ( .D(n8280), .E(n95), .CK(clk), .Q(
        \registers[648][5] ) );
  EDFFX1 \registers_reg[648][4]  ( .D(n8222), .E(n95), .CK(clk), .Q(
        \registers[648][4] ) );
  EDFFX1 \registers_reg[648][3]  ( .D(n8167), .E(n95), .CK(clk), .Q(
        \registers[648][3] ) );
  EDFFX1 \registers_reg[648][2]  ( .D(n8105), .E(n95), .CK(clk), .Q(
        \registers[648][2] ) );
  EDFFX1 \registers_reg[648][1]  ( .D(n8049), .E(n95), .CK(clk), .Q(
        \registers[648][1] ) );
  EDFFX1 \registers_reg[648][0]  ( .D(n8669), .E(n95), .CK(clk), .Q(
        \registers[648][0] ) );
  EDFFX1 \registers_reg[644][7]  ( .D(n8395), .E(n291), .CK(clk), .Q(
        \registers[644][7] ) );
  EDFFX1 \registers_reg[644][6]  ( .D(n8337), .E(n291), .CK(clk), .Q(
        \registers[644][6] ) );
  EDFFX1 \registers_reg[644][5]  ( .D(n8279), .E(n291), .CK(clk), .Q(
        \registers[644][5] ) );
  EDFFX1 \registers_reg[644][4]  ( .D(n8221), .E(n291), .CK(clk), .Q(
        \registers[644][4] ) );
  EDFFX1 \registers_reg[644][3]  ( .D(n8168), .E(n291), .CK(clk), .Q(
        \registers[644][3] ) );
  EDFFX1 \registers_reg[644][2]  ( .D(n8106), .E(n291), .CK(clk), .Q(
        \registers[644][2] ) );
  EDFFX1 \registers_reg[644][1]  ( .D(n8050), .E(n291), .CK(clk), .Q(
        \registers[644][1] ) );
  EDFFX1 \registers_reg[644][0]  ( .D(n8667), .E(n291), .CK(clk), .Q(
        \registers[644][0] ) );
  EDFFX1 \registers_reg[640][7]  ( .D(n8378), .E(n1002), .CK(clk), .Q(
        \registers[640][7] ) );
  EDFFX1 \registers_reg[640][6]  ( .D(n8320), .E(n1002), .CK(clk), .Q(
        \registers[640][6] ) );
  EDFFX1 \registers_reg[640][5]  ( .D(n8262), .E(n1002), .CK(clk), .Q(
        \registers[640][5] ) );
  EDFFX1 \registers_reg[640][4]  ( .D(n8204), .E(n1002), .CK(clk), .Q(
        \registers[640][4] ) );
  EDFFX1 \registers_reg[640][3]  ( .D(n8751), .E(n1002), .CK(clk), .Q(
        \registers[640][3] ) );
  EDFFX1 \registers_reg[640][2]  ( .D(n8110), .E(n1002), .CK(clk), .Q(
        \registers[640][2] ) );
  EDFFX1 \registers_reg[640][1]  ( .D(n8054), .E(n1002), .CK(clk), .Q(
        \registers[640][1] ) );
  EDFFX1 \registers_reg[640][0]  ( .D(n8009), .E(n1002), .CK(clk), .Q(
        \registers[640][0] ) );
  EDFFX1 \registers_reg[636][7]  ( .D(n8389), .E(n786), .CK(clk), .Q(
        \registers[636][7] ) );
  EDFFX1 \registers_reg[636][6]  ( .D(n8331), .E(n786), .CK(clk), .Q(
        \registers[636][6] ) );
  EDFFX1 \registers_reg[636][5]  ( .D(n8273), .E(n786), .CK(clk), .Q(
        \registers[636][5] ) );
  EDFFX1 \registers_reg[636][4]  ( .D(n8215), .E(n786), .CK(clk), .Q(
        \registers[636][4] ) );
  EDFFX1 \registers_reg[636][3]  ( .D(n8171), .E(n786), .CK(clk), .Q(
        \registers[636][3] ) );
  EDFFX1 \registers_reg[636][2]  ( .D(n8120), .E(n786), .CK(clk), .Q(
        \registers[636][2] ) );
  EDFFX1 \registers_reg[636][1]  ( .D(n8064), .E(n786), .CK(clk), .Q(
        \registers[636][1] ) );
  EDFFX1 \registers_reg[636][0]  ( .D(n8005), .E(n786), .CK(clk), .Q(
        \registers[636][0] ) );
  EDFFX1 \registers_reg[632][7]  ( .D(n8390), .E(n782), .CK(clk), .Q(
        \registers[632][7] ) );
  EDFFX1 \registers_reg[632][6]  ( .D(n8332), .E(n782), .CK(clk), .Q(
        \registers[632][6] ) );
  EDFFX1 \registers_reg[632][5]  ( .D(n8274), .E(n782), .CK(clk), .Q(
        \registers[632][5] ) );
  EDFFX1 \registers_reg[632][4]  ( .D(n8216), .E(n782), .CK(clk), .Q(
        \registers[632][4] ) );
  EDFFX1 \registers_reg[632][3]  ( .D(n8172), .E(n782), .CK(clk), .Q(
        \registers[632][3] ) );
  EDFFX1 \registers_reg[632][2]  ( .D(n8121), .E(n782), .CK(clk), .Q(
        \registers[632][2] ) );
  EDFFX1 \registers_reg[632][1]  ( .D(n8065), .E(n782), .CK(clk), .Q(
        \registers[632][1] ) );
  EDFFX1 \registers_reg[632][0]  ( .D(n8006), .E(n782), .CK(clk), .Q(
        \registers[632][0] ) );
  EDFFX1 \registers_reg[628][7]  ( .D(n8391), .E(n778), .CK(clk), .Q(
        \registers[628][7] ) );
  EDFFX1 \registers_reg[628][6]  ( .D(n8333), .E(n778), .CK(clk), .Q(
        \registers[628][6] ) );
  EDFFX1 \registers_reg[628][5]  ( .D(n8275), .E(n778), .CK(clk), .Q(
        \registers[628][5] ) );
  EDFFX1 \registers_reg[628][4]  ( .D(n8217), .E(n778), .CK(clk), .Q(
        \registers[628][4] ) );
  EDFFX1 \registers_reg[628][3]  ( .D(n8170), .E(n778), .CK(clk), .Q(
        \registers[628][3] ) );
  EDFFX1 \registers_reg[628][2]  ( .D(n8119), .E(n778), .CK(clk), .Q(
        \registers[628][2] ) );
  EDFFX1 \registers_reg[628][1]  ( .D(n8063), .E(n778), .CK(clk), .Q(
        \registers[628][1] ) );
  EDFFX1 \registers_reg[628][0]  ( .D(n8001), .E(n778), .CK(clk), .Q(
        \registers[628][0] ) );
  EDFFX1 \registers_reg[624][7]  ( .D(n8387), .E(n91), .CK(clk), .Q(
        \registers[624][7] ) );
  EDFFX1 \registers_reg[624][6]  ( .D(n8329), .E(n91), .CK(clk), .Q(
        \registers[624][6] ) );
  EDFFX1 \registers_reg[624][5]  ( .D(n8271), .E(n91), .CK(clk), .Q(
        \registers[624][5] ) );
  EDFFX1 \registers_reg[624][4]  ( .D(n8213), .E(n91), .CK(clk), .Q(
        \registers[624][4] ) );
  EDFFX1 \registers_reg[624][3]  ( .D(n8168), .E(n91), .CK(clk), .Q(
        \registers[624][3] ) );
  EDFFX1 \registers_reg[624][2]  ( .D(n8117), .E(n91), .CK(clk), .Q(
        \registers[624][2] ) );
  EDFFX1 \registers_reg[624][1]  ( .D(n8061), .E(n91), .CK(clk), .Q(
        \registers[624][1] ) );
  EDFFX1 \registers_reg[624][0]  ( .D(n8002), .E(n91), .CK(clk), .Q(
        \registers[624][0] ) );
  EDFFX1 \registers_reg[620][7]  ( .D(n8388), .E(n87), .CK(clk), .Q(
        \registers[620][7] ) );
  EDFFX1 \registers_reg[620][6]  ( .D(n8330), .E(n87), .CK(clk), .Q(
        \registers[620][6] ) );
  EDFFX1 \registers_reg[620][5]  ( .D(n8272), .E(n87), .CK(clk), .Q(
        \registers[620][5] ) );
  EDFFX1 \registers_reg[620][4]  ( .D(n8214), .E(n87), .CK(clk), .Q(
        \registers[620][4] ) );
  EDFFX1 \registers_reg[620][3]  ( .D(n8169), .E(n87), .CK(clk), .Q(
        \registers[620][3] ) );
  EDFFX1 \registers_reg[620][2]  ( .D(n8118), .E(n87), .CK(clk), .Q(
        \registers[620][2] ) );
  EDFFX1 \registers_reg[620][1]  ( .D(n8062), .E(n87), .CK(clk), .Q(
        \registers[620][1] ) );
  EDFFX1 \registers_reg[620][0]  ( .D(n8003), .E(n87), .CK(clk), .Q(
        \registers[620][0] ) );
  EDFFX1 \registers_reg[616][7]  ( .D(n8386), .E(n83), .CK(clk), .Q(
        \registers[616][7] ) );
  EDFFX1 \registers_reg[616][6]  ( .D(n8328), .E(n83), .CK(clk), .Q(
        \registers[616][6] ) );
  EDFFX1 \registers_reg[616][5]  ( .D(n8270), .E(n83), .CK(clk), .Q(
        \registers[616][5] ) );
  EDFFX1 \registers_reg[616][4]  ( .D(n8212), .E(n83), .CK(clk), .Q(
        \registers[616][4] ) );
  EDFFX1 \registers_reg[616][3]  ( .D(n8167), .E(n83), .CK(clk), .Q(
        \registers[616][3] ) );
  EDFFX1 \registers_reg[616][2]  ( .D(n8119), .E(n83), .CK(clk), .Q(
        \registers[616][2] ) );
  EDFFX1 \registers_reg[616][1]  ( .D(n8063), .E(n83), .CK(clk), .Q(
        \registers[616][1] ) );
  EDFFX1 \registers_reg[616][0]  ( .D(n8001), .E(n83), .CK(clk), .Q(
        \registers[616][0] ) );
  EDFFX1 \registers_reg[612][7]  ( .D(n8387), .E(n284), .CK(clk), .Q(
        \registers[612][7] ) );
  EDFFX1 \registers_reg[612][6]  ( .D(n8329), .E(n284), .CK(clk), .Q(
        \registers[612][6] ) );
  EDFFX1 \registers_reg[612][5]  ( .D(n8271), .E(n284), .CK(clk), .Q(
        \registers[612][5] ) );
  EDFFX1 \registers_reg[612][4]  ( .D(n8213), .E(n284), .CK(clk), .Q(
        \registers[612][4] ) );
  EDFFX1 \registers_reg[612][3]  ( .D(n8168), .E(n284), .CK(clk), .Q(
        \registers[612][3] ) );
  EDFFX1 \registers_reg[612][2]  ( .D(n8117), .E(n284), .CK(clk), .Q(
        \registers[612][2] ) );
  EDFFX1 \registers_reg[612][1]  ( .D(n8061), .E(n284), .CK(clk), .Q(
        \registers[612][1] ) );
  EDFFX1 \registers_reg[612][0]  ( .D(n8002), .E(n284), .CK(clk), .Q(
        \registers[612][0] ) );
  EDFFX1 \registers_reg[608][7]  ( .D(n8388), .E(n341), .CK(clk), .Q(
        \registers[608][7] ) );
  EDFFX1 \registers_reg[608][6]  ( .D(n8330), .E(n341), .CK(clk), .Q(
        \registers[608][6] ) );
  EDFFX1 \registers_reg[608][5]  ( .D(n8272), .E(n341), .CK(clk), .Q(
        \registers[608][5] ) );
  EDFFX1 \registers_reg[608][4]  ( .D(n8214), .E(n341), .CK(clk), .Q(
        \registers[608][4] ) );
  EDFFX1 \registers_reg[608][3]  ( .D(n8169), .E(n341), .CK(clk), .Q(
        \registers[608][3] ) );
  EDFFX1 \registers_reg[608][2]  ( .D(n8118), .E(n341), .CK(clk), .Q(
        \registers[608][2] ) );
  EDFFX1 \registers_reg[608][1]  ( .D(n8062), .E(n341), .CK(clk), .Q(
        \registers[608][1] ) );
  EDFFX1 \registers_reg[608][0]  ( .D(n8003), .E(n341), .CK(clk), .Q(
        \registers[608][0] ) );
  EDFFX1 \registers_reg[604][7]  ( .D(n8386), .E(n774), .CK(clk), .Q(
        \registers[604][7] ) );
  EDFFX1 \registers_reg[604][6]  ( .D(n8328), .E(n774), .CK(clk), .Q(
        \registers[604][6] ) );
  EDFFX1 \registers_reg[604][5]  ( .D(n8270), .E(n774), .CK(clk), .Q(
        \registers[604][5] ) );
  EDFFX1 \registers_reg[604][4]  ( .D(n8212), .E(n774), .CK(clk), .Q(
        \registers[604][4] ) );
  EDFFX1 \registers_reg[604][3]  ( .D(n8167), .E(n774), .CK(clk), .Q(
        \registers[604][3] ) );
  EDFFX1 \registers_reg[604][2]  ( .D(n8119), .E(n774), .CK(clk), .Q(
        \registers[604][2] ) );
  EDFFX1 \registers_reg[604][1]  ( .D(n8063), .E(n774), .CK(clk), .Q(
        \registers[604][1] ) );
  EDFFX1 \registers_reg[604][0]  ( .D(n8001), .E(n774), .CK(clk), .Q(
        \registers[604][0] ) );
  EDFFX1 \registers_reg[600][7]  ( .D(n8387), .E(n770), .CK(clk), .Q(
        \registers[600][7] ) );
  EDFFX1 \registers_reg[600][6]  ( .D(n8329), .E(n770), .CK(clk), .Q(
        \registers[600][6] ) );
  EDFFX1 \registers_reg[600][5]  ( .D(n8271), .E(n770), .CK(clk), .Q(
        \registers[600][5] ) );
  EDFFX1 \registers_reg[600][4]  ( .D(n8213), .E(n770), .CK(clk), .Q(
        \registers[600][4] ) );
  EDFFX1 \registers_reg[600][3]  ( .D(n8168), .E(n770), .CK(clk), .Q(
        \registers[600][3] ) );
  EDFFX1 \registers_reg[600][2]  ( .D(n8117), .E(n770), .CK(clk), .Q(
        \registers[600][2] ) );
  EDFFX1 \registers_reg[600][1]  ( .D(n8061), .E(n770), .CK(clk), .Q(
        \registers[600][1] ) );
  EDFFX1 \registers_reg[600][0]  ( .D(n8002), .E(n770), .CK(clk), .Q(
        \registers[600][0] ) );
  EDFFX1 \registers_reg[596][7]  ( .D(n8388), .E(n766), .CK(clk), .Q(
        \registers[596][7] ) );
  EDFFX1 \registers_reg[596][6]  ( .D(n8330), .E(n766), .CK(clk), .Q(
        \registers[596][6] ) );
  EDFFX1 \registers_reg[596][5]  ( .D(n8272), .E(n766), .CK(clk), .Q(
        \registers[596][5] ) );
  EDFFX1 \registers_reg[596][4]  ( .D(n8214), .E(n766), .CK(clk), .Q(
        \registers[596][4] ) );
  EDFFX1 \registers_reg[596][3]  ( .D(n8169), .E(n766), .CK(clk), .Q(
        \registers[596][3] ) );
  EDFFX1 \registers_reg[596][2]  ( .D(n8118), .E(n766), .CK(clk), .Q(
        \registers[596][2] ) );
  EDFFX1 \registers_reg[596][1]  ( .D(n8062), .E(n766), .CK(clk), .Q(
        \registers[596][1] ) );
  EDFFX1 \registers_reg[596][0]  ( .D(n8003), .E(n766), .CK(clk), .Q(
        \registers[596][0] ) );
  EDFFX1 \registers_reg[592][7]  ( .D(n8386), .E(n79), .CK(clk), .Q(
        \registers[592][7] ) );
  EDFFX1 \registers_reg[592][6]  ( .D(n8328), .E(n79), .CK(clk), .Q(
        \registers[592][6] ) );
  EDFFX1 \registers_reg[592][5]  ( .D(n8270), .E(n79), .CK(clk), .Q(
        \registers[592][5] ) );
  EDFFX1 \registers_reg[592][4]  ( .D(n8212), .E(n79), .CK(clk), .Q(
        \registers[592][4] ) );
  EDFFX1 \registers_reg[592][3]  ( .D(n8167), .E(n79), .CK(clk), .Q(
        \registers[592][3] ) );
  EDFFX1 \registers_reg[592][2]  ( .D(n8119), .E(n79), .CK(clk), .Q(
        \registers[592][2] ) );
  EDFFX1 \registers_reg[592][1]  ( .D(n8063), .E(n79), .CK(clk), .Q(
        \registers[592][1] ) );
  EDFFX1 \registers_reg[592][0]  ( .D(n8001), .E(n79), .CK(clk), .Q(
        \registers[592][0] ) );
  EDFFX1 \registers_reg[588][7]  ( .D(n8387), .E(n75), .CK(clk), .Q(
        \registers[588][7] ) );
  EDFFX1 \registers_reg[588][6]  ( .D(n8329), .E(n75), .CK(clk), .Q(
        \registers[588][6] ) );
  EDFFX1 \registers_reg[588][5]  ( .D(n8271), .E(n75), .CK(clk), .Q(
        \registers[588][5] ) );
  EDFFX1 \registers_reg[588][4]  ( .D(n8213), .E(n75), .CK(clk), .Q(
        \registers[588][4] ) );
  EDFFX1 \registers_reg[588][3]  ( .D(n8168), .E(n75), .CK(clk), .Q(
        \registers[588][3] ) );
  EDFFX1 \registers_reg[588][2]  ( .D(n8117), .E(n75), .CK(clk), .Q(
        \registers[588][2] ) );
  EDFFX1 \registers_reg[588][1]  ( .D(n8061), .E(n75), .CK(clk), .Q(
        \registers[588][1] ) );
  EDFFX1 \registers_reg[588][0]  ( .D(n8002), .E(n75), .CK(clk), .Q(
        \registers[588][0] ) );
  EDFFX1 \registers_reg[584][7]  ( .D(n8388), .E(n71), .CK(clk), .Q(
        \registers[584][7] ) );
  EDFFX1 \registers_reg[584][6]  ( .D(n8330), .E(n71), .CK(clk), .Q(
        \registers[584][6] ) );
  EDFFX1 \registers_reg[584][5]  ( .D(n8272), .E(n71), .CK(clk), .Q(
        \registers[584][5] ) );
  EDFFX1 \registers_reg[584][4]  ( .D(n8214), .E(n71), .CK(clk), .Q(
        \registers[584][4] ) );
  EDFFX1 \registers_reg[584][3]  ( .D(n8169), .E(n71), .CK(clk), .Q(
        \registers[584][3] ) );
  EDFFX1 \registers_reg[584][2]  ( .D(n8118), .E(n71), .CK(clk), .Q(
        \registers[584][2] ) );
  EDFFX1 \registers_reg[584][1]  ( .D(n8062), .E(n71), .CK(clk), .Q(
        \registers[584][1] ) );
  EDFFX1 \registers_reg[584][0]  ( .D(n8003), .E(n71), .CK(clk), .Q(
        \registers[584][0] ) );
  EDFFX1 \registers_reg[580][7]  ( .D(n8386), .E(n277), .CK(clk), .Q(
        \registers[580][7] ) );
  EDFFX1 \registers_reg[580][6]  ( .D(n8328), .E(n277), .CK(clk), .Q(
        \registers[580][6] ) );
  EDFFX1 \registers_reg[580][5]  ( .D(n8270), .E(n277), .CK(clk), .Q(
        \registers[580][5] ) );
  EDFFX1 \registers_reg[580][4]  ( .D(n8212), .E(n277), .CK(clk), .Q(
        \registers[580][4] ) );
  EDFFX1 \registers_reg[580][3]  ( .D(n8167), .E(n277), .CK(clk), .Q(
        \registers[580][3] ) );
  EDFFX1 \registers_reg[580][2]  ( .D(n8119), .E(n277), .CK(clk), .Q(
        \registers[580][2] ) );
  EDFFX1 \registers_reg[580][1]  ( .D(n8063), .E(n277), .CK(clk), .Q(
        \registers[580][1] ) );
  EDFFX1 \registers_reg[580][0]  ( .D(n8001), .E(n277), .CK(clk), .Q(
        \registers[580][0] ) );
  EDFFX1 \registers_reg[576][7]  ( .D(n8384), .E(n340), .CK(clk), .Q(
        \registers[576][7] ) );
  EDFFX1 \registers_reg[576][6]  ( .D(n8326), .E(n340), .CK(clk), .Q(
        \registers[576][6] ) );
  EDFFX1 \registers_reg[576][5]  ( .D(n8268), .E(n340), .CK(clk), .Q(
        \registers[576][5] ) );
  EDFFX1 \registers_reg[576][4]  ( .D(n8210), .E(n340), .CK(clk), .Q(
        \registers[576][4] ) );
  EDFFX1 \registers_reg[576][3]  ( .D(n8169), .E(n340), .CK(clk), .Q(
        \registers[576][3] ) );
  EDFFX1 \registers_reg[576][2]  ( .D(n8115), .E(n340), .CK(clk), .Q(
        \registers[576][2] ) );
  EDFFX1 \registers_reg[576][1]  ( .D(n8059), .E(n340), .CK(clk), .Q(
        \registers[576][1] ) );
  EDFFX1 \registers_reg[576][0]  ( .D(n7999), .E(n340), .CK(clk), .Q(
        \registers[576][0] ) );
  EDFFX1 \registers_reg[572][7]  ( .D(n8430), .E(n762), .CK(clk), .Q(
        \registers[572][7] ) );
  EDFFX1 \registers_reg[572][6]  ( .D(n8372), .E(n762), .CK(clk), .Q(
        \registers[572][6] ) );
  EDFFX1 \registers_reg[572][5]  ( .D(n8314), .E(n762), .CK(clk), .Q(
        \registers[572][5] ) );
  EDFFX1 \registers_reg[572][4]  ( .D(n8256), .E(n762), .CK(clk), .Q(
        \registers[572][4] ) );
  EDFFX1 \registers_reg[572][3]  ( .D(n8167), .E(n762), .CK(clk), .Q(
        \registers[572][3] ) );
  EDFFX1 \registers_reg[572][2]  ( .D(n8116), .E(n762), .CK(clk), .Q(
        \registers[572][2] ) );
  EDFFX1 \registers_reg[572][1]  ( .D(n8060), .E(n762), .CK(clk), .Q(
        \registers[572][1] ) );
  EDFFX1 \registers_reg[572][0]  ( .D(n7998), .E(n762), .CK(clk), .Q(
        \registers[572][0] ) );
  EDFFX1 \registers_reg[568][7]  ( .D(n8385), .E(n758), .CK(clk), .Q(
        \registers[568][7] ) );
  EDFFX1 \registers_reg[568][6]  ( .D(n8327), .E(n758), .CK(clk), .Q(
        \registers[568][6] ) );
  EDFFX1 \registers_reg[568][5]  ( .D(n8269), .E(n758), .CK(clk), .Q(
        \registers[568][5] ) );
  EDFFX1 \registers_reg[568][4]  ( .D(n8211), .E(n758), .CK(clk), .Q(
        \registers[568][4] ) );
  EDFFX1 \registers_reg[568][3]  ( .D(n8168), .E(n758), .CK(clk), .Q(
        \registers[568][3] ) );
  EDFFX1 \registers_reg[568][2]  ( .D(n8114), .E(n758), .CK(clk), .Q(
        \registers[568][2] ) );
  EDFFX1 \registers_reg[568][1]  ( .D(n8058), .E(n758), .CK(clk), .Q(
        \registers[568][1] ) );
  EDFFX1 \registers_reg[568][0]  ( .D(n7999), .E(n758), .CK(clk), .Q(
        \registers[568][0] ) );
  EDFFX1 \registers_reg[564][7]  ( .D(n8384), .E(n754), .CK(clk), .Q(
        \registers[564][7] ) );
  EDFFX1 \registers_reg[564][6]  ( .D(n8326), .E(n754), .CK(clk), .Q(
        \registers[564][6] ) );
  EDFFX1 \registers_reg[564][5]  ( .D(n8268), .E(n754), .CK(clk), .Q(
        \registers[564][5] ) );
  EDFFX1 \registers_reg[564][4]  ( .D(n8210), .E(n754), .CK(clk), .Q(
        \registers[564][4] ) );
  EDFFX1 \registers_reg[564][3]  ( .D(n8169), .E(n754), .CK(clk), .Q(
        \registers[564][3] ) );
  EDFFX1 \registers_reg[564][2]  ( .D(n8115), .E(n754), .CK(clk), .Q(
        \registers[564][2] ) );
  EDFFX1 \registers_reg[564][1]  ( .D(n8059), .E(n754), .CK(clk), .Q(
        \registers[564][1] ) );
  EDFFX1 \registers_reg[564][0]  ( .D(n8000), .E(n754), .CK(clk), .Q(
        \registers[564][0] ) );
  EDFFX1 \registers_reg[560][7]  ( .D(n8431), .E(n67), .CK(clk), .Q(
        \registers[560][7] ) );
  EDFFX1 \registers_reg[560][6]  ( .D(n8373), .E(n67), .CK(clk), .Q(
        \registers[560][6] ) );
  EDFFX1 \registers_reg[560][5]  ( .D(n8315), .E(n67), .CK(clk), .Q(
        \registers[560][5] ) );
  EDFFX1 \registers_reg[560][4]  ( .D(n8257), .E(n67), .CK(clk), .Q(
        \registers[560][4] ) );
  EDFFX1 \registers_reg[560][3]  ( .D(n8164), .E(n67), .CK(clk), .Q(
        \registers[560][3] ) );
  EDFFX1 \registers_reg[560][2]  ( .D(n8116), .E(n67), .CK(clk), .Q(
        \registers[560][2] ) );
  EDFFX1 \registers_reg[560][1]  ( .D(n8060), .E(n67), .CK(clk), .Q(
        \registers[560][1] ) );
  EDFFX1 \registers_reg[560][0]  ( .D(n7998), .E(n67), .CK(clk), .Q(
        \registers[560][0] ) );
  EDFFX1 \registers_reg[556][7]  ( .D(n8385), .E(n63), .CK(clk), .Q(
        \registers[556][7] ) );
  EDFFX1 \registers_reg[556][6]  ( .D(n8327), .E(n63), .CK(clk), .Q(
        \registers[556][6] ) );
  EDFFX1 \registers_reg[556][5]  ( .D(n8269), .E(n63), .CK(clk), .Q(
        \registers[556][5] ) );
  EDFFX1 \registers_reg[556][4]  ( .D(n8211), .E(n63), .CK(clk), .Q(
        \registers[556][4] ) );
  EDFFX1 \registers_reg[556][3]  ( .D(n8165), .E(n63), .CK(clk), .Q(
        \registers[556][3] ) );
  EDFFX1 \registers_reg[556][2]  ( .D(n8114), .E(n63), .CK(clk), .Q(
        \registers[556][2] ) );
  EDFFX1 \registers_reg[556][1]  ( .D(n8058), .E(n63), .CK(clk), .Q(
        \registers[556][1] ) );
  EDFFX1 \registers_reg[556][0]  ( .D(n7999), .E(n63), .CK(clk), .Q(
        \registers[556][0] ) );
  EDFFX1 \registers_reg[552][7]  ( .D(n8384), .E(n59), .CK(clk), .Q(
        \registers[552][7] ) );
  EDFFX1 \registers_reg[552][6]  ( .D(n8326), .E(n59), .CK(clk), .Q(
        \registers[552][6] ) );
  EDFFX1 \registers_reg[552][5]  ( .D(n8268), .E(n59), .CK(clk), .Q(
        \registers[552][5] ) );
  EDFFX1 \registers_reg[552][4]  ( .D(n8210), .E(n59), .CK(clk), .Q(
        \registers[552][4] ) );
  EDFFX1 \registers_reg[552][3]  ( .D(n8166), .E(n59), .CK(clk), .Q(
        \registers[552][3] ) );
  EDFFX1 \registers_reg[552][2]  ( .D(n8115), .E(n59), .CK(clk), .Q(
        \registers[552][2] ) );
  EDFFX1 \registers_reg[552][1]  ( .D(n8059), .E(n59), .CK(clk), .Q(
        \registers[552][1] ) );
  EDFFX1 \registers_reg[552][0]  ( .D(n8000), .E(n59), .CK(clk), .Q(
        \registers[552][0] ) );
  EDFFX1 \registers_reg[548][7]  ( .D(n8383), .E(n270), .CK(clk), .Q(
        \registers[548][7] ) );
  EDFFX1 \registers_reg[548][6]  ( .D(n8325), .E(n270), .CK(clk), .Q(
        \registers[548][6] ) );
  EDFFX1 \registers_reg[548][5]  ( .D(n8267), .E(n270), .CK(clk), .Q(
        \registers[548][5] ) );
  EDFFX1 \registers_reg[548][4]  ( .D(n8209), .E(n270), .CK(clk), .Q(
        \registers[548][4] ) );
  EDFFX1 \registers_reg[548][3]  ( .D(n8164), .E(n270), .CK(clk), .Q(
        \registers[548][3] ) );
  EDFFX1 \registers_reg[548][2]  ( .D(n8116), .E(n270), .CK(clk), .Q(
        \registers[548][2] ) );
  EDFFX1 \registers_reg[548][1]  ( .D(n8060), .E(n270), .CK(clk), .Q(
        \registers[548][1] ) );
  EDFFX1 \registers_reg[548][0]  ( .D(n7998), .E(n270), .CK(clk), .Q(
        \registers[548][0] ) );
  EDFFX1 \registers_reg[544][7]  ( .D(n8385), .E(n339), .CK(clk), .Q(
        \registers[544][7] ) );
  EDFFX1 \registers_reg[544][6]  ( .D(n8327), .E(n339), .CK(clk), .Q(
        \registers[544][6] ) );
  EDFFX1 \registers_reg[544][5]  ( .D(n8269), .E(n339), .CK(clk), .Q(
        \registers[544][5] ) );
  EDFFX1 \registers_reg[544][4]  ( .D(n8211), .E(n339), .CK(clk), .Q(
        \registers[544][4] ) );
  EDFFX1 \registers_reg[544][3]  ( .D(n8165), .E(n339), .CK(clk), .Q(
        \registers[544][3] ) );
  EDFFX1 \registers_reg[544][2]  ( .D(n8114), .E(n339), .CK(clk), .Q(
        \registers[544][2] ) );
  EDFFX1 \registers_reg[544][1]  ( .D(n8058), .E(n339), .CK(clk), .Q(
        \registers[544][1] ) );
  EDFFX1 \registers_reg[544][0]  ( .D(n7999), .E(n339), .CK(clk), .Q(
        \registers[544][0] ) );
  EDFFX1 \registers_reg[540][7]  ( .D(n8384), .E(n750), .CK(clk), .Q(
        \registers[540][7] ) );
  EDFFX1 \registers_reg[540][6]  ( .D(n8326), .E(n750), .CK(clk), .Q(
        \registers[540][6] ) );
  EDFFX1 \registers_reg[540][5]  ( .D(n8268), .E(n750), .CK(clk), .Q(
        \registers[540][5] ) );
  EDFFX1 \registers_reg[540][4]  ( .D(n8210), .E(n750), .CK(clk), .Q(
        \registers[540][4] ) );
  EDFFX1 \registers_reg[540][3]  ( .D(n8166), .E(n750), .CK(clk), .Q(
        \registers[540][3] ) );
  EDFFX1 \registers_reg[540][2]  ( .D(n8115), .E(n750), .CK(clk), .Q(
        \registers[540][2] ) );
  EDFFX1 \registers_reg[540][1]  ( .D(n8059), .E(n750), .CK(clk), .Q(
        \registers[540][1] ) );
  EDFFX1 \registers_reg[540][0]  ( .D(n8000), .E(n750), .CK(clk), .Q(
        \registers[540][0] ) );
  EDFFX1 \registers_reg[536][7]  ( .D(n8406), .E(n746), .CK(clk), .Q(
        \registers[536][7] ) );
  EDFFX1 \registers_reg[536][6]  ( .D(n8348), .E(n746), .CK(clk), .Q(
        \registers[536][6] ) );
  EDFFX1 \registers_reg[536][5]  ( .D(n8290), .E(n746), .CK(clk), .Q(
        \registers[536][5] ) );
  EDFFX1 \registers_reg[536][4]  ( .D(n8232), .E(n746), .CK(clk), .Q(
        \registers[536][4] ) );
  EDFFX1 \registers_reg[536][3]  ( .D(n8164), .E(n746), .CK(clk), .Q(
        \registers[536][3] ) );
  EDFFX1 \registers_reg[536][2]  ( .D(n8116), .E(n746), .CK(clk), .Q(
        \registers[536][2] ) );
  EDFFX1 \registers_reg[536][1]  ( .D(n8060), .E(n746), .CK(clk), .Q(
        \registers[536][1] ) );
  EDFFX1 \registers_reg[536][0]  ( .D(n7998), .E(n746), .CK(clk), .Q(
        \registers[536][0] ) );
  EDFFX1 \registers_reg[532][7]  ( .D(n8385), .E(n742), .CK(clk), .Q(
        \registers[532][7] ) );
  EDFFX1 \registers_reg[532][6]  ( .D(n8327), .E(n742), .CK(clk), .Q(
        \registers[532][6] ) );
  EDFFX1 \registers_reg[532][5]  ( .D(n8269), .E(n742), .CK(clk), .Q(
        \registers[532][5] ) );
  EDFFX1 \registers_reg[532][4]  ( .D(n8211), .E(n742), .CK(clk), .Q(
        \registers[532][4] ) );
  EDFFX1 \registers_reg[532][3]  ( .D(n8165), .E(n742), .CK(clk), .Q(
        \registers[532][3] ) );
  EDFFX1 \registers_reg[532][2]  ( .D(n8114), .E(n742), .CK(clk), .Q(
        \registers[532][2] ) );
  EDFFX1 \registers_reg[532][1]  ( .D(n8058), .E(n742), .CK(clk), .Q(
        \registers[532][1] ) );
  EDFFX1 \registers_reg[532][0]  ( .D(n7999), .E(n742), .CK(clk), .Q(
        \registers[532][0] ) );
  EDFFX1 \registers_reg[528][7]  ( .D(n8384), .E(n55), .CK(clk), .Q(
        \registers[528][7] ) );
  EDFFX1 \registers_reg[528][6]  ( .D(n8326), .E(n55), .CK(clk), .Q(
        \registers[528][6] ) );
  EDFFX1 \registers_reg[528][5]  ( .D(n8268), .E(n55), .CK(clk), .Q(
        \registers[528][5] ) );
  EDFFX1 \registers_reg[528][4]  ( .D(n8210), .E(n55), .CK(clk), .Q(
        \registers[528][4] ) );
  EDFFX1 \registers_reg[528][3]  ( .D(n8166), .E(n55), .CK(clk), .Q(
        \registers[528][3] ) );
  EDFFX1 \registers_reg[528][2]  ( .D(n8112), .E(n55), .CK(clk), .Q(
        \registers[528][2] ) );
  EDFFX1 \registers_reg[528][1]  ( .D(n8056), .E(n55), .CK(clk), .Q(
        \registers[528][1] ) );
  EDFFX1 \registers_reg[528][0]  ( .D(n8000), .E(n55), .CK(clk), .Q(
        \registers[528][0] ) );
  EDFFX1 \registers_reg[524][7]  ( .D(n8383), .E(n50), .CK(clk), .Q(
        \registers[524][7] ) );
  EDFFX1 \registers_reg[524][6]  ( .D(n8325), .E(n50), .CK(clk), .Q(
        \registers[524][6] ) );
  EDFFX1 \registers_reg[524][5]  ( .D(n8267), .E(n50), .CK(clk), .Q(
        \registers[524][5] ) );
  EDFFX1 \registers_reg[524][4]  ( .D(n8209), .E(n50), .CK(clk), .Q(
        \registers[524][4] ) );
  EDFFX1 \registers_reg[524][3]  ( .D(n8164), .E(n50), .CK(clk), .Q(
        \registers[524][3] ) );
  EDFFX1 \registers_reg[524][2]  ( .D(n8113), .E(n50), .CK(clk), .Q(
        \registers[524][2] ) );
  EDFFX1 \registers_reg[524][1]  ( .D(n8057), .E(n50), .CK(clk), .Q(
        \registers[524][1] ) );
  EDFFX1 \registers_reg[524][0]  ( .D(n7996), .E(n50), .CK(clk), .Q(
        \registers[524][0] ) );
  EDFFX1 \registers_reg[520][7]  ( .D(n8381), .E(n46), .CK(clk), .Q(
        \registers[520][7] ) );
  EDFFX1 \registers_reg[520][6]  ( .D(n8323), .E(n46), .CK(clk), .Q(
        \registers[520][6] ) );
  EDFFX1 \registers_reg[520][5]  ( .D(n8265), .E(n46), .CK(clk), .Q(
        \registers[520][5] ) );
  EDFFX1 \registers_reg[520][4]  ( .D(n8207), .E(n46), .CK(clk), .Q(
        \registers[520][4] ) );
  EDFFX1 \registers_reg[520][3]  ( .D(n8165), .E(n46), .CK(clk), .Q(
        \registers[520][3] ) );
  EDFFX1 \registers_reg[520][2]  ( .D(n8111), .E(n46), .CK(clk), .Q(
        \registers[520][2] ) );
  EDFFX1 \registers_reg[520][1]  ( .D(n8055), .E(n46), .CK(clk), .Q(
        \registers[520][1] ) );
  EDFFX1 \registers_reg[520][0]  ( .D(n7997), .E(n46), .CK(clk), .Q(
        \registers[520][0] ) );
  EDFFX1 \registers_reg[516][7]  ( .D(n8382), .E(n263), .CK(clk), .Q(
        \registers[516][7] ) );
  EDFFX1 \registers_reg[516][6]  ( .D(n8324), .E(n263), .CK(clk), .Q(
        \registers[516][6] ) );
  EDFFX1 \registers_reg[516][5]  ( .D(n8266), .E(n263), .CK(clk), .Q(
        \registers[516][5] ) );
  EDFFX1 \registers_reg[516][4]  ( .D(n8208), .E(n263), .CK(clk), .Q(
        \registers[516][4] ) );
  EDFFX1 \registers_reg[516][3]  ( .D(n8166), .E(n263), .CK(clk), .Q(
        \registers[516][3] ) );
  EDFFX1 \registers_reg[516][2]  ( .D(n8112), .E(n263), .CK(clk), .Q(
        \registers[516][2] ) );
  EDFFX1 \registers_reg[516][1]  ( .D(n8056), .E(n263), .CK(clk), .Q(
        \registers[516][1] ) );
  EDFFX1 \registers_reg[516][0]  ( .D(n8671), .E(n263), .CK(clk), .Q(
        \registers[516][0] ) );
  EDFFX1 \registers_reg[512][7]  ( .D(n8391), .E(n338), .CK(clk), .Q(
        \registers[512][7] ) );
  EDFFX1 \registers_reg[512][6]  ( .D(n8333), .E(n338), .CK(clk), .Q(
        \registers[512][6] ) );
  EDFFX1 \registers_reg[512][5]  ( .D(n8275), .E(n338), .CK(clk), .Q(
        \registers[512][5] ) );
  EDFFX1 \registers_reg[512][4]  ( .D(n8217), .E(n338), .CK(clk), .Q(
        \registers[512][4] ) );
  EDFFX1 \registers_reg[512][3]  ( .D(n8170), .E(n338), .CK(clk), .Q(
        \registers[512][3] ) );
  EDFFX1 \registers_reg[512][2]  ( .D(n8122), .E(n338), .CK(clk), .Q(
        \registers[512][2] ) );
  EDFFX1 \registers_reg[512][1]  ( .D(n8066), .E(n338), .CK(clk), .Q(
        \registers[512][1] ) );
  EDFFX1 \registers_reg[512][0]  ( .D(n8000), .E(n338), .CK(clk), .Q(
        \registers[512][0] ) );
  EDFFX1 \registers_reg[508][7]  ( .D(n8428), .E(n738), .CK(clk), .Q(
        \registers[508][7] ) );
  EDFFX1 \registers_reg[508][6]  ( .D(n8370), .E(n738), .CK(clk), .Q(
        \registers[508][6] ) );
  EDFFX1 \registers_reg[508][5]  ( .D(n8312), .E(n738), .CK(clk), .Q(
        \registers[508][5] ) );
  EDFFX1 \registers_reg[508][4]  ( .D(n8254), .E(n738), .CK(clk), .Q(
        \registers[508][4] ) );
  EDFFX1 \registers_reg[508][3]  ( .D(n8202), .E(n738), .CK(clk), .Q(
        \registers[508][3] ) );
  EDFFX1 \registers_reg[508][2]  ( .D(n8156), .E(n738), .CK(clk), .Q(
        \registers[508][2] ) );
  EDFFX1 \registers_reg[508][1]  ( .D(n8100), .E(n738), .CK(clk), .Q(
        \registers[508][1] ) );
  EDFFX1 \registers_reg[508][0]  ( .D(n8040), .E(n738), .CK(clk), .Q(
        \registers[508][0] ) );
  EDFFX1 \registers_reg[504][7]  ( .D(n8427), .E(n734), .CK(clk), .Q(
        \registers[504][7] ) );
  EDFFX1 \registers_reg[504][6]  ( .D(n8369), .E(n734), .CK(clk), .Q(
        \registers[504][6] ) );
  EDFFX1 \registers_reg[504][5]  ( .D(n8311), .E(n734), .CK(clk), .Q(
        \registers[504][5] ) );
  EDFFX1 \registers_reg[504][4]  ( .D(n8253), .E(n734), .CK(clk), .Q(
        \registers[504][4] ) );
  EDFFX1 \registers_reg[504][3]  ( .D(n8200), .E(n734), .CK(clk), .Q(
        \registers[504][3] ) );
  EDFFX1 \registers_reg[504][2]  ( .D(n8157), .E(n734), .CK(clk), .Q(
        \registers[504][2] ) );
  EDFFX1 \registers_reg[504][1]  ( .D(n8101), .E(n734), .CK(clk), .Q(
        \registers[504][1] ) );
  EDFFX1 \registers_reg[504][0]  ( .D(n8041), .E(n734), .CK(clk), .Q(
        \registers[504][0] ) );
  EDFFX1 \registers_reg[500][7]  ( .D(n8425), .E(n730), .CK(clk), .Q(
        \registers[500][7] ) );
  EDFFX1 \registers_reg[500][6]  ( .D(n8367), .E(n730), .CK(clk), .Q(
        \registers[500][6] ) );
  EDFFX1 \registers_reg[500][5]  ( .D(n8309), .E(n730), .CK(clk), .Q(
        \registers[500][5] ) );
  EDFFX1 \registers_reg[500][4]  ( .D(n8251), .E(n730), .CK(clk), .Q(
        \registers[500][4] ) );
  EDFFX1 \registers_reg[500][3]  ( .D(n8201), .E(n730), .CK(clk), .Q(
        \registers[500][3] ) );
  EDFFX1 \registers_reg[500][2]  ( .D(n8155), .E(n730), .CK(clk), .Q(
        \registers[500][2] ) );
  EDFFX1 \registers_reg[500][1]  ( .D(n8099), .E(n730), .CK(clk), .Q(
        \registers[500][1] ) );
  EDFFX1 \registers_reg[500][0]  ( .D(n8042), .E(n730), .CK(clk), .Q(
        \registers[500][0] ) );
  EDFFX1 \registers_reg[496][7]  ( .D(n8426), .E(n42), .CK(clk), .Q(
        \registers[496][7] ) );
  EDFFX1 \registers_reg[496][6]  ( .D(n8368), .E(n42), .CK(clk), .Q(
        \registers[496][6] ) );
  EDFFX1 \registers_reg[496][5]  ( .D(n8310), .E(n42), .CK(clk), .Q(
        \registers[496][5] ) );
  EDFFX1 \registers_reg[496][4]  ( .D(n8252), .E(n42), .CK(clk), .Q(
        \registers[496][4] ) );
  EDFFX1 \registers_reg[496][3]  ( .D(n8202), .E(n42), .CK(clk), .Q(
        \registers[496][3] ) );
  EDFFX1 \registers_reg[496][2]  ( .D(n8156), .E(n42), .CK(clk), .Q(
        \registers[496][2] ) );
  EDFFX1 \registers_reg[496][1]  ( .D(n8100), .E(n42), .CK(clk), .Q(
        \registers[496][1] ) );
  EDFFX1 \registers_reg[496][0]  ( .D(n8040), .E(n42), .CK(clk), .Q(
        \registers[496][0] ) );
  EDFFX1 \registers_reg[492][7]  ( .D(n8427), .E(n38), .CK(clk), .Q(
        \registers[492][7] ) );
  EDFFX1 \registers_reg[492][6]  ( .D(n8369), .E(n38), .CK(clk), .Q(
        \registers[492][6] ) );
  EDFFX1 \registers_reg[492][5]  ( .D(n8311), .E(n38), .CK(clk), .Q(
        \registers[492][5] ) );
  EDFFX1 \registers_reg[492][4]  ( .D(n8253), .E(n38), .CK(clk), .Q(
        \registers[492][4] ) );
  EDFFX1 \registers_reg[492][3]  ( .D(n8200), .E(n38), .CK(clk), .Q(
        \registers[492][3] ) );
  EDFFX1 \registers_reg[492][2]  ( .D(n8157), .E(n38), .CK(clk), .Q(
        \registers[492][2] ) );
  EDFFX1 \registers_reg[492][1]  ( .D(n8101), .E(n38), .CK(clk), .Q(
        \registers[492][1] ) );
  EDFFX1 \registers_reg[492][0]  ( .D(n8041), .E(n38), .CK(clk), .Q(
        \registers[492][0] ) );
  EDFFX1 \registers_reg[488][7]  ( .D(n8425), .E(n34), .CK(clk), .Q(
        \registers[488][7] ) );
  EDFFX1 \registers_reg[488][6]  ( .D(n8367), .E(n34), .CK(clk), .Q(
        \registers[488][6] ) );
  EDFFX1 \registers_reg[488][5]  ( .D(n8309), .E(n34), .CK(clk), .Q(
        \registers[488][5] ) );
  EDFFX1 \registers_reg[488][4]  ( .D(n8251), .E(n34), .CK(clk), .Q(
        \registers[488][4] ) );
  EDFFX1 \registers_reg[488][3]  ( .D(n8201), .E(n34), .CK(clk), .Q(
        \registers[488][3] ) );
  EDFFX1 \registers_reg[488][2]  ( .D(n8155), .E(n34), .CK(clk), .Q(
        \registers[488][2] ) );
  EDFFX1 \registers_reg[488][1]  ( .D(n8099), .E(n34), .CK(clk), .Q(
        \registers[488][1] ) );
  EDFFX1 \registers_reg[488][0]  ( .D(n8042), .E(n34), .CK(clk), .Q(
        \registers[488][0] ) );
  EDFFX1 \registers_reg[484][7]  ( .D(n8426), .E(n256), .CK(clk), .Q(
        \registers[484][7] ) );
  EDFFX1 \registers_reg[484][6]  ( .D(n8368), .E(n256), .CK(clk), .Q(
        \registers[484][6] ) );
  EDFFX1 \registers_reg[484][5]  ( .D(n8310), .E(n256), .CK(clk), .Q(
        \registers[484][5] ) );
  EDFFX1 \registers_reg[484][4]  ( .D(n8252), .E(n256), .CK(clk), .Q(
        \registers[484][4] ) );
  EDFFX1 \registers_reg[484][3]  ( .D(n8199), .E(n256), .CK(clk), .Q(
        \registers[484][3] ) );
  EDFFX1 \registers_reg[484][2]  ( .D(n8156), .E(n256), .CK(clk), .Q(
        \registers[484][2] ) );
  EDFFX1 \registers_reg[484][1]  ( .D(n8100), .E(n256), .CK(clk), .Q(
        \registers[484][1] ) );
  EDFFX1 \registers_reg[484][0]  ( .D(n8040), .E(n256), .CK(clk), .Q(
        \registers[484][0] ) );
  EDFFX1 \registers_reg[480][7]  ( .D(n8427), .E(n337), .CK(clk), .Q(
        \registers[480][7] ) );
  EDFFX1 \registers_reg[480][6]  ( .D(n8369), .E(n337), .CK(clk), .Q(
        \registers[480][6] ) );
  EDFFX1 \registers_reg[480][5]  ( .D(n8311), .E(n337), .CK(clk), .Q(
        \registers[480][5] ) );
  EDFFX1 \registers_reg[480][4]  ( .D(n8253), .E(n337), .CK(clk), .Q(
        \registers[480][4] ) );
  EDFFX1 \registers_reg[480][3]  ( .D(n8197), .E(n337), .CK(clk), .Q(
        \registers[480][3] ) );
  EDFFX1 \registers_reg[480][2]  ( .D(n8157), .E(n337), .CK(clk), .Q(
        \registers[480][2] ) );
  EDFFX1 \registers_reg[480][1]  ( .D(n8101), .E(n337), .CK(clk), .Q(
        \registers[480][1] ) );
  EDFFX1 \registers_reg[480][0]  ( .D(n8041), .E(n337), .CK(clk), .Q(
        \registers[480][0] ) );
  EDFFX1 \registers_reg[476][7]  ( .D(n8425), .E(n726), .CK(clk), .Q(
        \registers[476][7] ) );
  EDFFX1 \registers_reg[476][6]  ( .D(n8367), .E(n726), .CK(clk), .Q(
        \registers[476][6] ) );
  EDFFX1 \registers_reg[476][5]  ( .D(n8309), .E(n726), .CK(clk), .Q(
        \registers[476][5] ) );
  EDFFX1 \registers_reg[476][4]  ( .D(n8251), .E(n726), .CK(clk), .Q(
        \registers[476][4] ) );
  EDFFX1 \registers_reg[476][3]  ( .D(n8198), .E(n726), .CK(clk), .Q(
        \registers[476][3] ) );
  EDFFX1 \registers_reg[476][2]  ( .D(n8155), .E(n726), .CK(clk), .Q(
        \registers[476][2] ) );
  EDFFX1 \registers_reg[476][1]  ( .D(n8099), .E(n726), .CK(clk), .Q(
        \registers[476][1] ) );
  EDFFX1 \registers_reg[476][0]  ( .D(n8042), .E(n726), .CK(clk), .Q(
        \registers[476][0] ) );
  EDFFX1 \registers_reg[472][7]  ( .D(n8426), .E(n722), .CK(clk), .Q(
        \registers[472][7] ) );
  EDFFX1 \registers_reg[472][6]  ( .D(n8368), .E(n722), .CK(clk), .Q(
        \registers[472][6] ) );
  EDFFX1 \registers_reg[472][5]  ( .D(n8310), .E(n722), .CK(clk), .Q(
        \registers[472][5] ) );
  EDFFX1 \registers_reg[472][4]  ( .D(n8252), .E(n722), .CK(clk), .Q(
        \registers[472][4] ) );
  EDFFX1 \registers_reg[472][3]  ( .D(n8199), .E(n722), .CK(clk), .Q(
        \registers[472][3] ) );
  EDFFX1 \registers_reg[472][2]  ( .D(n8153), .E(n722), .CK(clk), .Q(
        \registers[472][2] ) );
  EDFFX1 \registers_reg[472][1]  ( .D(n8097), .E(n722), .CK(clk), .Q(
        \registers[472][1] ) );
  EDFFX1 \registers_reg[472][0]  ( .D(n8037), .E(n722), .CK(clk), .Q(
        \registers[472][0] ) );
  EDFFX1 \registers_reg[468][7]  ( .D(n8427), .E(n718), .CK(clk), .Q(
        \registers[468][7] ) );
  EDFFX1 \registers_reg[468][6]  ( .D(n8369), .E(n718), .CK(clk), .Q(
        \registers[468][6] ) );
  EDFFX1 \registers_reg[468][5]  ( .D(n8311), .E(n718), .CK(clk), .Q(
        \registers[468][5] ) );
  EDFFX1 \registers_reg[468][4]  ( .D(n8253), .E(n718), .CK(clk), .Q(
        \registers[468][4] ) );
  EDFFX1 \registers_reg[468][3]  ( .D(n8197), .E(n718), .CK(clk), .Q(
        \registers[468][3] ) );
  EDFFX1 \registers_reg[468][2]  ( .D(n8154), .E(n718), .CK(clk), .Q(
        \registers[468][2] ) );
  EDFFX1 \registers_reg[468][1]  ( .D(n8098), .E(n718), .CK(clk), .Q(
        \registers[468][1] ) );
  EDFFX1 \registers_reg[468][0]  ( .D(n8038), .E(n718), .CK(clk), .Q(
        \registers[468][0] ) );
  EDFFX1 \registers_reg[464][7]  ( .D(n8425), .E(n30), .CK(clk), .Q(
        \registers[464][7] ) );
  EDFFX1 \registers_reg[464][6]  ( .D(n8367), .E(n30), .CK(clk), .Q(
        \registers[464][6] ) );
  EDFFX1 \registers_reg[464][5]  ( .D(n8309), .E(n30), .CK(clk), .Q(
        \registers[464][5] ) );
  EDFFX1 \registers_reg[464][4]  ( .D(n8251), .E(n30), .CK(clk), .Q(
        \registers[464][4] ) );
  EDFFX1 \registers_reg[464][3]  ( .D(n8198), .E(n30), .CK(clk), .Q(
        \registers[464][3] ) );
  EDFFX1 \registers_reg[464][2]  ( .D(n8152), .E(n30), .CK(clk), .Q(
        \registers[464][2] ) );
  EDFFX1 \registers_reg[464][1]  ( .D(n8096), .E(n30), .CK(clk), .Q(
        \registers[464][1] ) );
  EDFFX1 \registers_reg[464][0]  ( .D(n8039), .E(n30), .CK(clk), .Q(
        \registers[464][0] ) );
  EDFFX1 \registers_reg[460][7]  ( .D(n8426), .E(n26), .CK(clk), .Q(
        \registers[460][7] ) );
  EDFFX1 \registers_reg[460][6]  ( .D(n8368), .E(n26), .CK(clk), .Q(
        \registers[460][6] ) );
  EDFFX1 \registers_reg[460][5]  ( .D(n8310), .E(n26), .CK(clk), .Q(
        \registers[460][5] ) );
  EDFFX1 \registers_reg[460][4]  ( .D(n8252), .E(n26), .CK(clk), .Q(
        \registers[460][4] ) );
  EDFFX1 \registers_reg[460][3]  ( .D(n8199), .E(n26), .CK(clk), .Q(
        \registers[460][3] ) );
  EDFFX1 \registers_reg[460][2]  ( .D(n8153), .E(n26), .CK(clk), .Q(
        \registers[460][2] ) );
  EDFFX1 \registers_reg[460][1]  ( .D(n8097), .E(n26), .CK(clk), .Q(
        \registers[460][1] ) );
  EDFFX1 \registers_reg[460][0]  ( .D(n8037), .E(n26), .CK(clk), .Q(
        \registers[460][0] ) );
  EDFFX1 \registers_reg[456][7]  ( .D(n8422), .E(n22), .CK(clk), .Q(
        \registers[456][7] ) );
  EDFFX1 \registers_reg[456][6]  ( .D(n8364), .E(n22), .CK(clk), .Q(
        \registers[456][6] ) );
  EDFFX1 \registers_reg[456][5]  ( .D(n8306), .E(n22), .CK(clk), .Q(
        \registers[456][5] ) );
  EDFFX1 \registers_reg[456][4]  ( .D(n8248), .E(n22), .CK(clk), .Q(
        \registers[456][4] ) );
  EDFFX1 \registers_reg[456][3]  ( .D(n8197), .E(n22), .CK(clk), .Q(
        \registers[456][3] ) );
  EDFFX1 \registers_reg[456][2]  ( .D(n8154), .E(n22), .CK(clk), .Q(
        \registers[456][2] ) );
  EDFFX1 \registers_reg[456][1]  ( .D(n8098), .E(n22), .CK(clk), .Q(
        \registers[456][1] ) );
  EDFFX1 \registers_reg[456][0]  ( .D(n8038), .E(n22), .CK(clk), .Q(
        \registers[456][0] ) );
  EDFFX1 \registers_reg[452][7]  ( .D(n8423), .E(n249), .CK(clk), .Q(
        \registers[452][7] ) );
  EDFFX1 \registers_reg[452][6]  ( .D(n8365), .E(n249), .CK(clk), .Q(
        \registers[452][6] ) );
  EDFFX1 \registers_reg[452][5]  ( .D(n8307), .E(n249), .CK(clk), .Q(
        \registers[452][5] ) );
  EDFFX1 \registers_reg[452][4]  ( .D(n8249), .E(n249), .CK(clk), .Q(
        \registers[452][4] ) );
  EDFFX1 \registers_reg[452][3]  ( .D(n8198), .E(n249), .CK(clk), .Q(
        \registers[452][3] ) );
  EDFFX1 \registers_reg[452][2]  ( .D(n8152), .E(n249), .CK(clk), .Q(
        \registers[452][2] ) );
  EDFFX1 \registers_reg[452][1]  ( .D(n8096), .E(n249), .CK(clk), .Q(
        \registers[452][1] ) );
  EDFFX1 \registers_reg[452][0]  ( .D(n8039), .E(n249), .CK(clk), .Q(
        \registers[452][0] ) );
  EDFFX1 \registers_reg[448][7]  ( .D(n8424), .E(n336), .CK(clk), .Q(
        \registers[448][7] ) );
  EDFFX1 \registers_reg[448][6]  ( .D(n8366), .E(n336), .CK(clk), .Q(
        \registers[448][6] ) );
  EDFFX1 \registers_reg[448][5]  ( .D(n8308), .E(n336), .CK(clk), .Q(
        \registers[448][5] ) );
  EDFFX1 \registers_reg[448][4]  ( .D(n8250), .E(n336), .CK(clk), .Q(
        \registers[448][4] ) );
  EDFFX1 \registers_reg[448][3]  ( .D(n8199), .E(n336), .CK(clk), .Q(
        \registers[448][3] ) );
  EDFFX1 \registers_reg[448][2]  ( .D(n8153), .E(n336), .CK(clk), .Q(
        \registers[448][2] ) );
  EDFFX1 \registers_reg[448][1]  ( .D(n8097), .E(n336), .CK(clk), .Q(
        \registers[448][1] ) );
  EDFFX1 \registers_reg[448][0]  ( .D(n8037), .E(n336), .CK(clk), .Q(
        \registers[448][0] ) );
  EDFFX1 \registers_reg[444][7]  ( .D(n8423), .E(n714), .CK(clk), .Q(
        \registers[444][7] ) );
  EDFFX1 \registers_reg[444][6]  ( .D(n8365), .E(n714), .CK(clk), .Q(
        \registers[444][6] ) );
  EDFFX1 \registers_reg[444][5]  ( .D(n8307), .E(n714), .CK(clk), .Q(
        \registers[444][5] ) );
  EDFFX1 \registers_reg[444][4]  ( .D(n8249), .E(n714), .CK(clk), .Q(
        \registers[444][4] ) );
  EDFFX1 \registers_reg[444][3]  ( .D(n8198), .E(n714), .CK(clk), .Q(
        \registers[444][3] ) );
  EDFFX1 \registers_reg[444][2]  ( .D(n8152), .E(n714), .CK(clk), .Q(
        \registers[444][2] ) );
  EDFFX1 \registers_reg[444][1]  ( .D(n8096), .E(n714), .CK(clk), .Q(
        \registers[444][1] ) );
  EDFFX1 \registers_reg[444][0]  ( .D(n8039), .E(n714), .CK(clk), .Q(
        \registers[444][0] ) );
  EDFFX1 \registers_reg[440][7]  ( .D(n8424), .E(n710), .CK(clk), .Q(
        \registers[440][7] ) );
  EDFFX1 \registers_reg[440][6]  ( .D(n8366), .E(n710), .CK(clk), .Q(
        \registers[440][6] ) );
  EDFFX1 \registers_reg[440][5]  ( .D(n8308), .E(n710), .CK(clk), .Q(
        \registers[440][5] ) );
  EDFFX1 \registers_reg[440][4]  ( .D(n8250), .E(n710), .CK(clk), .Q(
        \registers[440][4] ) );
  EDFFX1 \registers_reg[440][3]  ( .D(n8199), .E(n710), .CK(clk), .Q(
        \registers[440][3] ) );
  EDFFX1 \registers_reg[440][2]  ( .D(n8153), .E(n710), .CK(clk), .Q(
        \registers[440][2] ) );
  EDFFX1 \registers_reg[440][1]  ( .D(n8097), .E(n710), .CK(clk), .Q(
        \registers[440][1] ) );
  EDFFX1 \registers_reg[440][0]  ( .D(n8037), .E(n710), .CK(clk), .Q(
        \registers[440][0] ) );
  EDFFX1 \registers_reg[436][7]  ( .D(n8422), .E(n706), .CK(clk), .Q(
        \registers[436][7] ) );
  EDFFX1 \registers_reg[436][6]  ( .D(n8364), .E(n706), .CK(clk), .Q(
        \registers[436][6] ) );
  EDFFX1 \registers_reg[436][5]  ( .D(n8306), .E(n706), .CK(clk), .Q(
        \registers[436][5] ) );
  EDFFX1 \registers_reg[436][4]  ( .D(n8248), .E(n706), .CK(clk), .Q(
        \registers[436][4] ) );
  EDFFX1 \registers_reg[436][3]  ( .D(n8197), .E(n706), .CK(clk), .Q(
        \registers[436][3] ) );
  EDFFX1 \registers_reg[436][2]  ( .D(n8154), .E(n706), .CK(clk), .Q(
        \registers[436][2] ) );
  EDFFX1 \registers_reg[436][1]  ( .D(n8098), .E(n706), .CK(clk), .Q(
        \registers[436][1] ) );
  EDFFX1 \registers_reg[436][0]  ( .D(n8038), .E(n706), .CK(clk), .Q(
        \registers[436][0] ) );
  EDFFX1 \registers_reg[432][7]  ( .D(n8423), .E(n18), .CK(clk), .Q(
        \registers[432][7] ) );
  EDFFX1 \registers_reg[432][6]  ( .D(n8365), .E(n18), .CK(clk), .Q(
        \registers[432][6] ) );
  EDFFX1 \registers_reg[432][5]  ( .D(n8307), .E(n18), .CK(clk), .Q(
        \registers[432][5] ) );
  EDFFX1 \registers_reg[432][4]  ( .D(n8249), .E(n18), .CK(clk), .Q(
        \registers[432][4] ) );
  EDFFX1 \registers_reg[432][3]  ( .D(n8198), .E(n18), .CK(clk), .Q(
        \registers[432][3] ) );
  EDFFX1 \registers_reg[432][2]  ( .D(n8152), .E(n18), .CK(clk), .Q(
        \registers[432][2] ) );
  EDFFX1 \registers_reg[432][1]  ( .D(n8096), .E(n18), .CK(clk), .Q(
        \registers[432][1] ) );
  EDFFX1 \registers_reg[432][0]  ( .D(n8039), .E(n18), .CK(clk), .Q(
        \registers[432][0] ) );
  EDFFX1 \registers_reg[428][7]  ( .D(n8424), .E(n14), .CK(clk), .Q(
        \registers[428][7] ) );
  EDFFX1 \registers_reg[428][6]  ( .D(n8366), .E(n14), .CK(clk), .Q(
        \registers[428][6] ) );
  EDFFX1 \registers_reg[428][5]  ( .D(n8308), .E(n14), .CK(clk), .Q(
        \registers[428][5] ) );
  EDFFX1 \registers_reg[428][4]  ( .D(n8250), .E(n14), .CK(clk), .Q(
        \registers[428][4] ) );
  EDFFX1 \registers_reg[428][3]  ( .D(n8199), .E(n14), .CK(clk), .Q(
        \registers[428][3] ) );
  EDFFX1 \registers_reg[428][2]  ( .D(n8153), .E(n14), .CK(clk), .Q(
        \registers[428][2] ) );
  EDFFX1 \registers_reg[428][1]  ( .D(n8097), .E(n14), .CK(clk), .Q(
        \registers[428][1] ) );
  EDFFX1 \registers_reg[428][0]  ( .D(n8037), .E(n14), .CK(clk), .Q(
        \registers[428][0] ) );
  EDFFX1 \registers_reg[424][7]  ( .D(n8422), .E(n10), .CK(clk), .Q(
        \registers[424][7] ) );
  EDFFX1 \registers_reg[424][6]  ( .D(n8364), .E(n10), .CK(clk), .Q(
        \registers[424][6] ) );
  EDFFX1 \registers_reg[424][5]  ( .D(n8306), .E(n10), .CK(clk), .Q(
        \registers[424][5] ) );
  EDFFX1 \registers_reg[424][4]  ( .D(n8248), .E(n10), .CK(clk), .Q(
        \registers[424][4] ) );
  EDFFX1 \registers_reg[424][3]  ( .D(n8194), .E(n10), .CK(clk), .Q(
        \registers[424][3] ) );
  EDFFX1 \registers_reg[424][2]  ( .D(n8154), .E(n10), .CK(clk), .Q(
        \registers[424][2] ) );
  EDFFX1 \registers_reg[424][1]  ( .D(n8098), .E(n10), .CK(clk), .Q(
        \registers[424][1] ) );
  EDFFX1 \registers_reg[424][0]  ( .D(n8038), .E(n10), .CK(clk), .Q(
        \registers[424][0] ) );
  EDFFX1 \registers_reg[420][7]  ( .D(n8423), .E(n242), .CK(clk), .Q(
        \registers[420][7] ) );
  EDFFX1 \registers_reg[420][6]  ( .D(n8365), .E(n242), .CK(clk), .Q(
        \registers[420][6] ) );
  EDFFX1 \registers_reg[420][5]  ( .D(n8307), .E(n242), .CK(clk), .Q(
        \registers[420][5] ) );
  EDFFX1 \registers_reg[420][4]  ( .D(n8249), .E(n242), .CK(clk), .Q(
        \registers[420][4] ) );
  EDFFX1 \registers_reg[420][3]  ( .D(n8195), .E(n242), .CK(clk), .Q(
        \registers[420][3] ) );
  EDFFX1 \registers_reg[420][2]  ( .D(n8150), .E(n242), .CK(clk), .Q(
        \registers[420][2] ) );
  EDFFX1 \registers_reg[420][1]  ( .D(n8094), .E(n242), .CK(clk), .Q(
        \registers[420][1] ) );
  EDFFX1 \registers_reg[420][0]  ( .D(n8036), .E(n242), .CK(clk), .Q(
        \registers[420][0] ) );
  EDFFX1 \registers_reg[416][7]  ( .D(n8424), .E(n335), .CK(clk), .Q(
        \registers[416][7] ) );
  EDFFX1 \registers_reg[416][6]  ( .D(n8366), .E(n335), .CK(clk), .Q(
        \registers[416][6] ) );
  EDFFX1 \registers_reg[416][5]  ( .D(n8308), .E(n335), .CK(clk), .Q(
        \registers[416][5] ) );
  EDFFX1 \registers_reg[416][4]  ( .D(n8250), .E(n335), .CK(clk), .Q(
        \registers[416][4] ) );
  EDFFX1 \registers_reg[416][3]  ( .D(n8196), .E(n335), .CK(clk), .Q(
        \registers[416][3] ) );
  EDFFX1 \registers_reg[416][2]  ( .D(n8151), .E(n335), .CK(clk), .Q(
        \registers[416][2] ) );
  EDFFX1 \registers_reg[416][1]  ( .D(n8095), .E(n335), .CK(clk), .Q(
        \registers[416][1] ) );
  EDFFX1 \registers_reg[416][0]  ( .D(n8034), .E(n335), .CK(clk), .Q(
        \registers[416][0] ) );
  EDFFX1 \registers_reg[412][7]  ( .D(n8422), .E(n702), .CK(clk), .Q(
        \registers[412][7] ) );
  EDFFX1 \registers_reg[412][6]  ( .D(n8364), .E(n702), .CK(clk), .Q(
        \registers[412][6] ) );
  EDFFX1 \registers_reg[412][5]  ( .D(n8306), .E(n702), .CK(clk), .Q(
        \registers[412][5] ) );
  EDFFX1 \registers_reg[412][4]  ( .D(n8248), .E(n702), .CK(clk), .Q(
        \registers[412][4] ) );
  EDFFX1 \registers_reg[412][3]  ( .D(n8194), .E(n702), .CK(clk), .Q(
        \registers[412][3] ) );
  EDFFX1 \registers_reg[412][2]  ( .D(n8736), .E(n702), .CK(clk), .Q(
        \registers[412][2] ) );
  EDFFX1 \registers_reg[412][1]  ( .D(n8708), .E(n702), .CK(clk), .Q(
        \registers[412][1] ) );
  EDFFX1 \registers_reg[412][0]  ( .D(n8035), .E(n702), .CK(clk), .Q(
        \registers[412][0] ) );
  EDFFX1 \registers_reg[408][7]  ( .D(n8423), .E(n698), .CK(clk), .Q(
        \registers[408][7] ) );
  EDFFX1 \registers_reg[408][6]  ( .D(n8365), .E(n698), .CK(clk), .Q(
        \registers[408][6] ) );
  EDFFX1 \registers_reg[408][5]  ( .D(n8307), .E(n698), .CK(clk), .Q(
        \registers[408][5] ) );
  EDFFX1 \registers_reg[408][4]  ( .D(n8249), .E(n698), .CK(clk), .Q(
        \registers[408][4] ) );
  EDFFX1 \registers_reg[408][3]  ( .D(n8195), .E(n698), .CK(clk), .Q(
        \registers[408][3] ) );
  EDFFX1 \registers_reg[408][2]  ( .D(n8150), .E(n698), .CK(clk), .Q(
        \registers[408][2] ) );
  EDFFX1 \registers_reg[408][1]  ( .D(n8094), .E(n698), .CK(clk), .Q(
        \registers[408][1] ) );
  EDFFX1 \registers_reg[408][0]  ( .D(n8036), .E(n698), .CK(clk), .Q(
        \registers[408][0] ) );
  EDFFX1 \registers_reg[404][7]  ( .D(n8419), .E(n694), .CK(clk), .Q(
        \registers[404][7] ) );
  EDFFX1 \registers_reg[404][6]  ( .D(n8361), .E(n694), .CK(clk), .Q(
        \registers[404][6] ) );
  EDFFX1 \registers_reg[404][5]  ( .D(n8303), .E(n694), .CK(clk), .Q(
        \registers[404][5] ) );
  EDFFX1 \registers_reg[404][4]  ( .D(n8245), .E(n694), .CK(clk), .Q(
        \registers[404][4] ) );
  EDFFX1 \registers_reg[404][3]  ( .D(n8196), .E(n694), .CK(clk), .Q(
        \registers[404][3] ) );
  EDFFX1 \registers_reg[404][2]  ( .D(n8151), .E(n694), .CK(clk), .Q(
        \registers[404][2] ) );
  EDFFX1 \registers_reg[404][1]  ( .D(n8095), .E(n694), .CK(clk), .Q(
        \registers[404][1] ) );
  EDFFX1 \registers_reg[404][0]  ( .D(n8034), .E(n694), .CK(clk), .Q(
        \registers[404][0] ) );
  EDFFX1 \registers_reg[400][7]  ( .D(n8420), .E(n690), .CK(clk), .Q(
        \registers[400][7] ) );
  EDFFX1 \registers_reg[400][6]  ( .D(n8362), .E(n690), .CK(clk), .Q(
        \registers[400][6] ) );
  EDFFX1 \registers_reg[400][5]  ( .D(n8304), .E(n690), .CK(clk), .Q(
        \registers[400][5] ) );
  EDFFX1 \registers_reg[400][4]  ( .D(n8246), .E(n690), .CK(clk), .Q(
        \registers[400][4] ) );
  EDFFX1 \registers_reg[400][3]  ( .D(n8194), .E(n690), .CK(clk), .Q(
        \registers[400][3] ) );
  EDFFX1 \registers_reg[400][2]  ( .D(n8735), .E(n690), .CK(clk), .Q(
        \registers[400][2] ) );
  EDFFX1 \registers_reg[400][1]  ( .D(n8707), .E(n690), .CK(clk), .Q(
        \registers[400][1] ) );
  EDFFX1 \registers_reg[400][0]  ( .D(n8035), .E(n690), .CK(clk), .Q(
        \registers[400][0] ) );
  EDFFX1 \registers_reg[396][7]  ( .D(n8421), .E(n686), .CK(clk), .Q(
        \registers[396][7] ) );
  EDFFX1 \registers_reg[396][6]  ( .D(n8363), .E(n686), .CK(clk), .Q(
        \registers[396][6] ) );
  EDFFX1 \registers_reg[396][5]  ( .D(n8305), .E(n686), .CK(clk), .Q(
        \registers[396][5] ) );
  EDFFX1 \registers_reg[396][4]  ( .D(n8247), .E(n686), .CK(clk), .Q(
        \registers[396][4] ) );
  EDFFX1 \registers_reg[396][3]  ( .D(n8195), .E(n686), .CK(clk), .Q(
        \registers[396][3] ) );
  EDFFX1 \registers_reg[396][2]  ( .D(n8150), .E(n686), .CK(clk), .Q(
        \registers[396][2] ) );
  EDFFX1 \registers_reg[396][1]  ( .D(n8094), .E(n686), .CK(clk), .Q(
        \registers[396][1] ) );
  EDFFX1 \registers_reg[396][0]  ( .D(n8036), .E(n686), .CK(clk), .Q(
        \registers[396][0] ) );
  EDFFX1 \registers_reg[392][7]  ( .D(n8419), .E(n682), .CK(clk), .Q(
        \registers[392][7] ) );
  EDFFX1 \registers_reg[392][6]  ( .D(n8361), .E(n682), .CK(clk), .Q(
        \registers[392][6] ) );
  EDFFX1 \registers_reg[392][5]  ( .D(n8303), .E(n682), .CK(clk), .Q(
        \registers[392][5] ) );
  EDFFX1 \registers_reg[392][4]  ( .D(n8245), .E(n682), .CK(clk), .Q(
        \registers[392][4] ) );
  EDFFX1 \registers_reg[392][3]  ( .D(n8196), .E(n682), .CK(clk), .Q(
        \registers[392][3] ) );
  EDFFX1 \registers_reg[392][2]  ( .D(n8151), .E(n682), .CK(clk), .Q(
        \registers[392][2] ) );
  EDFFX1 \registers_reg[392][1]  ( .D(n8095), .E(n682), .CK(clk), .Q(
        \registers[392][1] ) );
  EDFFX1 \registers_reg[392][0]  ( .D(n8034), .E(n682), .CK(clk), .Q(
        \registers[392][0] ) );
  EDFFX1 \registers_reg[388][7]  ( .D(n8420), .E(n998), .CK(clk), .Q(
        \registers[388][7] ) );
  EDFFX1 \registers_reg[388][6]  ( .D(n8362), .E(n998), .CK(clk), .Q(
        \registers[388][6] ) );
  EDFFX1 \registers_reg[388][5]  ( .D(n8304), .E(n998), .CK(clk), .Q(
        \registers[388][5] ) );
  EDFFX1 \registers_reg[388][4]  ( .D(n8246), .E(n998), .CK(clk), .Q(
        \registers[388][4] ) );
  EDFFX1 \registers_reg[388][3]  ( .D(n8194), .E(n998), .CK(clk), .Q(
        \registers[388][3] ) );
  EDFFX1 \registers_reg[388][2]  ( .D(n8734), .E(n998), .CK(clk), .Q(
        \registers[388][2] ) );
  EDFFX1 \registers_reg[388][1]  ( .D(n8706), .E(n998), .CK(clk), .Q(
        \registers[388][1] ) );
  EDFFX1 \registers_reg[388][0]  ( .D(n8035), .E(n998), .CK(clk), .Q(
        \registers[388][0] ) );
  EDFFX1 \registers_reg[384][7]  ( .D(n8422), .E(n334), .CK(clk), .Q(
        \registers[384][7] ) );
  EDFFX1 \registers_reg[384][6]  ( .D(n8364), .E(n334), .CK(clk), .Q(
        \registers[384][6] ) );
  EDFFX1 \registers_reg[384][5]  ( .D(n8306), .E(n334), .CK(clk), .Q(
        \registers[384][5] ) );
  EDFFX1 \registers_reg[384][4]  ( .D(n8248), .E(n334), .CK(clk), .Q(
        \registers[384][4] ) );
  EDFFX1 \registers_reg[384][3]  ( .D(n8197), .E(n334), .CK(clk), .Q(
        \registers[384][3] ) );
  EDFFX1 \registers_reg[384][2]  ( .D(n8154), .E(n334), .CK(clk), .Q(
        \registers[384][2] ) );
  EDFFX1 \registers_reg[384][1]  ( .D(n8098), .E(n334), .CK(clk), .Q(
        \registers[384][1] ) );
  EDFFX1 \registers_reg[384][0]  ( .D(n8036), .E(n334), .CK(clk), .Q(
        \registers[384][0] ) );
  EDFFX1 \registers_reg[380][7]  ( .D(n8433), .E(n678), .CK(clk), .Q(
        \registers[380][7] ) );
  EDFFX1 \registers_reg[380][6]  ( .D(n8375), .E(n678), .CK(clk), .Q(
        \registers[380][6] ) );
  EDFFX1 \registers_reg[380][5]  ( .D(n8317), .E(n678), .CK(clk), .Q(
        \registers[380][5] ) );
  EDFFX1 \registers_reg[380][4]  ( .D(n8259), .E(n678), .CK(clk), .Q(
        \registers[380][4] ) );
  EDFFX1 \registers_reg[380][3]  ( .D(n8194), .E(n678), .CK(clk), .Q(
        \registers[380][3] ) );
  EDFFX1 \registers_reg[380][2]  ( .D(n8112), .E(n678), .CK(clk), .Q(
        \registers[380][2] ) );
  EDFFX1 \registers_reg[380][1]  ( .D(n8056), .E(n678), .CK(clk), .Q(
        \registers[380][1] ) );
  EDFFX1 \registers_reg[380][0]  ( .D(n7998), .E(n678), .CK(clk), .Q(
        \registers[380][0] ) );
  EDFFX1 \registers_reg[376][7]  ( .D(n8434), .E(n674), .CK(clk), .Q(
        \registers[376][7] ) );
  EDFFX1 \registers_reg[376][6]  ( .D(n8376), .E(n674), .CK(clk), .Q(
        \registers[376][6] ) );
  EDFFX1 \registers_reg[376][5]  ( .D(n8318), .E(n674), .CK(clk), .Q(
        \registers[376][5] ) );
  EDFFX1 \registers_reg[376][4]  ( .D(n8260), .E(n674), .CK(clk), .Q(
        \registers[376][4] ) );
  EDFFX1 \registers_reg[376][3]  ( .D(n8195), .E(n674), .CK(clk), .Q(
        \registers[376][3] ) );
  EDFFX1 \registers_reg[376][2]  ( .D(n8113), .E(n674), .CK(clk), .Q(
        \registers[376][2] ) );
  EDFFX1 \registers_reg[376][1]  ( .D(n8057), .E(n674), .CK(clk), .Q(
        \registers[376][1] ) );
  EDFFX1 \registers_reg[376][0]  ( .D(n8004), .E(n674), .CK(clk), .Q(
        \registers[376][0] ) );
  EDFFX1 \registers_reg[372][7]  ( .D(n8434), .E(n670), .CK(clk), .Q(
        \registers[372][7] ) );
  EDFFX1 \registers_reg[372][6]  ( .D(n8376), .E(n670), .CK(clk), .Q(
        \registers[372][6] ) );
  EDFFX1 \registers_reg[372][5]  ( .D(n8318), .E(n670), .CK(clk), .Q(
        \registers[372][5] ) );
  EDFFX1 \registers_reg[372][4]  ( .D(n8260), .E(n670), .CK(clk), .Q(
        \registers[372][4] ) );
  EDFFX1 \registers_reg[372][3]  ( .D(n8196), .E(n670), .CK(clk), .Q(
        \registers[372][3] ) );
  EDFFX1 \registers_reg[372][2]  ( .D(n8111), .E(n670), .CK(clk), .Q(
        \registers[372][2] ) );
  EDFFX1 \registers_reg[372][1]  ( .D(n8055), .E(n670), .CK(clk), .Q(
        \registers[372][1] ) );
  EDFFX1 \registers_reg[372][0]  ( .D(n7999), .E(n670), .CK(clk), .Q(
        \registers[372][0] ) );
  EDFFX1 \registers_reg[368][7]  ( .D(n8433), .E(n666), .CK(clk), .Q(
        \registers[368][7] ) );
  EDFFX1 \registers_reg[368][6]  ( .D(n8375), .E(n666), .CK(clk), .Q(
        \registers[368][6] ) );
  EDFFX1 \registers_reg[368][5]  ( .D(n8317), .E(n666), .CK(clk), .Q(
        \registers[368][5] ) );
  EDFFX1 \registers_reg[368][4]  ( .D(n8259), .E(n666), .CK(clk), .Q(
        \registers[368][4] ) );
  EDFFX1 \registers_reg[368][3]  ( .D(n8191), .E(n666), .CK(clk), .Q(
        \registers[368][3] ) );
  EDFFX1 \registers_reg[368][2]  ( .D(n8138), .E(n666), .CK(clk), .Q(
        \registers[368][2] ) );
  EDFFX1 \registers_reg[368][1]  ( .D(n8082), .E(n666), .CK(clk), .Q(
        \registers[368][1] ) );
  EDFFX1 \registers_reg[368][0]  ( .D(n8048), .E(n666), .CK(clk), .Q(
        \registers[368][0] ) );
  EDFFX1 \registers_reg[364][7]  ( .D(n8434), .E(n662), .CK(clk), .Q(
        \registers[364][7] ) );
  EDFFX1 \registers_reg[364][6]  ( .D(n8376), .E(n662), .CK(clk), .Q(
        \registers[364][6] ) );
  EDFFX1 \registers_reg[364][5]  ( .D(n8318), .E(n662), .CK(clk), .Q(
        \registers[364][5] ) );
  EDFFX1 \registers_reg[364][4]  ( .D(n8260), .E(n662), .CK(clk), .Q(
        \registers[364][4] ) );
  EDFFX1 \registers_reg[364][3]  ( .D(n8192), .E(n662), .CK(clk), .Q(
        \registers[364][3] ) );
  EDFFX1 \registers_reg[364][2]  ( .D(n8157), .E(n662), .CK(clk), .Q(
        \registers[364][2] ) );
  EDFFX1 \registers_reg[364][1]  ( .D(n8101), .E(n662), .CK(clk), .Q(
        \registers[364][1] ) );
  EDFFX1 \registers_reg[364][0]  ( .D(n8046), .E(n662), .CK(clk), .Q(
        \registers[364][0] ) );
  EDFFX1 \registers_reg[360][7]  ( .D(n8433), .E(n658), .CK(clk), .Q(
        \registers[360][7] ) );
  EDFFX1 \registers_reg[360][6]  ( .D(n8375), .E(n658), .CK(clk), .Q(
        \registers[360][6] ) );
  EDFFX1 \registers_reg[360][5]  ( .D(n8317), .E(n658), .CK(clk), .Q(
        \registers[360][5] ) );
  EDFFX1 \registers_reg[360][4]  ( .D(n8259), .E(n658), .CK(clk), .Q(
        \registers[360][4] ) );
  EDFFX1 \registers_reg[360][3]  ( .D(n8193), .E(n658), .CK(clk), .Q(
        \registers[360][3] ) );
  EDFFX1 \registers_reg[360][2]  ( .D(n8125), .E(n658), .CK(clk), .Q(
        \registers[360][2] ) );
  EDFFX1 \registers_reg[360][1]  ( .D(n8069), .E(n658), .CK(clk), .Q(
        \registers[360][1] ) );
  EDFFX1 \registers_reg[360][0]  ( .D(n8047), .E(n658), .CK(clk), .Q(
        \registers[360][0] ) );
  EDFFX1 \registers_reg[356][7]  ( .D(n8433), .E(n991), .CK(clk), .Q(
        \registers[356][7] ) );
  EDFFX1 \registers_reg[356][6]  ( .D(n8375), .E(n991), .CK(clk), .Q(
        \registers[356][6] ) );
  EDFFX1 \registers_reg[356][5]  ( .D(n8317), .E(n991), .CK(clk), .Q(
        \registers[356][5] ) );
  EDFFX1 \registers_reg[356][4]  ( .D(n8259), .E(n991), .CK(clk), .Q(
        \registers[356][4] ) );
  EDFFX1 \registers_reg[356][3]  ( .D(n8200), .E(n991), .CK(clk), .Q(
        \registers[356][3] ) );
  EDFFX1 \registers_reg[356][2]  ( .D(n8139), .E(n991), .CK(clk), .Q(
        \registers[356][2] ) );
  EDFFX1 \registers_reg[356][1]  ( .D(n8083), .E(n991), .CK(clk), .Q(
        \registers[356][1] ) );
  EDFFX1 \registers_reg[356][0]  ( .D(n8048), .E(n991), .CK(clk), .Q(
        \registers[356][0] ) );
  EDFFX1 \registers_reg[352][7]  ( .D(n8434), .E(n333), .CK(clk), .Q(
        \registers[352][7] ) );
  EDFFX1 \registers_reg[352][6]  ( .D(n8376), .E(n333), .CK(clk), .Q(
        \registers[352][6] ) );
  EDFFX1 \registers_reg[352][5]  ( .D(n8318), .E(n333), .CK(clk), .Q(
        \registers[352][5] ) );
  EDFFX1 \registers_reg[352][4]  ( .D(n8260), .E(n333), .CK(clk), .Q(
        \registers[352][4] ) );
  EDFFX1 \registers_reg[352][3]  ( .D(n8165), .E(n333), .CK(clk), .Q(
        \registers[352][3] ) );
  EDFFX1 \registers_reg[352][2]  ( .D(n8155), .E(n333), .CK(clk), .Q(
        \registers[352][2] ) );
  EDFFX1 \registers_reg[352][1]  ( .D(n8099), .E(n333), .CK(clk), .Q(
        \registers[352][1] ) );
  EDFFX1 \registers_reg[352][0]  ( .D(n8046), .E(n333), .CK(clk), .Q(
        \registers[352][0] ) );
  EDFFX1 \registers_reg[348][7]  ( .D(n8430), .E(n654), .CK(clk), .Q(
        \registers[348][7] ) );
  EDFFX1 \registers_reg[348][6]  ( .D(n8372), .E(n654), .CK(clk), .Q(
        \registers[348][6] ) );
  EDFFX1 \registers_reg[348][5]  ( .D(n8314), .E(n654), .CK(clk), .Q(
        \registers[348][5] ) );
  EDFFX1 \registers_reg[348][4]  ( .D(n8256), .E(n654), .CK(clk), .Q(
        \registers[348][4] ) );
  EDFFX1 \registers_reg[348][3]  ( .D(n8181), .E(n654), .CK(clk), .Q(
        \registers[348][3] ) );
  EDFFX1 \registers_reg[348][2]  ( .D(n8120), .E(n654), .CK(clk), .Q(
        \registers[348][2] ) );
  EDFFX1 \registers_reg[348][1]  ( .D(n8064), .E(n654), .CK(clk), .Q(
        \registers[348][1] ) );
  EDFFX1 \registers_reg[348][0]  ( .D(n8047), .E(n654), .CK(clk), .Q(
        \registers[348][0] ) );
  EDFFX1 \registers_reg[344][7]  ( .D(n8431), .E(n650), .CK(clk), .Q(
        \registers[344][7] ) );
  EDFFX1 \registers_reg[344][6]  ( .D(n8373), .E(n650), .CK(clk), .Q(
        \registers[344][6] ) );
  EDFFX1 \registers_reg[344][5]  ( .D(n8315), .E(n650), .CK(clk), .Q(
        \registers[344][5] ) );
  EDFFX1 \registers_reg[344][4]  ( .D(n8257), .E(n650), .CK(clk), .Q(
        \registers[344][4] ) );
  EDFFX1 \registers_reg[344][3]  ( .D(n8201), .E(n650), .CK(clk), .Q(
        \registers[344][3] ) );
  EDFFX1 \registers_reg[344][2]  ( .D(n8140), .E(n650), .CK(clk), .Q(
        \registers[344][2] ) );
  EDFFX1 \registers_reg[344][1]  ( .D(n8084), .E(n650), .CK(clk), .Q(
        \registers[344][1] ) );
  EDFFX1 \registers_reg[344][0]  ( .D(n8048), .E(n650), .CK(clk), .Q(
        \registers[344][0] ) );
  EDFFX1 \registers_reg[340][7]  ( .D(n8432), .E(n646), .CK(clk), .Q(
        \registers[340][7] ) );
  EDFFX1 \registers_reg[340][6]  ( .D(n8374), .E(n646), .CK(clk), .Q(
        \registers[340][6] ) );
  EDFFX1 \registers_reg[340][5]  ( .D(n8316), .E(n646), .CK(clk), .Q(
        \registers[340][5] ) );
  EDFFX1 \registers_reg[340][4]  ( .D(n8258), .E(n646), .CK(clk), .Q(
        \registers[340][4] ) );
  EDFFX1 \registers_reg[340][3]  ( .D(n8187), .E(n646), .CK(clk), .Q(
        \registers[340][3] ) );
  EDFFX1 \registers_reg[340][2]  ( .D(n8159), .E(n646), .CK(clk), .Q(
        \registers[340][2] ) );
  EDFFX1 \registers_reg[340][1]  ( .D(n8103), .E(n646), .CK(clk), .Q(
        \registers[340][1] ) );
  EDFFX1 \registers_reg[340][0]  ( .D(n8046), .E(n646), .CK(clk), .Q(
        \registers[340][0] ) );
  EDFFX1 \registers_reg[336][7]  ( .D(n8430), .E(n642), .CK(clk), .Q(
        \registers[336][7] ) );
  EDFFX1 \registers_reg[336][6]  ( .D(n8372), .E(n642), .CK(clk), .Q(
        \registers[336][6] ) );
  EDFFX1 \registers_reg[336][5]  ( .D(n8314), .E(n642), .CK(clk), .Q(
        \registers[336][5] ) );
  EDFFX1 \registers_reg[336][4]  ( .D(n8256), .E(n642), .CK(clk), .Q(
        \registers[336][4] ) );
  EDFFX1 \registers_reg[336][3]  ( .D(n8177), .E(n642), .CK(clk), .Q(
        \registers[336][3] ) );
  EDFFX1 \registers_reg[336][2]  ( .D(n8121), .E(n642), .CK(clk), .Q(
        \registers[336][2] ) );
  EDFFX1 \registers_reg[336][1]  ( .D(n8065), .E(n642), .CK(clk), .Q(
        \registers[336][1] ) );
  EDFFX1 \registers_reg[336][0]  ( .D(n8047), .E(n642), .CK(clk), .Q(
        \registers[336][0] ) );
  EDFFX1 \registers_reg[332][7]  ( .D(n8431), .E(n638), .CK(clk), .Q(
        \registers[332][7] ) );
  EDFFX1 \registers_reg[332][6]  ( .D(n8373), .E(n638), .CK(clk), .Q(
        \registers[332][6] ) );
  EDFFX1 \registers_reg[332][5]  ( .D(n8315), .E(n638), .CK(clk), .Q(
        \registers[332][5] ) );
  EDFFX1 \registers_reg[332][4]  ( .D(n8257), .E(n638), .CK(clk), .Q(
        \registers[332][4] ) );
  EDFFX1 \registers_reg[332][3]  ( .D(n8197), .E(n638), .CK(clk), .Q(
        \registers[332][3] ) );
  EDFFX1 \registers_reg[332][2]  ( .D(n8147), .E(n638), .CK(clk), .Q(
        \registers[332][2] ) );
  EDFFX1 \registers_reg[332][1]  ( .D(n8091), .E(n638), .CK(clk), .Q(
        \registers[332][1] ) );
  EDFFX1 \registers_reg[332][0]  ( .D(n8048), .E(n638), .CK(clk), .Q(
        \registers[332][0] ) );
  EDFFX1 \registers_reg[328][7]  ( .D(n8432), .E(n634), .CK(clk), .Q(
        \registers[328][7] ) );
  EDFFX1 \registers_reg[328][6]  ( .D(n8374), .E(n634), .CK(clk), .Q(
        \registers[328][6] ) );
  EDFFX1 \registers_reg[328][5]  ( .D(n8316), .E(n634), .CK(clk), .Q(
        \registers[328][5] ) );
  EDFFX1 \registers_reg[328][4]  ( .D(n8258), .E(n634), .CK(clk), .Q(
        \registers[328][4] ) );
  EDFFX1 \registers_reg[328][3]  ( .D(n8170), .E(n634), .CK(clk), .Q(
        \registers[328][3] ) );
  EDFFX1 \registers_reg[328][2]  ( .D(n8160), .E(n634), .CK(clk), .Q(
        \registers[328][2] ) );
  EDFFX1 \registers_reg[328][1]  ( .D(n8104), .E(n634), .CK(clk), .Q(
        \registers[328][1] ) );
  EDFFX1 \registers_reg[328][0]  ( .D(n8046), .E(n634), .CK(clk), .Q(
        \registers[328][0] ) );
  EDFFX1 \registers_reg[324][7]  ( .D(n8430), .E(n984), .CK(clk), .Q(
        \registers[324][7] ) );
  EDFFX1 \registers_reg[324][6]  ( .D(n8372), .E(n984), .CK(clk), .Q(
        \registers[324][6] ) );
  EDFFX1 \registers_reg[324][5]  ( .D(n8314), .E(n984), .CK(clk), .Q(
        \registers[324][5] ) );
  EDFFX1 \registers_reg[324][4]  ( .D(n8256), .E(n984), .CK(clk), .Q(
        \registers[324][4] ) );
  EDFFX1 \registers_reg[324][3]  ( .D(n8178), .E(n984), .CK(clk), .Q(
        \registers[324][3] ) );
  EDFFX1 \registers_reg[324][2]  ( .D(n8122), .E(n984), .CK(clk), .Q(
        \registers[324][2] ) );
  EDFFX1 \registers_reg[324][1]  ( .D(n8066), .E(n984), .CK(clk), .Q(
        \registers[324][1] ) );
  EDFFX1 \registers_reg[324][0]  ( .D(n8047), .E(n984), .CK(clk), .Q(
        \registers[324][0] ) );
  EDFFX1 \registers_reg[320][7]  ( .D(n8432), .E(n332), .CK(clk), .Q(
        \registers[320][7] ) );
  EDFFX1 \registers_reg[320][6]  ( .D(n8374), .E(n332), .CK(clk), .Q(
        \registers[320][6] ) );
  EDFFX1 \registers_reg[320][5]  ( .D(n8316), .E(n332), .CK(clk), .Q(
        \registers[320][5] ) );
  EDFFX1 \registers_reg[320][4]  ( .D(n8258), .E(n332), .CK(clk), .Q(
        \registers[320][4] ) );
  EDFFX1 \registers_reg[320][3]  ( .D(n8171), .E(n332), .CK(clk), .Q(
        \registers[320][3] ) );
  EDFFX1 \registers_reg[320][2]  ( .D(n8159), .E(n332), .CK(clk), .Q(
        \registers[320][2] ) );
  EDFFX1 \registers_reg[320][1]  ( .D(n8103), .E(n332), .CK(clk), .Q(
        \registers[320][1] ) );
  EDFFX1 \registers_reg[320][0]  ( .D(n8048), .E(n332), .CK(clk), .Q(
        \registers[320][0] ) );
  EDFFX1 \registers_reg[316][7]  ( .D(n8430), .E(n630), .CK(clk), .Q(
        \registers[316][7] ) );
  EDFFX1 \registers_reg[316][6]  ( .D(n8372), .E(n630), .CK(clk), .Q(
        \registers[316][6] ) );
  EDFFX1 \registers_reg[316][5]  ( .D(n8314), .E(n630), .CK(clk), .Q(
        \registers[316][5] ) );
  EDFFX1 \registers_reg[316][4]  ( .D(n8256), .E(n630), .CK(clk), .Q(
        \registers[316][4] ) );
  EDFFX1 \registers_reg[316][3]  ( .D(n8176), .E(n630), .CK(clk), .Q(
        \registers[316][3] ) );
  EDFFX1 \registers_reg[316][2]  ( .D(n8160), .E(n630), .CK(clk), .Q(
        \registers[316][2] ) );
  EDFFX1 \registers_reg[316][1]  ( .D(n8104), .E(n630), .CK(clk), .Q(
        \registers[316][1] ) );
  EDFFX1 \registers_reg[316][0]  ( .D(n8044), .E(n630), .CK(clk), .Q(
        \registers[316][0] ) );
  EDFFX1 \registers_reg[312][7]  ( .D(n8431), .E(n626), .CK(clk), .Q(
        \registers[312][7] ) );
  EDFFX1 \registers_reg[312][6]  ( .D(n8373), .E(n626), .CK(clk), .Q(
        \registers[312][6] ) );
  EDFFX1 \registers_reg[312][5]  ( .D(n8315), .E(n626), .CK(clk), .Q(
        \registers[312][5] ) );
  EDFFX1 \registers_reg[312][4]  ( .D(n8257), .E(n626), .CK(clk), .Q(
        \registers[312][4] ) );
  EDFFX1 \registers_reg[312][3]  ( .D(n8198), .E(n626), .CK(clk), .Q(
        \registers[312][3] ) );
  EDFFX1 \registers_reg[312][2]  ( .D(n8158), .E(n626), .CK(clk), .Q(
        \registers[312][2] ) );
  EDFFX1 \registers_reg[312][1]  ( .D(n8102), .E(n626), .CK(clk), .Q(
        \registers[312][1] ) );
  EDFFX1 \registers_reg[312][0]  ( .D(n8045), .E(n626), .CK(clk), .Q(
        \registers[312][0] ) );
  EDFFX1 \registers_reg[308][7]  ( .D(n8432), .E(n622), .CK(clk), .Q(
        \registers[308][7] ) );
  EDFFX1 \registers_reg[308][6]  ( .D(n8374), .E(n622), .CK(clk), .Q(
        \registers[308][6] ) );
  EDFFX1 \registers_reg[308][5]  ( .D(n8316), .E(n622), .CK(clk), .Q(
        \registers[308][5] ) );
  EDFFX1 \registers_reg[308][4]  ( .D(n8258), .E(n622), .CK(clk), .Q(
        \registers[308][4] ) );
  EDFFX1 \registers_reg[308][3]  ( .D(n8172), .E(n622), .CK(clk), .Q(
        \registers[308][3] ) );
  EDFFX1 \registers_reg[308][2]  ( .D(n8159), .E(n622), .CK(clk), .Q(
        \registers[308][2] ) );
  EDFFX1 \registers_reg[308][1]  ( .D(n8103), .E(n622), .CK(clk), .Q(
        \registers[308][1] ) );
  EDFFX1 \registers_reg[308][0]  ( .D(n8043), .E(n622), .CK(clk), .Q(
        \registers[308][0] ) );
  EDFFX1 \registers_reg[304][7]  ( .D(n8430), .E(n618), .CK(clk), .Q(
        \registers[304][7] ) );
  EDFFX1 \registers_reg[304][6]  ( .D(n8372), .E(n618), .CK(clk), .Q(
        \registers[304][6] ) );
  EDFFX1 \registers_reg[304][5]  ( .D(n8314), .E(n618), .CK(clk), .Q(
        \registers[304][5] ) );
  EDFFX1 \registers_reg[304][4]  ( .D(n8256), .E(n618), .CK(clk), .Q(
        \registers[304][4] ) );
  EDFFX1 \registers_reg[304][3]  ( .D(n8173), .E(n618), .CK(clk), .Q(
        \registers[304][3] ) );
  EDFFX1 \registers_reg[304][2]  ( .D(n8160), .E(n618), .CK(clk), .Q(
        \registers[304][2] ) );
  EDFFX1 \registers_reg[304][1]  ( .D(n8104), .E(n618), .CK(clk), .Q(
        \registers[304][1] ) );
  EDFFX1 \registers_reg[304][0]  ( .D(n8044), .E(n618), .CK(clk), .Q(
        \registers[304][0] ) );
  EDFFX1 \registers_reg[300][7]  ( .D(n8434), .E(n614), .CK(clk), .Q(
        \registers[300][7] ) );
  EDFFX1 \registers_reg[300][6]  ( .D(n8376), .E(n614), .CK(clk), .Q(
        \registers[300][6] ) );
  EDFFX1 \registers_reg[300][5]  ( .D(n8318), .E(n614), .CK(clk), .Q(
        \registers[300][5] ) );
  EDFFX1 \registers_reg[300][4]  ( .D(n8260), .E(n614), .CK(clk), .Q(
        \registers[300][4] ) );
  EDFFX1 \registers_reg[300][3]  ( .D(n8174), .E(n614), .CK(clk), .Q(
        \registers[300][3] ) );
  EDFFX1 \registers_reg[300][2]  ( .D(n8158), .E(n614), .CK(clk), .Q(
        \registers[300][2] ) );
  EDFFX1 \registers_reg[300][1]  ( .D(n8102), .E(n614), .CK(clk), .Q(
        \registers[300][1] ) );
  EDFFX1 \registers_reg[300][0]  ( .D(n8045), .E(n614), .CK(clk), .Q(
        \registers[300][0] ) );
  EDFFX1 \registers_reg[296][7]  ( .D(n8428), .E(n610), .CK(clk), .Q(
        \registers[296][7] ) );
  EDFFX1 \registers_reg[296][6]  ( .D(n8370), .E(n610), .CK(clk), .Q(
        \registers[296][6] ) );
  EDFFX1 \registers_reg[296][5]  ( .D(n8312), .E(n610), .CK(clk), .Q(
        \registers[296][5] ) );
  EDFFX1 \registers_reg[296][4]  ( .D(n8254), .E(n610), .CK(clk), .Q(
        \registers[296][4] ) );
  EDFFX1 \registers_reg[296][3]  ( .D(n8167), .E(n610), .CK(clk), .Q(
        \registers[296][3] ) );
  EDFFX1 \registers_reg[296][2]  ( .D(n8159), .E(n610), .CK(clk), .Q(
        \registers[296][2] ) );
  EDFFX1 \registers_reg[296][1]  ( .D(n8103), .E(n610), .CK(clk), .Q(
        \registers[296][1] ) );
  EDFFX1 \registers_reg[296][0]  ( .D(n8043), .E(n610), .CK(clk), .Q(
        \registers[296][0] ) );
  EDFFX1 \registers_reg[292][7]  ( .D(n8429), .E(n977), .CK(clk), .Q(
        \registers[292][7] ) );
  EDFFX1 \registers_reg[292][6]  ( .D(n8371), .E(n977), .CK(clk), .Q(
        \registers[292][6] ) );
  EDFFX1 \registers_reg[292][5]  ( .D(n8313), .E(n977), .CK(clk), .Q(
        \registers[292][5] ) );
  EDFFX1 \registers_reg[292][4]  ( .D(n8255), .E(n977), .CK(clk), .Q(
        \registers[292][4] ) );
  EDFFX1 \registers_reg[292][3]  ( .D(n8200), .E(n977), .CK(clk), .Q(
        \registers[292][3] ) );
  EDFFX1 \registers_reg[292][2]  ( .D(n8160), .E(n977), .CK(clk), .Q(
        \registers[292][2] ) );
  EDFFX1 \registers_reg[292][1]  ( .D(n8104), .E(n977), .CK(clk), .Q(
        \registers[292][1] ) );
  EDFFX1 \registers_reg[292][0]  ( .D(n8044), .E(n977), .CK(clk), .Q(
        \registers[292][0] ) );
  EDFFX1 \registers_reg[288][7]  ( .D(n8425), .E(n331), .CK(clk), .Q(
        \registers[288][7] ) );
  EDFFX1 \registers_reg[288][6]  ( .D(n8367), .E(n331), .CK(clk), .Q(
        \registers[288][6] ) );
  EDFFX1 \registers_reg[288][5]  ( .D(n8309), .E(n331), .CK(clk), .Q(
        \registers[288][5] ) );
  EDFFX1 \registers_reg[288][4]  ( .D(n8251), .E(n331), .CK(clk), .Q(
        \registers[288][4] ) );
  EDFFX1 \registers_reg[288][3]  ( .D(n8201), .E(n331), .CK(clk), .Q(
        \registers[288][3] ) );
  EDFFX1 \registers_reg[288][2]  ( .D(n8158), .E(n331), .CK(clk), .Q(
        \registers[288][2] ) );
  EDFFX1 \registers_reg[288][1]  ( .D(n8102), .E(n331), .CK(clk), .Q(
        \registers[288][1] ) );
  EDFFX1 \registers_reg[288][0]  ( .D(n8045), .E(n331), .CK(clk), .Q(
        \registers[288][0] ) );
  EDFFX1 \registers_reg[284][7]  ( .D(n8428), .E(n606), .CK(clk), .Q(
        \registers[284][7] ) );
  EDFFX1 \registers_reg[284][6]  ( .D(n8370), .E(n606), .CK(clk), .Q(
        \registers[284][6] ) );
  EDFFX1 \registers_reg[284][5]  ( .D(n8312), .E(n606), .CK(clk), .Q(
        \registers[284][5] ) );
  EDFFX1 \registers_reg[284][4]  ( .D(n8254), .E(n606), .CK(clk), .Q(
        \registers[284][4] ) );
  EDFFX1 \registers_reg[284][3]  ( .D(n8202), .E(n606), .CK(clk), .Q(
        \registers[284][3] ) );
  EDFFX1 \registers_reg[284][2]  ( .D(n8159), .E(n606), .CK(clk), .Q(
        \registers[284][2] ) );
  EDFFX1 \registers_reg[284][1]  ( .D(n8103), .E(n606), .CK(clk), .Q(
        \registers[284][1] ) );
  EDFFX1 \registers_reg[284][0]  ( .D(n8043), .E(n606), .CK(clk), .Q(
        \registers[284][0] ) );
  EDFFX1 \registers_reg[280][7]  ( .D(n8429), .E(n602), .CK(clk), .Q(
        \registers[280][7] ) );
  EDFFX1 \registers_reg[280][6]  ( .D(n8371), .E(n602), .CK(clk), .Q(
        \registers[280][6] ) );
  EDFFX1 \registers_reg[280][5]  ( .D(n8313), .E(n602), .CK(clk), .Q(
        \registers[280][5] ) );
  EDFFX1 \registers_reg[280][4]  ( .D(n8255), .E(n602), .CK(clk), .Q(
        \registers[280][4] ) );
  EDFFX1 \registers_reg[280][3]  ( .D(n8200), .E(n602), .CK(clk), .Q(
        \registers[280][3] ) );
  EDFFX1 \registers_reg[280][2]  ( .D(n8160), .E(n602), .CK(clk), .Q(
        \registers[280][2] ) );
  EDFFX1 \registers_reg[280][1]  ( .D(n8104), .E(n602), .CK(clk), .Q(
        \registers[280][1] ) );
  EDFFX1 \registers_reg[280][0]  ( .D(n8044), .E(n602), .CK(clk), .Q(
        \registers[280][0] ) );
  EDFFX1 \registers_reg[276][7]  ( .D(n8426), .E(n598), .CK(clk), .Q(
        \registers[276][7] ) );
  EDFFX1 \registers_reg[276][6]  ( .D(n8368), .E(n598), .CK(clk), .Q(
        \registers[276][6] ) );
  EDFFX1 \registers_reg[276][5]  ( .D(n8310), .E(n598), .CK(clk), .Q(
        \registers[276][5] ) );
  EDFFX1 \registers_reg[276][4]  ( .D(n8252), .E(n598), .CK(clk), .Q(
        \registers[276][4] ) );
  EDFFX1 \registers_reg[276][3]  ( .D(n8201), .E(n598), .CK(clk), .Q(
        \registers[276][3] ) );
  EDFFX1 \registers_reg[276][2]  ( .D(n8158), .E(n598), .CK(clk), .Q(
        \registers[276][2] ) );
  EDFFX1 \registers_reg[276][1]  ( .D(n8102), .E(n598), .CK(clk), .Q(
        \registers[276][1] ) );
  EDFFX1 \registers_reg[276][0]  ( .D(n8045), .E(n598), .CK(clk), .Q(
        \registers[276][0] ) );
  EDFFX1 \registers_reg[272][7]  ( .D(n8428), .E(n594), .CK(clk), .Q(
        \registers[272][7] ) );
  EDFFX1 \registers_reg[272][6]  ( .D(n8370), .E(n594), .CK(clk), .Q(
        \registers[272][6] ) );
  EDFFX1 \registers_reg[272][5]  ( .D(n8312), .E(n594), .CK(clk), .Q(
        \registers[272][5] ) );
  EDFFX1 \registers_reg[272][4]  ( .D(n8254), .E(n594), .CK(clk), .Q(
        \registers[272][4] ) );
  EDFFX1 \registers_reg[272][3]  ( .D(n8202), .E(n594), .CK(clk), .Q(
        \registers[272][3] ) );
  EDFFX1 \registers_reg[272][2]  ( .D(n8159), .E(n594), .CK(clk), .Q(
        \registers[272][2] ) );
  EDFFX1 \registers_reg[272][1]  ( .D(n8103), .E(n594), .CK(clk), .Q(
        \registers[272][1] ) );
  EDFFX1 \registers_reg[272][0]  ( .D(n8043), .E(n594), .CK(clk), .Q(
        \registers[272][0] ) );
  EDFFX1 \registers_reg[268][7]  ( .D(n8429), .E(n590), .CK(clk), .Q(
        \registers[268][7] ) );
  EDFFX1 \registers_reg[268][6]  ( .D(n8371), .E(n590), .CK(clk), .Q(
        \registers[268][6] ) );
  EDFFX1 \registers_reg[268][5]  ( .D(n8313), .E(n590), .CK(clk), .Q(
        \registers[268][5] ) );
  EDFFX1 \registers_reg[268][4]  ( .D(n8255), .E(n590), .CK(clk), .Q(
        \registers[268][4] ) );
  EDFFX1 \registers_reg[268][3]  ( .D(n8200), .E(n590), .CK(clk), .Q(
        \registers[268][3] ) );
  EDFFX1 \registers_reg[268][2]  ( .D(n8157), .E(n590), .CK(clk), .Q(
        \registers[268][2] ) );
  EDFFX1 \registers_reg[268][1]  ( .D(n8101), .E(n590), .CK(clk), .Q(
        \registers[268][1] ) );
  EDFFX1 \registers_reg[268][0]  ( .D(n8041), .E(n590), .CK(clk), .Q(
        \registers[268][0] ) );
  EDFFX1 \registers_reg[264][7]  ( .D(n8427), .E(n586), .CK(clk), .Q(
        \registers[264][7] ) );
  EDFFX1 \registers_reg[264][6]  ( .D(n8369), .E(n586), .CK(clk), .Q(
        \registers[264][6] ) );
  EDFFX1 \registers_reg[264][5]  ( .D(n8311), .E(n586), .CK(clk), .Q(
        \registers[264][5] ) );
  EDFFX1 \registers_reg[264][4]  ( .D(n8253), .E(n586), .CK(clk), .Q(
        \registers[264][4] ) );
  EDFFX1 \registers_reg[264][3]  ( .D(n8201), .E(n586), .CK(clk), .Q(
        \registers[264][3] ) );
  EDFFX1 \registers_reg[264][2]  ( .D(n8155), .E(n586), .CK(clk), .Q(
        \registers[264][2] ) );
  EDFFX1 \registers_reg[264][1]  ( .D(n8099), .E(n586), .CK(clk), .Q(
        \registers[264][1] ) );
  EDFFX1 \registers_reg[264][0]  ( .D(n8042), .E(n586), .CK(clk), .Q(
        \registers[264][0] ) );
  EDFFX1 \registers_reg[260][7]  ( .D(n8428), .E(n970), .CK(clk), .Q(
        \registers[260][7] ) );
  EDFFX1 \registers_reg[260][6]  ( .D(n8370), .E(n970), .CK(clk), .Q(
        \registers[260][6] ) );
  EDFFX1 \registers_reg[260][5]  ( .D(n8312), .E(n970), .CK(clk), .Q(
        \registers[260][5] ) );
  EDFFX1 \registers_reg[260][4]  ( .D(n8254), .E(n970), .CK(clk), .Q(
        \registers[260][4] ) );
  EDFFX1 \registers_reg[260][3]  ( .D(n8202), .E(n970), .CK(clk), .Q(
        \registers[260][3] ) );
  EDFFX1 \registers_reg[260][2]  ( .D(n8156), .E(n970), .CK(clk), .Q(
        \registers[260][2] ) );
  EDFFX1 \registers_reg[260][1]  ( .D(n8100), .E(n970), .CK(clk), .Q(
        \registers[260][1] ) );
  EDFFX1 \registers_reg[260][0]  ( .D(n8040), .E(n970), .CK(clk), .Q(
        \registers[260][0] ) );
  EDFFX1 \registers_reg[256][7]  ( .D(n8411), .E(n330), .CK(clk), .Q(
        \registers[256][7] ) );
  EDFFX1 \registers_reg[256][6]  ( .D(n8353), .E(n330), .CK(clk), .Q(
        \registers[256][6] ) );
  EDFFX1 \registers_reg[256][5]  ( .D(n8295), .E(n330), .CK(clk), .Q(
        \registers[256][5] ) );
  EDFFX1 \registers_reg[256][4]  ( .D(n8237), .E(n330), .CK(clk), .Q(
        \registers[256][4] ) );
  EDFFX1 \registers_reg[256][3]  ( .D(n8188), .E(n330), .CK(clk), .Q(
        \registers[256][3] ) );
  EDFFX1 \registers_reg[256][2]  ( .D(n8143), .E(n330), .CK(clk), .Q(
        \registers[256][2] ) );
  EDFFX1 \registers_reg[256][1]  ( .D(n8087), .E(n330), .CK(clk), .Q(
        \registers[256][1] ) );
  EDFFX1 \registers_reg[256][0]  ( .D(n8043), .E(n330), .CK(clk), .Q(
        \registers[256][0] ) );
  EDFFX1 \registers_reg[252][7]  ( .D(n8412), .E(n582), .CK(clk), .Q(
        \registers[252][7] ) );
  EDFFX1 \registers_reg[252][6]  ( .D(n8354), .E(n582), .CK(clk), .Q(
        \registers[252][6] ) );
  EDFFX1 \registers_reg[252][5]  ( .D(n8296), .E(n582), .CK(clk), .Q(
        \registers[252][5] ) );
  EDFFX1 \registers_reg[252][4]  ( .D(n8238), .E(n582), .CK(clk), .Q(
        \registers[252][4] ) );
  EDFFX1 \registers_reg[252][3]  ( .D(n8189), .E(n582), .CK(clk), .Q(
        \registers[252][3] ) );
  EDFFX1 \registers_reg[252][2]  ( .D(n8141), .E(n582), .CK(clk), .Q(
        \registers[252][2] ) );
  EDFFX1 \registers_reg[252][1]  ( .D(n8085), .E(n582), .CK(clk), .Q(
        \registers[252][1] ) );
  EDFFX1 \registers_reg[252][0]  ( .D(n8027), .E(n582), .CK(clk), .Q(
        \registers[252][0] ) );
  EDFFX1 \registers_reg[248][7]  ( .D(n8410), .E(n578), .CK(clk), .Q(
        \registers[248][7] ) );
  EDFFX1 \registers_reg[248][6]  ( .D(n8352), .E(n578), .CK(clk), .Q(
        \registers[248][6] ) );
  EDFFX1 \registers_reg[248][5]  ( .D(n8294), .E(n578), .CK(clk), .Q(
        \registers[248][5] ) );
  EDFFX1 \registers_reg[248][4]  ( .D(n8236), .E(n578), .CK(clk), .Q(
        \registers[248][4] ) );
  EDFFX1 \registers_reg[248][3]  ( .D(n8190), .E(n578), .CK(clk), .Q(
        \registers[248][3] ) );
  EDFFX1 \registers_reg[248][2]  ( .D(n8142), .E(n578), .CK(clk), .Q(
        \registers[248][2] ) );
  EDFFX1 \registers_reg[248][1]  ( .D(n8086), .E(n578), .CK(clk), .Q(
        \registers[248][1] ) );
  EDFFX1 \registers_reg[248][0]  ( .D(n8025), .E(n578), .CK(clk), .Q(
        \registers[248][0] ) );
  EDFFX1 \registers_reg[244][7]  ( .D(n8411), .E(n574), .CK(clk), .Q(
        \registers[244][7] ) );
  EDFFX1 \registers_reg[244][6]  ( .D(n8353), .E(n574), .CK(clk), .Q(
        \registers[244][6] ) );
  EDFFX1 \registers_reg[244][5]  ( .D(n8295), .E(n574), .CK(clk), .Q(
        \registers[244][5] ) );
  EDFFX1 \registers_reg[244][4]  ( .D(n8237), .E(n574), .CK(clk), .Q(
        \registers[244][4] ) );
  EDFFX1 \registers_reg[244][3]  ( .D(n8188), .E(n574), .CK(clk), .Q(
        \registers[244][3] ) );
  EDFFX1 \registers_reg[244][2]  ( .D(n8143), .E(n574), .CK(clk), .Q(
        \registers[244][2] ) );
  EDFFX1 \registers_reg[244][1]  ( .D(n8087), .E(n574), .CK(clk), .Q(
        \registers[244][1] ) );
  EDFFX1 \registers_reg[244][0]  ( .D(n8026), .E(n574), .CK(clk), .Q(
        \registers[244][0] ) );
  EDFFX1 \registers_reg[240][7]  ( .D(n8412), .E(n570), .CK(clk), .Q(
        \registers[240][7] ) );
  EDFFX1 \registers_reg[240][6]  ( .D(n8354), .E(n570), .CK(clk), .Q(
        \registers[240][6] ) );
  EDFFX1 \registers_reg[240][5]  ( .D(n8296), .E(n570), .CK(clk), .Q(
        \registers[240][5] ) );
  EDFFX1 \registers_reg[240][4]  ( .D(n8238), .E(n570), .CK(clk), .Q(
        \registers[240][4] ) );
  EDFFX1 \registers_reg[240][3]  ( .D(n8189), .E(n570), .CK(clk), .Q(
        \registers[240][3] ) );
  EDFFX1 \registers_reg[240][2]  ( .D(n8141), .E(n570), .CK(clk), .Q(
        \registers[240][2] ) );
  EDFFX1 \registers_reg[240][1]  ( .D(n8085), .E(n570), .CK(clk), .Q(
        \registers[240][1] ) );
  EDFFX1 \registers_reg[240][0]  ( .D(n8027), .E(n570), .CK(clk), .Q(
        \registers[240][0] ) );
  EDFFX1 \registers_reg[236][7]  ( .D(n8410), .E(n566), .CK(clk), .Q(
        \registers[236][7] ) );
  EDFFX1 \registers_reg[236][6]  ( .D(n8352), .E(n566), .CK(clk), .Q(
        \registers[236][6] ) );
  EDFFX1 \registers_reg[236][5]  ( .D(n8294), .E(n566), .CK(clk), .Q(
        \registers[236][5] ) );
  EDFFX1 \registers_reg[236][4]  ( .D(n8236), .E(n566), .CK(clk), .Q(
        \registers[236][4] ) );
  EDFFX1 \registers_reg[236][3]  ( .D(n8190), .E(n566), .CK(clk), .Q(
        \registers[236][3] ) );
  EDFFX1 \registers_reg[236][2]  ( .D(n8142), .E(n566), .CK(clk), .Q(
        \registers[236][2] ) );
  EDFFX1 \registers_reg[236][1]  ( .D(n8086), .E(n566), .CK(clk), .Q(
        \registers[236][1] ) );
  EDFFX1 \registers_reg[236][0]  ( .D(n8025), .E(n566), .CK(clk), .Q(
        \registers[236][0] ) );
  EDFFX1 \registers_reg[232][7]  ( .D(n8411), .E(n562), .CK(clk), .Q(
        \registers[232][7] ) );
  EDFFX1 \registers_reg[232][6]  ( .D(n8353), .E(n562), .CK(clk), .Q(
        \registers[232][6] ) );
  EDFFX1 \registers_reg[232][5]  ( .D(n8295), .E(n562), .CK(clk), .Q(
        \registers[232][5] ) );
  EDFFX1 \registers_reg[232][4]  ( .D(n8237), .E(n562), .CK(clk), .Q(
        \registers[232][4] ) );
  EDFFX1 \registers_reg[232][3]  ( .D(n8185), .E(n562), .CK(clk), .Q(
        \registers[232][3] ) );
  EDFFX1 \registers_reg[232][2]  ( .D(n8143), .E(n562), .CK(clk), .Q(
        \registers[232][2] ) );
  EDFFX1 \registers_reg[232][1]  ( .D(n8087), .E(n562), .CK(clk), .Q(
        \registers[232][1] ) );
  EDFFX1 \registers_reg[232][0]  ( .D(n8026), .E(n562), .CK(clk), .Q(
        \registers[232][0] ) );
  EDFFX1 \registers_reg[228][7]  ( .D(n8412), .E(n1030), .CK(clk), .Q(
        \registers[228][7] ) );
  EDFFX1 \registers_reg[228][6]  ( .D(n8354), .E(n1030), .CK(clk), .Q(
        \registers[228][6] ) );
  EDFFX1 \registers_reg[228][5]  ( .D(n8296), .E(n1030), .CK(clk), .Q(
        \registers[228][5] ) );
  EDFFX1 \registers_reg[228][4]  ( .D(n8238), .E(n1030), .CK(clk), .Q(
        \registers[228][4] ) );
  EDFFX1 \registers_reg[228][3]  ( .D(n8186), .E(n1030), .CK(clk), .Q(
        \registers[228][3] ) );
  EDFFX1 \registers_reg[228][2]  ( .D(n8141), .E(n1030), .CK(clk), .Q(
        \registers[228][2] ) );
  EDFFX1 \registers_reg[228][1]  ( .D(n8085), .E(n1030), .CK(clk), .Q(
        \registers[228][1] ) );
  EDFFX1 \registers_reg[228][0]  ( .D(n8027), .E(n1030), .CK(clk), .Q(
        \registers[228][0] ) );
  EDFFX1 \registers_reg[224][7]  ( .D(n8410), .E(n390), .CK(clk), .Q(
        \registers[224][7] ) );
  EDFFX1 \registers_reg[224][6]  ( .D(n8352), .E(n390), .CK(clk), .Q(
        \registers[224][6] ) );
  EDFFX1 \registers_reg[224][5]  ( .D(n8294), .E(n390), .CK(clk), .Q(
        \registers[224][5] ) );
  EDFFX1 \registers_reg[224][4]  ( .D(n8236), .E(n390), .CK(clk), .Q(
        \registers[224][4] ) );
  EDFFX1 \registers_reg[224][3]  ( .D(n8187), .E(n390), .CK(clk), .Q(
        \registers[224][3] ) );
  EDFFX1 \registers_reg[224][2]  ( .D(n8142), .E(n390), .CK(clk), .Q(
        \registers[224][2] ) );
  EDFFX1 \registers_reg[224][1]  ( .D(n8086), .E(n390), .CK(clk), .Q(
        \registers[224][1] ) );
  EDFFX1 \registers_reg[224][0]  ( .D(n8025), .E(n390), .CK(clk), .Q(
        \registers[224][0] ) );
  EDFFX1 \registers_reg[220][7]  ( .D(n8411), .E(n558), .CK(clk), .Q(
        \registers[220][7] ) );
  EDFFX1 \registers_reg[220][6]  ( .D(n8353), .E(n558), .CK(clk), .Q(
        \registers[220][6] ) );
  EDFFX1 \registers_reg[220][5]  ( .D(n8295), .E(n558), .CK(clk), .Q(
        \registers[220][5] ) );
  EDFFX1 \registers_reg[220][4]  ( .D(n8237), .E(n558), .CK(clk), .Q(
        \registers[220][4] ) );
  EDFFX1 \registers_reg[220][3]  ( .D(n8185), .E(n558), .CK(clk), .Q(
        \registers[220][3] ) );
  EDFFX1 \registers_reg[220][2]  ( .D(n8143), .E(n558), .CK(clk), .Q(
        \registers[220][2] ) );
  EDFFX1 \registers_reg[220][1]  ( .D(n8087), .E(n558), .CK(clk), .Q(
        \registers[220][1] ) );
  EDFFX1 \registers_reg[220][0]  ( .D(n8026), .E(n558), .CK(clk), .Q(
        \registers[220][0] ) );
  EDFFX1 \registers_reg[216][7]  ( .D(n8412), .E(n554), .CK(clk), .Q(
        \registers[216][7] ) );
  EDFFX1 \registers_reg[216][6]  ( .D(n8354), .E(n554), .CK(clk), .Q(
        \registers[216][6] ) );
  EDFFX1 \registers_reg[216][5]  ( .D(n8296), .E(n554), .CK(clk), .Q(
        \registers[216][5] ) );
  EDFFX1 \registers_reg[216][4]  ( .D(n8238), .E(n554), .CK(clk), .Q(
        \registers[216][4] ) );
  EDFFX1 \registers_reg[216][3]  ( .D(n8186), .E(n554), .CK(clk), .Q(
        \registers[216][3] ) );
  EDFFX1 \registers_reg[216][2]  ( .D(n8138), .E(n554), .CK(clk), .Q(
        \registers[216][2] ) );
  EDFFX1 \registers_reg[216][1]  ( .D(n8082), .E(n554), .CK(clk), .Q(
        \registers[216][1] ) );
  EDFFX1 \registers_reg[216][0]  ( .D(n8024), .E(n554), .CK(clk), .Q(
        \registers[216][0] ) );
  EDFFX1 \registers_reg[212][7]  ( .D(n8410), .E(n550), .CK(clk), .Q(
        \registers[212][7] ) );
  EDFFX1 \registers_reg[212][6]  ( .D(n8352), .E(n550), .CK(clk), .Q(
        \registers[212][6] ) );
  EDFFX1 \registers_reg[212][5]  ( .D(n8294), .E(n550), .CK(clk), .Q(
        \registers[212][5] ) );
  EDFFX1 \registers_reg[212][4]  ( .D(n8236), .E(n550), .CK(clk), .Q(
        \registers[212][4] ) );
  EDFFX1 \registers_reg[212][3]  ( .D(n8187), .E(n550), .CK(clk), .Q(
        \registers[212][3] ) );
  EDFFX1 \registers_reg[212][2]  ( .D(n8139), .E(n550), .CK(clk), .Q(
        \registers[212][2] ) );
  EDFFX1 \registers_reg[212][1]  ( .D(n8083), .E(n550), .CK(clk), .Q(
        \registers[212][1] ) );
  EDFFX1 \registers_reg[212][0]  ( .D(n8022), .E(n550), .CK(clk), .Q(
        \registers[212][0] ) );
  EDFFX1 \registers_reg[208][7]  ( .D(n8411), .E(n546), .CK(clk), .Q(
        \registers[208][7] ) );
  EDFFX1 \registers_reg[208][6]  ( .D(n8353), .E(n546), .CK(clk), .Q(
        \registers[208][6] ) );
  EDFFX1 \registers_reg[208][5]  ( .D(n8295), .E(n546), .CK(clk), .Q(
        \registers[208][5] ) );
  EDFFX1 \registers_reg[208][4]  ( .D(n8237), .E(n546), .CK(clk), .Q(
        \registers[208][4] ) );
  EDFFX1 \registers_reg[208][3]  ( .D(n8185), .E(n546), .CK(clk), .Q(
        \registers[208][3] ) );
  EDFFX1 \registers_reg[208][2]  ( .D(n8140), .E(n546), .CK(clk), .Q(
        \registers[208][2] ) );
  EDFFX1 \registers_reg[208][1]  ( .D(n8084), .E(n546), .CK(clk), .Q(
        \registers[208][1] ) );
  EDFFX1 \registers_reg[208][0]  ( .D(n8023), .E(n546), .CK(clk), .Q(
        \registers[208][0] ) );
  EDFFX1 \registers_reg[204][7]  ( .D(n8407), .E(n542), .CK(clk), .Q(
        \registers[204][7] ) );
  EDFFX1 \registers_reg[204][6]  ( .D(n8349), .E(n542), .CK(clk), .Q(
        \registers[204][6] ) );
  EDFFX1 \registers_reg[204][5]  ( .D(n8291), .E(n542), .CK(clk), .Q(
        \registers[204][5] ) );
  EDFFX1 \registers_reg[204][4]  ( .D(n8233), .E(n542), .CK(clk), .Q(
        \registers[204][4] ) );
  EDFFX1 \registers_reg[204][3]  ( .D(n8186), .E(n542), .CK(clk), .Q(
        \registers[204][3] ) );
  EDFFX1 \registers_reg[204][2]  ( .D(n8138), .E(n542), .CK(clk), .Q(
        \registers[204][2] ) );
  EDFFX1 \registers_reg[204][1]  ( .D(n8082), .E(n542), .CK(clk), .Q(
        \registers[204][1] ) );
  EDFFX1 \registers_reg[204][0]  ( .D(n8024), .E(n542), .CK(clk), .Q(
        \registers[204][0] ) );
  EDFFX1 \registers_reg[200][7]  ( .D(n8408), .E(n538), .CK(clk), .Q(
        \registers[200][7] ) );
  EDFFX1 \registers_reg[200][6]  ( .D(n8350), .E(n538), .CK(clk), .Q(
        \registers[200][6] ) );
  EDFFX1 \registers_reg[200][5]  ( .D(n8292), .E(n538), .CK(clk), .Q(
        \registers[200][5] ) );
  EDFFX1 \registers_reg[200][4]  ( .D(n8234), .E(n538), .CK(clk), .Q(
        \registers[200][4] ) );
  EDFFX1 \registers_reg[200][3]  ( .D(n8187), .E(n538), .CK(clk), .Q(
        \registers[200][3] ) );
  EDFFX1 \registers_reg[200][2]  ( .D(n8139), .E(n538), .CK(clk), .Q(
        \registers[200][2] ) );
  EDFFX1 \registers_reg[200][1]  ( .D(n8083), .E(n538), .CK(clk), .Q(
        \registers[200][1] ) );
  EDFFX1 \registers_reg[200][0]  ( .D(n8022), .E(n538), .CK(clk), .Q(
        \registers[200][0] ) );
  EDFFX1 \registers_reg[196][7]  ( .D(n8409), .E(n1026), .CK(clk), .Q(
        \registers[196][7] ) );
  EDFFX1 \registers_reg[196][6]  ( .D(n8351), .E(n1026), .CK(clk), .Q(
        \registers[196][6] ) );
  EDFFX1 \registers_reg[196][5]  ( .D(n8293), .E(n1026), .CK(clk), .Q(
        \registers[196][5] ) );
  EDFFX1 \registers_reg[196][4]  ( .D(n8235), .E(n1026), .CK(clk), .Q(
        \registers[196][4] ) );
  EDFFX1 \registers_reg[196][3]  ( .D(n8185), .E(n1026), .CK(clk), .Q(
        \registers[196][3] ) );
  EDFFX1 \registers_reg[196][2]  ( .D(n8140), .E(n1026), .CK(clk), .Q(
        \registers[196][2] ) );
  EDFFX1 \registers_reg[196][1]  ( .D(n8084), .E(n1026), .CK(clk), .Q(
        \registers[196][1] ) );
  EDFFX1 \registers_reg[196][0]  ( .D(n8023), .E(n1026), .CK(clk), .Q(
        \registers[196][0] ) );
  EDFFX1 \registers_reg[192][7]  ( .D(n8408), .E(n389), .CK(clk), .Q(
        \registers[192][7] ) );
  EDFFX1 \registers_reg[192][6]  ( .D(n8350), .E(n389), .CK(clk), .Q(
        \registers[192][6] ) );
  EDFFX1 \registers_reg[192][5]  ( .D(n8292), .E(n389), .CK(clk), .Q(
        \registers[192][5] ) );
  EDFFX1 \registers_reg[192][4]  ( .D(n8234), .E(n389), .CK(clk), .Q(
        \registers[192][4] ) );
  EDFFX1 \registers_reg[192][3]  ( .D(n8187), .E(n389), .CK(clk), .Q(
        \registers[192][3] ) );
  EDFFX1 \registers_reg[192][2]  ( .D(n8139), .E(n389), .CK(clk), .Q(
        \registers[192][2] ) );
  EDFFX1 \registers_reg[192][1]  ( .D(n8083), .E(n389), .CK(clk), .Q(
        \registers[192][1] ) );
  EDFFX1 \registers_reg[192][0]  ( .D(n8024), .E(n389), .CK(clk), .Q(
        \registers[192][0] ) );
  EDFFX1 \registers_reg[188][7]  ( .D(n8409), .E(n534), .CK(clk), .Q(
        \registers[188][7] ) );
  EDFFX1 \registers_reg[188][6]  ( .D(n8351), .E(n534), .CK(clk), .Q(
        \registers[188][6] ) );
  EDFFX1 \registers_reg[188][5]  ( .D(n8293), .E(n534), .CK(clk), .Q(
        \registers[188][5] ) );
  EDFFX1 \registers_reg[188][4]  ( .D(n8235), .E(n534), .CK(clk), .Q(
        \registers[188][4] ) );
  EDFFX1 \registers_reg[188][3]  ( .D(n8185), .E(n534), .CK(clk), .Q(
        \registers[188][3] ) );
  EDFFX1 \registers_reg[188][2]  ( .D(n8140), .E(n534), .CK(clk), .Q(
        \registers[188][2] ) );
  EDFFX1 \registers_reg[188][1]  ( .D(n8084), .E(n534), .CK(clk), .Q(
        \registers[188][1] ) );
  EDFFX1 \registers_reg[188][0]  ( .D(n8023), .E(n534), .CK(clk), .Q(
        \registers[188][0] ) );
  EDFFX1 \registers_reg[184][7]  ( .D(n8407), .E(n530), .CK(clk), .Q(
        \registers[184][7] ) );
  EDFFX1 \registers_reg[184][6]  ( .D(n8349), .E(n530), .CK(clk), .Q(
        \registers[184][6] ) );
  EDFFX1 \registers_reg[184][5]  ( .D(n8291), .E(n530), .CK(clk), .Q(
        \registers[184][5] ) );
  EDFFX1 \registers_reg[184][4]  ( .D(n8233), .E(n530), .CK(clk), .Q(
        \registers[184][4] ) );
  EDFFX1 \registers_reg[184][3]  ( .D(n8186), .E(n530), .CK(clk), .Q(
        \registers[184][3] ) );
  EDFFX1 \registers_reg[184][2]  ( .D(n8138), .E(n530), .CK(clk), .Q(
        \registers[184][2] ) );
  EDFFX1 \registers_reg[184][1]  ( .D(n8082), .E(n530), .CK(clk), .Q(
        \registers[184][1] ) );
  EDFFX1 \registers_reg[184][0]  ( .D(n8024), .E(n530), .CK(clk), .Q(
        \registers[184][0] ) );
  EDFFX1 \registers_reg[180][7]  ( .D(n8408), .E(n526), .CK(clk), .Q(
        \registers[180][7] ) );
  EDFFX1 \registers_reg[180][6]  ( .D(n8350), .E(n526), .CK(clk), .Q(
        \registers[180][6] ) );
  EDFFX1 \registers_reg[180][5]  ( .D(n8292), .E(n526), .CK(clk), .Q(
        \registers[180][5] ) );
  EDFFX1 \registers_reg[180][4]  ( .D(n8234), .E(n526), .CK(clk), .Q(
        \registers[180][4] ) );
  EDFFX1 \registers_reg[180][3]  ( .D(n8187), .E(n526), .CK(clk), .Q(
        \registers[180][3] ) );
  EDFFX1 \registers_reg[180][2]  ( .D(n8139), .E(n526), .CK(clk), .Q(
        \registers[180][2] ) );
  EDFFX1 \registers_reg[180][1]  ( .D(n8083), .E(n526), .CK(clk), .Q(
        \registers[180][1] ) );
  EDFFX1 \registers_reg[180][0]  ( .D(n8022), .E(n526), .CK(clk), .Q(
        \registers[180][0] ) );
  EDFFX1 \registers_reg[176][7]  ( .D(n8409), .E(n522), .CK(clk), .Q(
        \registers[176][7] ) );
  EDFFX1 \registers_reg[176][6]  ( .D(n8351), .E(n522), .CK(clk), .Q(
        \registers[176][6] ) );
  EDFFX1 \registers_reg[176][5]  ( .D(n8293), .E(n522), .CK(clk), .Q(
        \registers[176][5] ) );
  EDFFX1 \registers_reg[176][4]  ( .D(n8235), .E(n522), .CK(clk), .Q(
        \registers[176][4] ) );
  EDFFX1 \registers_reg[176][3]  ( .D(n8185), .E(n522), .CK(clk), .Q(
        \registers[176][3] ) );
  EDFFX1 \registers_reg[176][2]  ( .D(n8140), .E(n522), .CK(clk), .Q(
        \registers[176][2] ) );
  EDFFX1 \registers_reg[176][1]  ( .D(n8084), .E(n522), .CK(clk), .Q(
        \registers[176][1] ) );
  EDFFX1 \registers_reg[176][0]  ( .D(n8023), .E(n522), .CK(clk), .Q(
        \registers[176][0] ) );
  EDFFX1 \registers_reg[172][7]  ( .D(n8407), .E(n518), .CK(clk), .Q(
        \registers[172][7] ) );
  EDFFX1 \registers_reg[172][6]  ( .D(n8349), .E(n518), .CK(clk), .Q(
        \registers[172][6] ) );
  EDFFX1 \registers_reg[172][5]  ( .D(n8291), .E(n518), .CK(clk), .Q(
        \registers[172][5] ) );
  EDFFX1 \registers_reg[172][4]  ( .D(n8233), .E(n518), .CK(clk), .Q(
        \registers[172][4] ) );
  EDFFX1 \registers_reg[172][3]  ( .D(n8183), .E(n518), .CK(clk), .Q(
        \registers[172][3] ) );
  EDFFX1 \registers_reg[172][2]  ( .D(n8138), .E(n518), .CK(clk), .Q(
        \registers[172][2] ) );
  EDFFX1 \registers_reg[172][1]  ( .D(n8082), .E(n518), .CK(clk), .Q(
        \registers[172][1] ) );
  EDFFX1 \registers_reg[172][0]  ( .D(n8024), .E(n518), .CK(clk), .Q(
        \registers[172][0] ) );
  EDFFX1 \registers_reg[168][7]  ( .D(n8408), .E(n514), .CK(clk), .Q(
        \registers[168][7] ) );
  EDFFX1 \registers_reg[168][6]  ( .D(n8350), .E(n514), .CK(clk), .Q(
        \registers[168][6] ) );
  EDFFX1 \registers_reg[168][5]  ( .D(n8292), .E(n514), .CK(clk), .Q(
        \registers[168][5] ) );
  EDFFX1 \registers_reg[168][4]  ( .D(n8234), .E(n514), .CK(clk), .Q(
        \registers[168][4] ) );
  EDFFX1 \registers_reg[168][3]  ( .D(n8184), .E(n514), .CK(clk), .Q(
        \registers[168][3] ) );
  EDFFX1 \registers_reg[168][2]  ( .D(n8136), .E(n514), .CK(clk), .Q(
        \registers[168][2] ) );
  EDFFX1 \registers_reg[168][1]  ( .D(n8080), .E(n514), .CK(clk), .Q(
        \registers[168][1] ) );
  EDFFX1 \registers_reg[168][0]  ( .D(n8019), .E(n514), .CK(clk), .Q(
        \registers[168][0] ) );
  EDFFX1 \registers_reg[164][7]  ( .D(n8409), .E(n1022), .CK(clk), .Q(
        \registers[164][7] ) );
  EDFFX1 \registers_reg[164][6]  ( .D(n8351), .E(n1022), .CK(clk), .Q(
        \registers[164][6] ) );
  EDFFX1 \registers_reg[164][5]  ( .D(n8293), .E(n1022), .CK(clk), .Q(
        \registers[164][5] ) );
  EDFFX1 \registers_reg[164][4]  ( .D(n8235), .E(n1022), .CK(clk), .Q(
        \registers[164][4] ) );
  EDFFX1 \registers_reg[164][3]  ( .D(n8182), .E(n1022), .CK(clk), .Q(
        \registers[164][3] ) );
  EDFFX1 \registers_reg[164][2]  ( .D(n8137), .E(n1022), .CK(clk), .Q(
        \registers[164][2] ) );
  EDFFX1 \registers_reg[164][1]  ( .D(n8081), .E(n1022), .CK(clk), .Q(
        \registers[164][1] ) );
  EDFFX1 \registers_reg[164][0]  ( .D(n8020), .E(n1022), .CK(clk), .Q(
        \registers[164][0] ) );
  EDFFX1 \registers_reg[160][7]  ( .D(n8407), .E(n388), .CK(clk), .Q(
        \registers[160][7] ) );
  EDFFX1 \registers_reg[160][6]  ( .D(n8349), .E(n388), .CK(clk), .Q(
        \registers[160][6] ) );
  EDFFX1 \registers_reg[160][5]  ( .D(n8291), .E(n388), .CK(clk), .Q(
        \registers[160][5] ) );
  EDFFX1 \registers_reg[160][4]  ( .D(n8233), .E(n388), .CK(clk), .Q(
        \registers[160][4] ) );
  EDFFX1 \registers_reg[160][3]  ( .D(n8183), .E(n388), .CK(clk), .Q(
        \registers[160][3] ) );
  EDFFX1 \registers_reg[160][2]  ( .D(n8135), .E(n388), .CK(clk), .Q(
        \registers[160][2] ) );
  EDFFX1 \registers_reg[160][1]  ( .D(n8079), .E(n388), .CK(clk), .Q(
        \registers[160][1] ) );
  EDFFX1 \registers_reg[160][0]  ( .D(n8021), .E(n388), .CK(clk), .Q(
        \registers[160][0] ) );
  EDFFX1 \registers_reg[156][7]  ( .D(n8406), .E(n510), .CK(clk), .Q(
        \registers[156][7] ) );
  EDFFX1 \registers_reg[156][6]  ( .D(n8348), .E(n510), .CK(clk), .Q(
        \registers[156][6] ) );
  EDFFX1 \registers_reg[156][5]  ( .D(n8290), .E(n510), .CK(clk), .Q(
        \registers[156][5] ) );
  EDFFX1 \registers_reg[156][4]  ( .D(n8232), .E(n510), .CK(clk), .Q(
        \registers[156][4] ) );
  EDFFX1 \registers_reg[156][3]  ( .D(n8184), .E(n510), .CK(clk), .Q(
        \registers[156][3] ) );
  EDFFX1 \registers_reg[156][2]  ( .D(n8136), .E(n510), .CK(clk), .Q(
        \registers[156][2] ) );
  EDFFX1 \registers_reg[156][1]  ( .D(n8080), .E(n510), .CK(clk), .Q(
        \registers[156][1] ) );
  EDFFX1 \registers_reg[156][0]  ( .D(n8019), .E(n510), .CK(clk), .Q(
        \registers[156][0] ) );
  EDFFX1 \registers_reg[152][7]  ( .D(n8404), .E(n506), .CK(clk), .Q(
        \registers[152][7] ) );
  EDFFX1 \registers_reg[152][6]  ( .D(n8346), .E(n506), .CK(clk), .Q(
        \registers[152][6] ) );
  EDFFX1 \registers_reg[152][5]  ( .D(n8288), .E(n506), .CK(clk), .Q(
        \registers[152][5] ) );
  EDFFX1 \registers_reg[152][4]  ( .D(n8230), .E(n506), .CK(clk), .Q(
        \registers[152][4] ) );
  EDFFX1 \registers_reg[152][3]  ( .D(n8182), .E(n506), .CK(clk), .Q(
        \registers[152][3] ) );
  EDFFX1 \registers_reg[152][2]  ( .D(n8137), .E(n506), .CK(clk), .Q(
        \registers[152][2] ) );
  EDFFX1 \registers_reg[152][1]  ( .D(n8081), .E(n506), .CK(clk), .Q(
        \registers[152][1] ) );
  EDFFX1 \registers_reg[152][0]  ( .D(n8020), .E(n506), .CK(clk), .Q(
        \registers[152][0] ) );
  EDFFX1 \registers_reg[148][7]  ( .D(n8405), .E(n502), .CK(clk), .Q(
        \registers[148][7] ) );
  EDFFX1 \registers_reg[148][6]  ( .D(n8347), .E(n502), .CK(clk), .Q(
        \registers[148][6] ) );
  EDFFX1 \registers_reg[148][5]  ( .D(n8289), .E(n502), .CK(clk), .Q(
        \registers[148][5] ) );
  EDFFX1 \registers_reg[148][4]  ( .D(n8231), .E(n502), .CK(clk), .Q(
        \registers[148][4] ) );
  EDFFX1 \registers_reg[148][3]  ( .D(n8183), .E(n502), .CK(clk), .Q(
        \registers[148][3] ) );
  EDFFX1 \registers_reg[148][2]  ( .D(n8135), .E(n502), .CK(clk), .Q(
        \registers[148][2] ) );
  EDFFX1 \registers_reg[148][1]  ( .D(n8079), .E(n502), .CK(clk), .Q(
        \registers[148][1] ) );
  EDFFX1 \registers_reg[148][0]  ( .D(n8021), .E(n502), .CK(clk), .Q(
        \registers[148][0] ) );
  EDFFX1 \registers_reg[144][7]  ( .D(n8406), .E(n498), .CK(clk), .Q(
        \registers[144][7] ) );
  EDFFX1 \registers_reg[144][6]  ( .D(n8348), .E(n498), .CK(clk), .Q(
        \registers[144][6] ) );
  EDFFX1 \registers_reg[144][5]  ( .D(n8290), .E(n498), .CK(clk), .Q(
        \registers[144][5] ) );
  EDFFX1 \registers_reg[144][4]  ( .D(n8232), .E(n498), .CK(clk), .Q(
        \registers[144][4] ) );
  EDFFX1 \registers_reg[144][3]  ( .D(n8184), .E(n498), .CK(clk), .Q(
        \registers[144][3] ) );
  EDFFX1 \registers_reg[144][2]  ( .D(n8136), .E(n498), .CK(clk), .Q(
        \registers[144][2] ) );
  EDFFX1 \registers_reg[144][1]  ( .D(n8080), .E(n498), .CK(clk), .Q(
        \registers[144][1] ) );
  EDFFX1 \registers_reg[144][0]  ( .D(n8019), .E(n498), .CK(clk), .Q(
        \registers[144][0] ) );
  EDFFX1 \registers_reg[140][7]  ( .D(n8404), .E(n494), .CK(clk), .Q(
        \registers[140][7] ) );
  EDFFX1 \registers_reg[140][6]  ( .D(n8346), .E(n494), .CK(clk), .Q(
        \registers[140][6] ) );
  EDFFX1 \registers_reg[140][5]  ( .D(n8288), .E(n494), .CK(clk), .Q(
        \registers[140][5] ) );
  EDFFX1 \registers_reg[140][4]  ( .D(n8230), .E(n494), .CK(clk), .Q(
        \registers[140][4] ) );
  EDFFX1 \registers_reg[140][3]  ( .D(n8182), .E(n494), .CK(clk), .Q(
        \registers[140][3] ) );
  EDFFX1 \registers_reg[140][2]  ( .D(n8137), .E(n494), .CK(clk), .Q(
        \registers[140][2] ) );
  EDFFX1 \registers_reg[140][1]  ( .D(n8081), .E(n494), .CK(clk), .Q(
        \registers[140][1] ) );
  EDFFX1 \registers_reg[140][0]  ( .D(n8020), .E(n494), .CK(clk), .Q(
        \registers[140][0] ) );
  EDFFX1 \registers_reg[136][7]  ( .D(n8405), .E(n490), .CK(clk), .Q(
        \registers[136][7] ) );
  EDFFX1 \registers_reg[136][6]  ( .D(n8347), .E(n490), .CK(clk), .Q(
        \registers[136][6] ) );
  EDFFX1 \registers_reg[136][5]  ( .D(n8289), .E(n490), .CK(clk), .Q(
        \registers[136][5] ) );
  EDFFX1 \registers_reg[136][4]  ( .D(n8231), .E(n490), .CK(clk), .Q(
        \registers[136][4] ) );
  EDFFX1 \registers_reg[136][3]  ( .D(n8183), .E(n490), .CK(clk), .Q(
        \registers[136][3] ) );
  EDFFX1 \registers_reg[136][2]  ( .D(n8135), .E(n490), .CK(clk), .Q(
        \registers[136][2] ) );
  EDFFX1 \registers_reg[136][1]  ( .D(n8079), .E(n490), .CK(clk), .Q(
        \registers[136][1] ) );
  EDFFX1 \registers_reg[136][0]  ( .D(n8021), .E(n490), .CK(clk), .Q(
        \registers[136][0] ) );
  EDFFX1 \registers_reg[132][7]  ( .D(n8406), .E(n1018), .CK(clk), .Q(
        \registers[132][7] ) );
  EDFFX1 \registers_reg[132][6]  ( .D(n8348), .E(n1018), .CK(clk), .Q(
        \registers[132][6] ) );
  EDFFX1 \registers_reg[132][5]  ( .D(n8290), .E(n1018), .CK(clk), .Q(
        \registers[132][5] ) );
  EDFFX1 \registers_reg[132][4]  ( .D(n8232), .E(n1018), .CK(clk), .Q(
        \registers[132][4] ) );
  EDFFX1 \registers_reg[132][3]  ( .D(n8184), .E(n1018), .CK(clk), .Q(
        \registers[132][3] ) );
  EDFFX1 \registers_reg[132][2]  ( .D(n8136), .E(n1018), .CK(clk), .Q(
        \registers[132][2] ) );
  EDFFX1 \registers_reg[132][1]  ( .D(n8080), .E(n1018), .CK(clk), .Q(
        \registers[132][1] ) );
  EDFFX1 \registers_reg[132][0]  ( .D(n8019), .E(n1018), .CK(clk), .Q(
        \registers[132][0] ) );
  EDFFX1 \registers_reg[128][7]  ( .D(n8421), .E(n387), .CK(clk), .Q(
        \registers[128][7] ) );
  EDFFX1 \registers_reg[128][6]  ( .D(n8363), .E(n387), .CK(clk), .Q(
        \registers[128][6] ) );
  EDFFX1 \registers_reg[128][5]  ( .D(n8305), .E(n387), .CK(clk), .Q(
        \registers[128][5] ) );
  EDFFX1 \registers_reg[128][4]  ( .D(n8247), .E(n387), .CK(clk), .Q(
        \registers[128][4] ) );
  EDFFX1 \registers_reg[128][3]  ( .D(n8195), .E(n387), .CK(clk), .Q(
        \registers[128][3] ) );
  EDFFX1 \registers_reg[128][2]  ( .D(n8150), .E(n387), .CK(clk), .Q(
        \registers[128][2] ) );
  EDFFX1 \registers_reg[128][1]  ( .D(n8094), .E(n387), .CK(clk), .Q(
        \registers[128][1] ) );
  EDFFX1 \registers_reg[128][0]  ( .D(n8035), .E(n387), .CK(clk), .Q(
        \registers[128][0] ) );
  EDFFX1 \registers_reg[124][7]  ( .D(n8419), .E(n486), .CK(clk), .Q(
        \registers[124][7] ) );
  EDFFX1 \registers_reg[124][6]  ( .D(n8361), .E(n486), .CK(clk), .Q(
        \registers[124][6] ) );
  EDFFX1 \registers_reg[124][5]  ( .D(n8303), .E(n486), .CK(clk), .Q(
        \registers[124][5] ) );
  EDFFX1 \registers_reg[124][4]  ( .D(n8245), .E(n486), .CK(clk), .Q(
        \registers[124][4] ) );
  EDFFX1 \registers_reg[124][3]  ( .D(n8196), .E(n486), .CK(clk), .Q(
        \registers[124][3] ) );
  EDFFX1 \registers_reg[124][2]  ( .D(n8151), .E(n486), .CK(clk), .Q(
        \registers[124][2] ) );
  EDFFX1 \registers_reg[124][1]  ( .D(n8095), .E(n486), .CK(clk), .Q(
        \registers[124][1] ) );
  EDFFX1 \registers_reg[124][0]  ( .D(n8035), .E(n486), .CK(clk), .Q(
        \registers[124][0] ) );
  EDFFX1 \registers_reg[120][7]  ( .D(n8420), .E(n482), .CK(clk), .Q(
        \registers[120][7] ) );
  EDFFX1 \registers_reg[120][6]  ( .D(n8362), .E(n482), .CK(clk), .Q(
        \registers[120][6] ) );
  EDFFX1 \registers_reg[120][5]  ( .D(n8304), .E(n482), .CK(clk), .Q(
        \registers[120][5] ) );
  EDFFX1 \registers_reg[120][4]  ( .D(n8246), .E(n482), .CK(clk), .Q(
        \registers[120][4] ) );
  EDFFX1 \registers_reg[120][3]  ( .D(n8194), .E(n482), .CK(clk), .Q(
        \registers[120][3] ) );
  EDFFX1 \registers_reg[120][2]  ( .D(n8730), .E(n482), .CK(clk), .Q(
        \registers[120][2] ) );
  EDFFX1 \registers_reg[120][1]  ( .D(n8702), .E(n482), .CK(clk), .Q(
        \registers[120][1] ) );
  EDFFX1 \registers_reg[120][0]  ( .D(n8036), .E(n482), .CK(clk), .Q(
        \registers[120][0] ) );
  EDFFX1 \registers_reg[116][7]  ( .D(n8421), .E(n478), .CK(clk), .Q(
        \registers[116][7] ) );
  EDFFX1 \registers_reg[116][6]  ( .D(n8363), .E(n478), .CK(clk), .Q(
        \registers[116][6] ) );
  EDFFX1 \registers_reg[116][5]  ( .D(n8305), .E(n478), .CK(clk), .Q(
        \registers[116][5] ) );
  EDFFX1 \registers_reg[116][4]  ( .D(n8247), .E(n478), .CK(clk), .Q(
        \registers[116][4] ) );
  EDFFX1 \registers_reg[116][3]  ( .D(n8195), .E(n478), .CK(clk), .Q(
        \registers[116][3] ) );
  EDFFX1 \registers_reg[116][2]  ( .D(n8147), .E(n478), .CK(clk), .Q(
        \registers[116][2] ) );
  EDFFX1 \registers_reg[116][1]  ( .D(n8091), .E(n478), .CK(clk), .Q(
        \registers[116][1] ) );
  EDFFX1 \registers_reg[116][0]  ( .D(n8031), .E(n478), .CK(clk), .Q(
        \registers[116][0] ) );
  EDFFX1 \registers_reg[112][7]  ( .D(n8419), .E(n474), .CK(clk), .Q(
        \registers[112][7] ) );
  EDFFX1 \registers_reg[112][6]  ( .D(n8361), .E(n474), .CK(clk), .Q(
        \registers[112][6] ) );
  EDFFX1 \registers_reg[112][5]  ( .D(n8303), .E(n474), .CK(clk), .Q(
        \registers[112][5] ) );
  EDFFX1 \registers_reg[112][4]  ( .D(n8245), .E(n474), .CK(clk), .Q(
        \registers[112][4] ) );
  EDFFX1 \registers_reg[112][3]  ( .D(n8196), .E(n474), .CK(clk), .Q(
        \registers[112][3] ) );
  EDFFX1 \registers_reg[112][2]  ( .D(n8148), .E(n474), .CK(clk), .Q(
        \registers[112][2] ) );
  EDFFX1 \registers_reg[112][1]  ( .D(n8092), .E(n474), .CK(clk), .Q(
        \registers[112][1] ) );
  EDFFX1 \registers_reg[112][0]  ( .D(n8032), .E(n474), .CK(clk), .Q(
        \registers[112][0] ) );
  EDFFX1 \registers_reg[108][7]  ( .D(n8420), .E(n470), .CK(clk), .Q(
        \registers[108][7] ) );
  EDFFX1 \registers_reg[108][6]  ( .D(n8362), .E(n470), .CK(clk), .Q(
        \registers[108][6] ) );
  EDFFX1 \registers_reg[108][5]  ( .D(n8304), .E(n470), .CK(clk), .Q(
        \registers[108][5] ) );
  EDFFX1 \registers_reg[108][4]  ( .D(n8246), .E(n470), .CK(clk), .Q(
        \registers[108][4] ) );
  EDFFX1 \registers_reg[108][3]  ( .D(n8194), .E(n470), .CK(clk), .Q(
        \registers[108][3] ) );
  EDFFX1 \registers_reg[108][2]  ( .D(n8149), .E(n470), .CK(clk), .Q(
        \registers[108][2] ) );
  EDFFX1 \registers_reg[108][1]  ( .D(n8093), .E(n470), .CK(clk), .Q(
        \registers[108][1] ) );
  EDFFX1 \registers_reg[108][0]  ( .D(n8033), .E(n470), .CK(clk), .Q(
        \registers[108][0] ) );
  EDFFX1 \registers_reg[104][7]  ( .D(n8421), .E(n466), .CK(clk), .Q(
        \registers[104][7] ) );
  EDFFX1 \registers_reg[104][6]  ( .D(n8363), .E(n466), .CK(clk), .Q(
        \registers[104][6] ) );
  EDFFX1 \registers_reg[104][5]  ( .D(n8305), .E(n466), .CK(clk), .Q(
        \registers[104][5] ) );
  EDFFX1 \registers_reg[104][4]  ( .D(n8247), .E(n466), .CK(clk), .Q(
        \registers[104][4] ) );
  EDFFX1 \registers_reg[104][3]  ( .D(n8192), .E(n466), .CK(clk), .Q(
        \registers[104][3] ) );
  EDFFX1 \registers_reg[104][2]  ( .D(n8147), .E(n466), .CK(clk), .Q(
        \registers[104][2] ) );
  EDFFX1 \registers_reg[104][1]  ( .D(n8091), .E(n466), .CK(clk), .Q(
        \registers[104][1] ) );
  EDFFX1 \registers_reg[104][0]  ( .D(n8031), .E(n466), .CK(clk), .Q(
        \registers[104][0] ) );
  EDFFX1 \registers_reg[100][7]  ( .D(n8417), .E(n951), .CK(clk), .Q(
        \registers[100][7] ) );
  EDFFX1 \registers_reg[100][6]  ( .D(n8359), .E(n951), .CK(clk), .Q(
        \registers[100][6] ) );
  EDFFX1 \registers_reg[100][5]  ( .D(n8301), .E(n951), .CK(clk), .Q(
        \registers[100][5] ) );
  EDFFX1 \registers_reg[100][4]  ( .D(n8243), .E(n951), .CK(clk), .Q(
        \registers[100][4] ) );
  EDFFX1 \registers_reg[100][3]  ( .D(n8193), .E(n951), .CK(clk), .Q(
        \registers[100][3] ) );
  EDFFX1 \registers_reg[100][2]  ( .D(n8148), .E(n951), .CK(clk), .Q(
        \registers[100][2] ) );
  EDFFX1 \registers_reg[100][1]  ( .D(n8092), .E(n951), .CK(clk), .Q(
        \registers[100][1] ) );
  EDFFX1 \registers_reg[100][0]  ( .D(n8032), .E(n951), .CK(clk), .Q(
        \registers[100][0] ) );
  EDFFX1 \registers_reg[96][7]  ( .D(n8418), .E(n344), .CK(clk), .Q(
        \registers[96][7] ) );
  EDFFX1 \registers_reg[96][6]  ( .D(n8360), .E(n344), .CK(clk), .Q(
        \registers[96][6] ) );
  EDFFX1 \registers_reg[96][5]  ( .D(n8302), .E(n344), .CK(clk), .Q(
        \registers[96][5] ) );
  EDFFX1 \registers_reg[96][4]  ( .D(n8244), .E(n344), .CK(clk), .Q(
        \registers[96][4] ) );
  EDFFX1 \registers_reg[96][3]  ( .D(n8191), .E(n344), .CK(clk), .Q(
        \registers[96][3] ) );
  EDFFX1 \registers_reg[96][2]  ( .D(n8149), .E(n344), .CK(clk), .Q(
        \registers[96][2] ) );
  EDFFX1 \registers_reg[96][1]  ( .D(n8093), .E(n344), .CK(clk), .Q(
        \registers[96][1] ) );
  EDFFX1 \registers_reg[96][0]  ( .D(n8033), .E(n344), .CK(clk), .Q(
        \registers[96][0] ) );
  EDFFX1 \registers_reg[92][7]  ( .D(n8416), .E(n462), .CK(clk), .Q(
        \registers[92][7] ) );
  EDFFX1 \registers_reg[92][6]  ( .D(n8358), .E(n462), .CK(clk), .Q(
        \registers[92][6] ) );
  EDFFX1 \registers_reg[92][5]  ( .D(n8300), .E(n462), .CK(clk), .Q(
        \registers[92][5] ) );
  EDFFX1 \registers_reg[92][4]  ( .D(n8242), .E(n462), .CK(clk), .Q(
        \registers[92][4] ) );
  EDFFX1 \registers_reg[92][3]  ( .D(n8192), .E(n462), .CK(clk), .Q(
        \registers[92][3] ) );
  EDFFX1 \registers_reg[92][2]  ( .D(n8147), .E(n462), .CK(clk), .Q(
        \registers[92][2] ) );
  EDFFX1 \registers_reg[92][1]  ( .D(n8091), .E(n462), .CK(clk), .Q(
        \registers[92][1] ) );
  EDFFX1 \registers_reg[92][0]  ( .D(n8031), .E(n462), .CK(clk), .Q(
        \registers[92][0] ) );
  EDFFX1 \registers_reg[88][7]  ( .D(n8417), .E(n458), .CK(clk), .Q(
        \registers[88][7] ) );
  EDFFX1 \registers_reg[88][6]  ( .D(n8359), .E(n458), .CK(clk), .Q(
        \registers[88][6] ) );
  EDFFX1 \registers_reg[88][5]  ( .D(n8301), .E(n458), .CK(clk), .Q(
        \registers[88][5] ) );
  EDFFX1 \registers_reg[88][4]  ( .D(n8243), .E(n458), .CK(clk), .Q(
        \registers[88][4] ) );
  EDFFX1 \registers_reg[88][3]  ( .D(n8193), .E(n458), .CK(clk), .Q(
        \registers[88][3] ) );
  EDFFX1 \registers_reg[88][2]  ( .D(n8148), .E(n458), .CK(clk), .Q(
        \registers[88][2] ) );
  EDFFX1 \registers_reg[88][1]  ( .D(n8092), .E(n458), .CK(clk), .Q(
        \registers[88][1] ) );
  EDFFX1 \registers_reg[88][0]  ( .D(n8032), .E(n458), .CK(clk), .Q(
        \registers[88][0] ) );
  EDFFX1 \registers_reg[84][7]  ( .D(n8418), .E(n454), .CK(clk), .Q(
        \registers[84][7] ) );
  EDFFX1 \registers_reg[84][6]  ( .D(n8360), .E(n454), .CK(clk), .Q(
        \registers[84][6] ) );
  EDFFX1 \registers_reg[84][5]  ( .D(n8302), .E(n454), .CK(clk), .Q(
        \registers[84][5] ) );
  EDFFX1 \registers_reg[84][4]  ( .D(n8244), .E(n454), .CK(clk), .Q(
        \registers[84][4] ) );
  EDFFX1 \registers_reg[84][3]  ( .D(n8191), .E(n454), .CK(clk), .Q(
        \registers[84][3] ) );
  EDFFX1 \registers_reg[84][2]  ( .D(n8149), .E(n454), .CK(clk), .Q(
        \registers[84][2] ) );
  EDFFX1 \registers_reg[84][1]  ( .D(n8093), .E(n454), .CK(clk), .Q(
        \registers[84][1] ) );
  EDFFX1 \registers_reg[84][0]  ( .D(n8033), .E(n454), .CK(clk), .Q(
        \registers[84][0] ) );
  EDFFX1 \registers_reg[80][7]  ( .D(n8416), .E(n450), .CK(clk), .Q(
        \registers[80][7] ) );
  EDFFX1 \registers_reg[80][6]  ( .D(n8358), .E(n450), .CK(clk), .Q(
        \registers[80][6] ) );
  EDFFX1 \registers_reg[80][5]  ( .D(n8300), .E(n450), .CK(clk), .Q(
        \registers[80][5] ) );
  EDFFX1 \registers_reg[80][4]  ( .D(n8242), .E(n450), .CK(clk), .Q(
        \registers[80][4] ) );
  EDFFX1 \registers_reg[80][3]  ( .D(n8192), .E(n450), .CK(clk), .Q(
        \registers[80][3] ) );
  EDFFX1 \registers_reg[80][2]  ( .D(n8147), .E(n450), .CK(clk), .Q(
        \registers[80][2] ) );
  EDFFX1 \registers_reg[80][1]  ( .D(n8091), .E(n450), .CK(clk), .Q(
        \registers[80][1] ) );
  EDFFX1 \registers_reg[80][0]  ( .D(n8031), .E(n450), .CK(clk), .Q(
        \registers[80][0] ) );
  EDFFX1 \registers_reg[76][7]  ( .D(n8417), .E(n446), .CK(clk), .Q(
        \registers[76][7] ) );
  EDFFX1 \registers_reg[76][6]  ( .D(n8359), .E(n446), .CK(clk), .Q(
        \registers[76][6] ) );
  EDFFX1 \registers_reg[76][5]  ( .D(n8301), .E(n446), .CK(clk), .Q(
        \registers[76][5] ) );
  EDFFX1 \registers_reg[76][4]  ( .D(n8243), .E(n446), .CK(clk), .Q(
        \registers[76][4] ) );
  EDFFX1 \registers_reg[76][3]  ( .D(n8193), .E(n446), .CK(clk), .Q(
        \registers[76][3] ) );
  EDFFX1 \registers_reg[76][2]  ( .D(n8148), .E(n446), .CK(clk), .Q(
        \registers[76][2] ) );
  EDFFX1 \registers_reg[76][1]  ( .D(n8092), .E(n446), .CK(clk), .Q(
        \registers[76][1] ) );
  EDFFX1 \registers_reg[76][0]  ( .D(n8032), .E(n446), .CK(clk), .Q(
        \registers[76][0] ) );
  EDFFX1 \registers_reg[72][7]  ( .D(n8418), .E(n442), .CK(clk), .Q(
        \registers[72][7] ) );
  EDFFX1 \registers_reg[72][6]  ( .D(n8360), .E(n442), .CK(clk), .Q(
        \registers[72][6] ) );
  EDFFX1 \registers_reg[72][5]  ( .D(n8302), .E(n442), .CK(clk), .Q(
        \registers[72][5] ) );
  EDFFX1 \registers_reg[72][4]  ( .D(n8244), .E(n442), .CK(clk), .Q(
        \registers[72][4] ) );
  EDFFX1 \registers_reg[72][3]  ( .D(n8191), .E(n442), .CK(clk), .Q(
        \registers[72][3] ) );
  EDFFX1 \registers_reg[72][2]  ( .D(n8149), .E(n442), .CK(clk), .Q(
        \registers[72][2] ) );
  EDFFX1 \registers_reg[72][1]  ( .D(n8093), .E(n442), .CK(clk), .Q(
        \registers[72][1] ) );
  EDFFX1 \registers_reg[72][0]  ( .D(n8033), .E(n442), .CK(clk), .Q(
        \registers[72][0] ) );
  EDFFX1 \registers_reg[68][7]  ( .D(n8416), .E(n944), .CK(clk), .Q(
        \registers[68][7] ) );
  EDFFX1 \registers_reg[68][6]  ( .D(n8358), .E(n944), .CK(clk), .Q(
        \registers[68][6] ) );
  EDFFX1 \registers_reg[68][5]  ( .D(n8300), .E(n944), .CK(clk), .Q(
        \registers[68][5] ) );
  EDFFX1 \registers_reg[68][4]  ( .D(n8242), .E(n944), .CK(clk), .Q(
        \registers[68][4] ) );
  EDFFX1 \registers_reg[68][3]  ( .D(n8192), .E(n944), .CK(clk), .Q(
        \registers[68][3] ) );
  EDFFX1 \registers_reg[68][2]  ( .D(n8147), .E(n944), .CK(clk), .Q(
        \registers[68][2] ) );
  EDFFX1 \registers_reg[68][1]  ( .D(n8091), .E(n944), .CK(clk), .Q(
        \registers[68][1] ) );
  EDFFX1 \registers_reg[68][0]  ( .D(n8031), .E(n944), .CK(clk), .Q(
        \registers[68][0] ) );
  EDFFX1 \registers_reg[64][7]  ( .D(n8418), .E(n343), .CK(clk), .Q(
        \registers[64][7] ) );
  EDFFX1 \registers_reg[64][6]  ( .D(n8360), .E(n343), .CK(clk), .Q(
        \registers[64][6] ) );
  EDFFX1 \registers_reg[64][5]  ( .D(n8302), .E(n343), .CK(clk), .Q(
        \registers[64][5] ) );
  EDFFX1 \registers_reg[64][4]  ( .D(n8244), .E(n343), .CK(clk), .Q(
        \registers[64][4] ) );
  EDFFX1 \registers_reg[64][3]  ( .D(n8191), .E(n343), .CK(clk), .Q(
        \registers[64][3] ) );
  EDFFX1 \registers_reg[64][2]  ( .D(n8146), .E(n343), .CK(clk), .Q(
        \registers[64][2] ) );
  EDFFX1 \registers_reg[64][1]  ( .D(n8090), .E(n343), .CK(clk), .Q(
        \registers[64][1] ) );
  EDFFX1 \registers_reg[64][0]  ( .D(n8030), .E(n343), .CK(clk), .Q(
        \registers[64][0] ) );
  EDFFX1 \registers_reg[60][7]  ( .D(n8416), .E(n438), .CK(clk), .Q(
        \registers[60][7] ) );
  EDFFX1 \registers_reg[60][6]  ( .D(n8358), .E(n438), .CK(clk), .Q(
        \registers[60][6] ) );
  EDFFX1 \registers_reg[60][5]  ( .D(n8300), .E(n438), .CK(clk), .Q(
        \registers[60][5] ) );
  EDFFX1 \registers_reg[60][4]  ( .D(n8242), .E(n438), .CK(clk), .Q(
        \registers[60][4] ) );
  EDFFX1 \registers_reg[60][3]  ( .D(n8192), .E(n438), .CK(clk), .Q(
        \registers[60][3] ) );
  EDFFX1 \registers_reg[60][2]  ( .D(n8144), .E(n438), .CK(clk), .Q(
        \registers[60][2] ) );
  EDFFX1 \registers_reg[60][1]  ( .D(n8088), .E(n438), .CK(clk), .Q(
        \registers[60][1] ) );
  EDFFX1 \registers_reg[60][0]  ( .D(n8028), .E(n438), .CK(clk), .Q(
        \registers[60][0] ) );
  EDFFX1 \registers_reg[56][7]  ( .D(n8417), .E(n434), .CK(clk), .Q(
        \registers[56][7] ) );
  EDFFX1 \registers_reg[56][6]  ( .D(n8359), .E(n434), .CK(clk), .Q(
        \registers[56][6] ) );
  EDFFX1 \registers_reg[56][5]  ( .D(n8301), .E(n434), .CK(clk), .Q(
        \registers[56][5] ) );
  EDFFX1 \registers_reg[56][4]  ( .D(n8243), .E(n434), .CK(clk), .Q(
        \registers[56][4] ) );
  EDFFX1 \registers_reg[56][3]  ( .D(n8193), .E(n434), .CK(clk), .Q(
        \registers[56][3] ) );
  EDFFX1 \registers_reg[56][2]  ( .D(n8145), .E(n434), .CK(clk), .Q(
        \registers[56][2] ) );
  EDFFX1 \registers_reg[56][1]  ( .D(n8089), .E(n434), .CK(clk), .Q(
        \registers[56][1] ) );
  EDFFX1 \registers_reg[56][0]  ( .D(n8029), .E(n434), .CK(clk), .Q(
        \registers[56][0] ) );
  EDFFX1 \registers_reg[52][7]  ( .D(n8413), .E(n430), .CK(clk), .Q(
        \registers[52][7] ) );
  EDFFX1 \registers_reg[52][6]  ( .D(n8355), .E(n430), .CK(clk), .Q(
        \registers[52][6] ) );
  EDFFX1 \registers_reg[52][5]  ( .D(n8297), .E(n430), .CK(clk), .Q(
        \registers[52][5] ) );
  EDFFX1 \registers_reg[52][4]  ( .D(n8239), .E(n430), .CK(clk), .Q(
        \registers[52][4] ) );
  EDFFX1 \registers_reg[52][3]  ( .D(n8191), .E(n430), .CK(clk), .Q(
        \registers[52][3] ) );
  EDFFX1 \registers_reg[52][2]  ( .D(n8146), .E(n430), .CK(clk), .Q(
        \registers[52][2] ) );
  EDFFX1 \registers_reg[52][1]  ( .D(n8090), .E(n430), .CK(clk), .Q(
        \registers[52][1] ) );
  EDFFX1 \registers_reg[52][0]  ( .D(n8030), .E(n430), .CK(clk), .Q(
        \registers[52][0] ) );
  EDFFX1 \registers_reg[48][7]  ( .D(n8414), .E(n426), .CK(clk), .Q(
        \registers[48][7] ) );
  EDFFX1 \registers_reg[48][6]  ( .D(n8356), .E(n426), .CK(clk), .Q(
        \registers[48][6] ) );
  EDFFX1 \registers_reg[48][5]  ( .D(n8298), .E(n426), .CK(clk), .Q(
        \registers[48][5] ) );
  EDFFX1 \registers_reg[48][4]  ( .D(n8240), .E(n426), .CK(clk), .Q(
        \registers[48][4] ) );
  EDFFX1 \registers_reg[48][3]  ( .D(n8192), .E(n426), .CK(clk), .Q(
        \registers[48][3] ) );
  EDFFX1 \registers_reg[48][2]  ( .D(n8144), .E(n426), .CK(clk), .Q(
        \registers[48][2] ) );
  EDFFX1 \registers_reg[48][1]  ( .D(n8088), .E(n426), .CK(clk), .Q(
        \registers[48][1] ) );
  EDFFX1 \registers_reg[48][0]  ( .D(n8028), .E(n426), .CK(clk), .Q(
        \registers[48][0] ) );
  EDFFX1 \registers_reg[44][7]  ( .D(n8415), .E(n422), .CK(clk), .Q(
        \registers[44][7] ) );
  EDFFX1 \registers_reg[44][6]  ( .D(n8357), .E(n422), .CK(clk), .Q(
        \registers[44][6] ) );
  EDFFX1 \registers_reg[44][5]  ( .D(n8299), .E(n422), .CK(clk), .Q(
        \registers[44][5] ) );
  EDFFX1 \registers_reg[44][4]  ( .D(n8241), .E(n422), .CK(clk), .Q(
        \registers[44][4] ) );
  EDFFX1 \registers_reg[44][3]  ( .D(n8193), .E(n422), .CK(clk), .Q(
        \registers[44][3] ) );
  EDFFX1 \registers_reg[44][2]  ( .D(n8145), .E(n422), .CK(clk), .Q(
        \registers[44][2] ) );
  EDFFX1 \registers_reg[44][1]  ( .D(n8089), .E(n422), .CK(clk), .Q(
        \registers[44][1] ) );
  EDFFX1 \registers_reg[44][0]  ( .D(n8029), .E(n422), .CK(clk), .Q(
        \registers[44][0] ) );
  EDFFX1 \registers_reg[40][7]  ( .D(n8413), .E(n418), .CK(clk), .Q(
        \registers[40][7] ) );
  EDFFX1 \registers_reg[40][6]  ( .D(n8355), .E(n418), .CK(clk), .Q(
        \registers[40][6] ) );
  EDFFX1 \registers_reg[40][5]  ( .D(n8297), .E(n418), .CK(clk), .Q(
        \registers[40][5] ) );
  EDFFX1 \registers_reg[40][4]  ( .D(n8239), .E(n418), .CK(clk), .Q(
        \registers[40][4] ) );
  EDFFX1 \registers_reg[40][3]  ( .D(n8188), .E(n418), .CK(clk), .Q(
        \registers[40][3] ) );
  EDFFX1 \registers_reg[40][2]  ( .D(n8146), .E(n418), .CK(clk), .Q(
        \registers[40][2] ) );
  EDFFX1 \registers_reg[40][1]  ( .D(n8090), .E(n418), .CK(clk), .Q(
        \registers[40][1] ) );
  EDFFX1 \registers_reg[40][0]  ( .D(n8030), .E(n418), .CK(clk), .Q(
        \registers[40][0] ) );
  EDFFX1 \registers_reg[36][7]  ( .D(n8414), .E(n937), .CK(clk), .Q(
        \registers[36][7] ) );
  EDFFX1 \registers_reg[36][6]  ( .D(n8356), .E(n937), .CK(clk), .Q(
        \registers[36][6] ) );
  EDFFX1 \registers_reg[36][5]  ( .D(n8298), .E(n937), .CK(clk), .Q(
        \registers[36][5] ) );
  EDFFX1 \registers_reg[36][4]  ( .D(n8240), .E(n937), .CK(clk), .Q(
        \registers[36][4] ) );
  EDFFX1 \registers_reg[36][3]  ( .D(n8189), .E(n937), .CK(clk), .Q(
        \registers[36][3] ) );
  EDFFX1 \registers_reg[36][2]  ( .D(n8144), .E(n937), .CK(clk), .Q(
        \registers[36][2] ) );
  EDFFX1 \registers_reg[36][1]  ( .D(n8088), .E(n937), .CK(clk), .Q(
        \registers[36][1] ) );
  EDFFX1 \registers_reg[36][0]  ( .D(n8028), .E(n937), .CK(clk), .Q(
        \registers[36][0] ) );
  EDFFX1 \registers_reg[32][7]  ( .D(n8415), .E(n342), .CK(clk), .Q(
        \registers[32][7] ) );
  EDFFX1 \registers_reg[32][6]  ( .D(n8357), .E(n342), .CK(clk), .Q(
        \registers[32][6] ) );
  EDFFX1 \registers_reg[32][5]  ( .D(n8299), .E(n342), .CK(clk), .Q(
        \registers[32][5] ) );
  EDFFX1 \registers_reg[32][4]  ( .D(n8241), .E(n342), .CK(clk), .Q(
        \registers[32][4] ) );
  EDFFX1 \registers_reg[32][3]  ( .D(n8190), .E(n342), .CK(clk), .Q(
        \registers[32][3] ) );
  EDFFX1 \registers_reg[32][2]  ( .D(n8145), .E(n342), .CK(clk), .Q(
        \registers[32][2] ) );
  EDFFX1 \registers_reg[32][1]  ( .D(n8089), .E(n342), .CK(clk), .Q(
        \registers[32][1] ) );
  EDFFX1 \registers_reg[32][0]  ( .D(n8029), .E(n342), .CK(clk), .Q(
        \registers[32][0] ) );
  EDFFX1 \registers_reg[28][7]  ( .D(n8413), .E(n414), .CK(clk), .Q(
        \registers[28][7] ) );
  EDFFX1 \registers_reg[28][6]  ( .D(n8355), .E(n414), .CK(clk), .Q(
        \registers[28][6] ) );
  EDFFX1 \registers_reg[28][5]  ( .D(n8297), .E(n414), .CK(clk), .Q(
        \registers[28][5] ) );
  EDFFX1 \registers_reg[28][4]  ( .D(n8239), .E(n414), .CK(clk), .Q(
        \registers[28][4] ) );
  EDFFX1 \registers_reg[28][3]  ( .D(n8188), .E(n414), .CK(clk), .Q(
        \registers[28][3] ) );
  EDFFX1 \registers_reg[28][2]  ( .D(n8146), .E(n414), .CK(clk), .Q(
        \registers[28][2] ) );
  EDFFX1 \registers_reg[28][1]  ( .D(n8090), .E(n414), .CK(clk), .Q(
        \registers[28][1] ) );
  EDFFX1 \registers_reg[28][0]  ( .D(n8030), .E(n414), .CK(clk), .Q(
        \registers[28][0] ) );
  EDFFX1 \registers_reg[24][7]  ( .D(n8414), .E(n410), .CK(clk), .Q(
        \registers[24][7] ) );
  EDFFX1 \registers_reg[24][6]  ( .D(n8356), .E(n410), .CK(clk), .Q(
        \registers[24][6] ) );
  EDFFX1 \registers_reg[24][5]  ( .D(n8298), .E(n410), .CK(clk), .Q(
        \registers[24][5] ) );
  EDFFX1 \registers_reg[24][4]  ( .D(n8240), .E(n410), .CK(clk), .Q(
        \registers[24][4] ) );
  EDFFX1 \registers_reg[24][3]  ( .D(n8189), .E(n410), .CK(clk), .Q(
        \registers[24][3] ) );
  EDFFX1 \registers_reg[24][2]  ( .D(n8144), .E(n410), .CK(clk), .Q(
        \registers[24][2] ) );
  EDFFX1 \registers_reg[24][1]  ( .D(n8088), .E(n410), .CK(clk), .Q(
        \registers[24][1] ) );
  EDFFX1 \registers_reg[24][0]  ( .D(n8028), .E(n410), .CK(clk), .Q(
        \registers[24][0] ) );
  EDFFX1 \registers_reg[20][7]  ( .D(n8415), .E(n406), .CK(clk), .Q(
        \registers[20][7] ) );
  EDFFX1 \registers_reg[20][6]  ( .D(n8357), .E(n406), .CK(clk), .Q(
        \registers[20][6] ) );
  EDFFX1 \registers_reg[20][5]  ( .D(n8299), .E(n406), .CK(clk), .Q(
        \registers[20][5] ) );
  EDFFX1 \registers_reg[20][4]  ( .D(n8241), .E(n406), .CK(clk), .Q(
        \registers[20][4] ) );
  EDFFX1 \registers_reg[20][3]  ( .D(n8190), .E(n406), .CK(clk), .Q(
        \registers[20][3] ) );
  EDFFX1 \registers_reg[20][2]  ( .D(n8145), .E(n406), .CK(clk), .Q(
        \registers[20][2] ) );
  EDFFX1 \registers_reg[20][1]  ( .D(n8089), .E(n406), .CK(clk), .Q(
        \registers[20][1] ) );
  EDFFX1 \registers_reg[20][0]  ( .D(n8029), .E(n406), .CK(clk), .Q(
        \registers[20][0] ) );
  EDFFX1 \registers_reg[16][7]  ( .D(n8413), .E(n402), .CK(clk), .Q(
        \registers[16][7] ) );
  EDFFX1 \registers_reg[16][6]  ( .D(n8355), .E(n402), .CK(clk), .Q(
        \registers[16][6] ) );
  EDFFX1 \registers_reg[16][5]  ( .D(n8297), .E(n402), .CK(clk), .Q(
        \registers[16][5] ) );
  EDFFX1 \registers_reg[16][4]  ( .D(n8239), .E(n402), .CK(clk), .Q(
        \registers[16][4] ) );
  EDFFX1 \registers_reg[16][3]  ( .D(n8188), .E(n402), .CK(clk), .Q(
        \registers[16][3] ) );
  EDFFX1 \registers_reg[16][2]  ( .D(n8146), .E(n402), .CK(clk), .Q(
        \registers[16][2] ) );
  EDFFX1 \registers_reg[16][1]  ( .D(n8090), .E(n402), .CK(clk), .Q(
        \registers[16][1] ) );
  EDFFX1 \registers_reg[16][0]  ( .D(n8030), .E(n402), .CK(clk), .Q(
        \registers[16][0] ) );
  EDFFX1 \registers_reg[12][7]  ( .D(n8414), .E(n398), .CK(clk), .Q(
        \registers[12][7] ) );
  EDFFX1 \registers_reg[12][6]  ( .D(n8356), .E(n398), .CK(clk), .Q(
        \registers[12][6] ) );
  EDFFX1 \registers_reg[12][5]  ( .D(n8298), .E(n398), .CK(clk), .Q(
        \registers[12][5] ) );
  EDFFX1 \registers_reg[12][4]  ( .D(n8240), .E(n398), .CK(clk), .Q(
        \registers[12][4] ) );
  EDFFX1 \registers_reg[12][3]  ( .D(n8189), .E(n398), .CK(clk), .Q(
        \registers[12][3] ) );
  EDFFX1 \registers_reg[12][2]  ( .D(n8141), .E(n398), .CK(clk), .Q(
        \registers[12][2] ) );
  EDFFX1 \registers_reg[12][1]  ( .D(n8085), .E(n398), .CK(clk), .Q(
        \registers[12][1] ) );
  EDFFX1 \registers_reg[12][0]  ( .D(n8025), .E(n398), .CK(clk), .Q(
        \registers[12][0] ) );
  EDFFX1 \registers_reg[8][7]  ( .D(n8415), .E(n394), .CK(clk), .Q(
        \registers[8][7] ) );
  EDFFX1 \registers_reg[8][6]  ( .D(n8357), .E(n394), .CK(clk), .Q(
        \registers[8][6] ) );
  EDFFX1 \registers_reg[8][5]  ( .D(n8299), .E(n394), .CK(clk), .Q(
        \registers[8][5] ), .QN(n1114) );
  EDFFX1 \registers_reg[8][4]  ( .D(n8241), .E(n394), .CK(clk), .Q(
        \registers[8][4] ), .QN(n1115) );
  EDFFX1 \registers_reg[8][3]  ( .D(n8190), .E(n394), .CK(clk), .Q(
        \registers[8][3] ), .QN(n1116) );
  EDFFX1 \registers_reg[8][2]  ( .D(n8142), .E(n394), .CK(clk), .Q(
        \registers[8][2] ), .QN(n1117) );
  EDFFX1 \registers_reg[8][1]  ( .D(n8086), .E(n394), .CK(clk), .Q(
        \registers[8][1] ), .QN(n1118) );
  EDFFX1 \registers_reg[8][0]  ( .D(n8026), .E(n394), .CK(clk), .Q(
        \registers[8][0] ), .QN(n1119) );
  EDFFX1 \registers_reg[4][7]  ( .D(n8413), .E(n1014), .CK(clk), .Q(
        \registers[4][7] ) );
  EDFFX1 \registers_reg[4][6]  ( .D(n8355), .E(n1014), .CK(clk), .Q(
        \registers[4][6] ) );
  EDFFX1 \registers_reg[4][5]  ( .D(n8297), .E(n1014), .CK(clk), .Q(
        \registers[4][5] ) );
  EDFFX1 \registers_reg[4][4]  ( .D(n8239), .E(n1014), .CK(clk), .Q(
        \registers[4][4] ) );
  EDFFX1 \registers_reg[4][3]  ( .D(n8188), .E(n1014), .CK(clk), .Q(
        \registers[4][3] ) );
  EDFFX1 \registers_reg[4][2]  ( .D(n8143), .E(n1014), .CK(clk), .Q(
        \registers[4][2] ) );
  EDFFX1 \registers_reg[1022][7]  ( .D(n8400), .E(n932), .CK(clk), .Q(
        \registers[1022][7] ) );
  EDFFX1 \registers_reg[1022][6]  ( .D(n8342), .E(n932), .CK(clk), .Q(
        \registers[1022][6] ) );
  EDFFX1 \registers_reg[1022][5]  ( .D(n8284), .E(n932), .CK(clk), .Q(
        \registers[1022][5] ) );
  EDFFX1 \registers_reg[1022][4]  ( .D(n8226), .E(n932), .CK(clk), .Q(
        \registers[1022][4] ) );
  EDFFX1 \registers_reg[1022][3]  ( .D(n8169), .E(n932), .CK(clk), .Q(
        \registers[1022][3] ) );
  EDFFX1 \registers_reg[1022][2]  ( .D(n8107), .E(n932), .CK(clk), .Q(
        \registers[1022][2] ) );
  EDFFX1 \registers_reg[1022][1]  ( .D(n8051), .E(n932), .CK(clk), .Q(
        \registers[1022][1] ) );
  EDFFX1 \registers_reg[1022][0]  ( .D(n8666), .E(n932), .CK(clk), .Q(
        \registers[1022][0] ) );
  EDFFX1 \registers_reg[1018][7]  ( .D(n8396), .E(n928), .CK(clk), .Q(
        \registers[1018][7] ) );
  EDFFX1 \registers_reg[1018][6]  ( .D(n8338), .E(n928), .CK(clk), .Q(
        \registers[1018][6] ) );
  EDFFX1 \registers_reg[1018][5]  ( .D(n8280), .E(n928), .CK(clk), .Q(
        \registers[1018][5] ) );
  EDFFX1 \registers_reg[1018][4]  ( .D(n8222), .E(n928), .CK(clk), .Q(
        \registers[1018][4] ) );
  EDFFX1 \registers_reg[1018][3]  ( .D(n8177), .E(n928), .CK(clk), .Q(
        \registers[1018][3] ) );
  EDFFX1 \registers_reg[1018][2]  ( .D(n8126), .E(n928), .CK(clk), .Q(
        \registers[1018][2] ) );
  EDFFX1 \registers_reg[1018][1]  ( .D(n8070), .E(n928), .CK(clk), .Q(
        \registers[1018][1] ) );
  EDFFX1 \registers_reg[1018][0]  ( .D(n8012), .E(n928), .CK(clk), .Q(
        \registers[1018][0] ) );
  EDFFX1 \registers_reg[1014][7]  ( .D(n8397), .E(n924), .CK(clk), .Q(
        \registers[1014][7] ) );
  EDFFX1 \registers_reg[1014][6]  ( .D(n8339), .E(n924), .CK(clk), .Q(
        \registers[1014][6] ) );
  EDFFX1 \registers_reg[1014][5]  ( .D(n8281), .E(n924), .CK(clk), .Q(
        \registers[1014][5] ) );
  EDFFX1 \registers_reg[1014][4]  ( .D(n8223), .E(n924), .CK(clk), .Q(
        \registers[1014][4] ) );
  EDFFX1 \registers_reg[1014][3]  ( .D(n8178), .E(n924), .CK(clk), .Q(
        \registers[1014][3] ) );
  EDFFX1 \registers_reg[1014][2]  ( .D(n8127), .E(n924), .CK(clk), .Q(
        \registers[1014][2] ) );
  EDFFX1 \registers_reg[1014][1]  ( .D(n8071), .E(n924), .CK(clk), .Q(
        \registers[1014][1] ) );
  EDFFX1 \registers_reg[1014][0]  ( .D(n8010), .E(n924), .CK(clk), .Q(
        \registers[1014][0] ) );
  EDFFX1 \registers_reg[1010][7]  ( .D(n8395), .E(n237), .CK(clk), .Q(
        \registers[1010][7] ) );
  EDFFX1 \registers_reg[1010][6]  ( .D(n8337), .E(n237), .CK(clk), .Q(
        \registers[1010][6] ) );
  EDFFX1 \registers_reg[1010][5]  ( .D(n8279), .E(n237), .CK(clk), .Q(
        \registers[1010][5] ) );
  EDFFX1 \registers_reg[1010][4]  ( .D(n8221), .E(n237), .CK(clk), .Q(
        \registers[1010][4] ) );
  EDFFX1 \registers_reg[1010][3]  ( .D(n8176), .E(n237), .CK(clk), .Q(
        \registers[1010][3] ) );
  EDFFX1 \registers_reg[1010][2]  ( .D(n8128), .E(n237), .CK(clk), .Q(
        \registers[1010][2] ) );
  EDFFX1 \registers_reg[1010][1]  ( .D(n8072), .E(n237), .CK(clk), .Q(
        \registers[1010][1] ) );
  EDFFX1 \registers_reg[1010][0]  ( .D(n8011), .E(n237), .CK(clk), .Q(
        \registers[1010][0] ) );
  EDFFX1 \registers_reg[1006][7]  ( .D(n8396), .E(n233), .CK(clk), .Q(
        \registers[1006][7] ) );
  EDFFX1 \registers_reg[1006][6]  ( .D(n8338), .E(n233), .CK(clk), .Q(
        \registers[1006][6] ) );
  EDFFX1 \registers_reg[1006][5]  ( .D(n8280), .E(n233), .CK(clk), .Q(
        \registers[1006][5] ) );
  EDFFX1 \registers_reg[1006][4]  ( .D(n8222), .E(n233), .CK(clk), .Q(
        \registers[1006][4] ) );
  EDFFX1 \registers_reg[1006][3]  ( .D(n8177), .E(n233), .CK(clk), .Q(
        \registers[1006][3] ) );
  EDFFX1 \registers_reg[1006][2]  ( .D(n8126), .E(n233), .CK(clk), .Q(
        \registers[1006][2] ) );
  EDFFX1 \registers_reg[1006][1]  ( .D(n8070), .E(n233), .CK(clk), .Q(
        \registers[1006][1] ) );
  EDFFX1 \registers_reg[1006][0]  ( .D(n8012), .E(n233), .CK(clk), .Q(
        \registers[1006][0] ) );
  EDFFX1 \registers_reg[1002][7]  ( .D(n8397), .E(n229), .CK(clk), .Q(
        \registers[1002][7] ) );
  EDFFX1 \registers_reg[1002][6]  ( .D(n8339), .E(n229), .CK(clk), .Q(
        \registers[1002][6] ) );
  EDFFX1 \registers_reg[1002][5]  ( .D(n8281), .E(n229), .CK(clk), .Q(
        \registers[1002][5] ) );
  EDFFX1 \registers_reg[1002][4]  ( .D(n8223), .E(n229), .CK(clk), .Q(
        \registers[1002][4] ) );
  EDFFX1 \registers_reg[1002][3]  ( .D(n8175), .E(n229), .CK(clk), .Q(
        \registers[1002][3] ) );
  EDFFX1 \registers_reg[1002][2]  ( .D(n8127), .E(n229), .CK(clk), .Q(
        \registers[1002][2] ) );
  EDFFX1 \registers_reg[1002][1]  ( .D(n8071), .E(n229), .CK(clk), .Q(
        \registers[1002][1] ) );
  EDFFX1 \registers_reg[1002][0]  ( .D(n8010), .E(n229), .CK(clk), .Q(
        \registers[1002][0] ) );
  EDFFX1 \registers_reg[998][7]  ( .D(n8395), .E(n385), .CK(clk), .Q(
        \registers[998][7] ) );
  EDFFX1 \registers_reg[998][6]  ( .D(n8337), .E(n385), .CK(clk), .Q(
        \registers[998][6] ) );
  EDFFX1 \registers_reg[998][5]  ( .D(n8279), .E(n385), .CK(clk), .Q(
        \registers[998][5] ) );
  EDFFX1 \registers_reg[998][4]  ( .D(n8221), .E(n385), .CK(clk), .Q(
        \registers[998][4] ) );
  EDFFX1 \registers_reg[998][3]  ( .D(n8173), .E(n385), .CK(clk), .Q(
        \registers[998][3] ) );
  EDFFX1 \registers_reg[998][2]  ( .D(n8128), .E(n385), .CK(clk), .Q(
        \registers[998][2] ) );
  EDFFX1 \registers_reg[998][1]  ( .D(n8072), .E(n385), .CK(clk), .Q(
        \registers[998][1] ) );
  EDFFX1 \registers_reg[998][0]  ( .D(n8011), .E(n385), .CK(clk), .Q(
        \registers[998][0] ) );
  EDFFX1 \registers_reg[994][7]  ( .D(n8396), .E(n381), .CK(clk), .Q(
        \registers[994][7] ) );
  EDFFX1 \registers_reg[994][6]  ( .D(n8338), .E(n381), .CK(clk), .Q(
        \registers[994][6] ) );
  EDFFX1 \registers_reg[994][5]  ( .D(n8280), .E(n381), .CK(clk), .Q(
        \registers[994][5] ) );
  EDFFX1 \registers_reg[994][4]  ( .D(n8222), .E(n381), .CK(clk), .Q(
        \registers[994][4] ) );
  EDFFX1 \registers_reg[994][3]  ( .D(n8174), .E(n381), .CK(clk), .Q(
        \registers[994][3] ) );
  EDFFX1 \registers_reg[994][2]  ( .D(n8126), .E(n381), .CK(clk), .Q(
        \registers[994][2] ) );
  EDFFX1 \registers_reg[994][1]  ( .D(n8070), .E(n381), .CK(clk), .Q(
        \registers[994][1] ) );
  EDFFX1 \registers_reg[994][0]  ( .D(n8012), .E(n381), .CK(clk), .Q(
        \registers[994][0] ) );
  EDFFX1 \registers_reg[990][7]  ( .D(n8397), .E(n920), .CK(clk), .Q(
        \registers[990][7] ) );
  EDFFX1 \registers_reg[990][6]  ( .D(n8339), .E(n920), .CK(clk), .Q(
        \registers[990][6] ) );
  EDFFX1 \registers_reg[990][5]  ( .D(n8281), .E(n920), .CK(clk), .Q(
        \registers[990][5] ) );
  EDFFX1 \registers_reg[990][4]  ( .D(n8223), .E(n920), .CK(clk), .Q(
        \registers[990][4] ) );
  EDFFX1 \registers_reg[990][3]  ( .D(n8175), .E(n920), .CK(clk), .Q(
        \registers[990][3] ) );
  EDFFX1 \registers_reg[990][2]  ( .D(n8127), .E(n920), .CK(clk), .Q(
        \registers[990][2] ) );
  EDFFX1 \registers_reg[990][1]  ( .D(n8071), .E(n920), .CK(clk), .Q(
        \registers[990][1] ) );
  EDFFX1 \registers_reg[990][0]  ( .D(n8010), .E(n920), .CK(clk), .Q(
        \registers[990][0] ) );
  EDFFX1 \registers_reg[986][7]  ( .D(n8395), .E(n916), .CK(clk), .Q(
        \registers[986][7] ) );
  EDFFX1 \registers_reg[986][6]  ( .D(n8337), .E(n916), .CK(clk), .Q(
        \registers[986][6] ) );
  EDFFX1 \registers_reg[986][5]  ( .D(n8279), .E(n916), .CK(clk), .Q(
        \registers[986][5] ) );
  EDFFX1 \registers_reg[986][4]  ( .D(n8221), .E(n916), .CK(clk), .Q(
        \registers[986][4] ) );
  EDFFX1 \registers_reg[986][3]  ( .D(n8173), .E(n916), .CK(clk), .Q(
        \registers[986][3] ) );
  EDFFX1 \registers_reg[986][2]  ( .D(n8128), .E(n916), .CK(clk), .Q(
        \registers[986][2] ) );
  EDFFX1 \registers_reg[986][1]  ( .D(n8072), .E(n916), .CK(clk), .Q(
        \registers[986][1] ) );
  EDFFX1 \registers_reg[986][0]  ( .D(n8011), .E(n916), .CK(clk), .Q(
        \registers[986][0] ) );
  EDFFX1 \registers_reg[982][7]  ( .D(n8396), .E(n912), .CK(clk), .Q(
        \registers[982][7] ) );
  EDFFX1 \registers_reg[982][6]  ( .D(n8338), .E(n912), .CK(clk), .Q(
        \registers[982][6] ) );
  EDFFX1 \registers_reg[982][5]  ( .D(n8280), .E(n912), .CK(clk), .Q(
        \registers[982][5] ) );
  EDFFX1 \registers_reg[982][4]  ( .D(n8222), .E(n912), .CK(clk), .Q(
        \registers[982][4] ) );
  EDFFX1 \registers_reg[982][3]  ( .D(n8174), .E(n912), .CK(clk), .Q(
        \registers[982][3] ) );
  EDFFX1 \registers_reg[982][2]  ( .D(n8123), .E(n912), .CK(clk), .Q(
        \registers[982][2] ) );
  EDFFX1 \registers_reg[982][1]  ( .D(n8067), .E(n912), .CK(clk), .Q(
        \registers[982][1] ) );
  EDFFX1 \registers_reg[982][0]  ( .D(n8009), .E(n912), .CK(clk), .Q(
        \registers[982][0] ) );
  EDFFX1 \registers_reg[978][7]  ( .D(n8392), .E(n225), .CK(clk), .Q(
        \registers[978][7] ) );
  EDFFX1 \registers_reg[978][6]  ( .D(n8334), .E(n225), .CK(clk), .Q(
        \registers[978][6] ) );
  EDFFX1 \registers_reg[978][5]  ( .D(n8276), .E(n225), .CK(clk), .Q(
        \registers[978][5] ) );
  EDFFX1 \registers_reg[978][4]  ( .D(n8218), .E(n225), .CK(clk), .Q(
        \registers[978][4] ) );
  EDFFX1 \registers_reg[978][3]  ( .D(n8175), .E(n225), .CK(clk), .Q(
        \registers[978][3] ) );
  EDFFX1 \registers_reg[978][2]  ( .D(n8124), .E(n225), .CK(clk), .Q(
        \registers[978][2] ) );
  EDFFX1 \registers_reg[978][1]  ( .D(n8068), .E(n225), .CK(clk), .Q(
        \registers[978][1] ) );
  EDFFX1 \registers_reg[978][0]  ( .D(n8007), .E(n225), .CK(clk), .Q(
        \registers[978][0] ) );
  EDFFX1 \registers_reg[974][7]  ( .D(n8393), .E(n221), .CK(clk), .Q(
        \registers[974][7] ) );
  EDFFX1 \registers_reg[974][6]  ( .D(n8335), .E(n221), .CK(clk), .Q(
        \registers[974][6] ) );
  EDFFX1 \registers_reg[974][5]  ( .D(n8277), .E(n221), .CK(clk), .Q(
        \registers[974][5] ) );
  EDFFX1 \registers_reg[974][4]  ( .D(n8219), .E(n221), .CK(clk), .Q(
        \registers[974][4] ) );
  EDFFX1 \registers_reg[974][3]  ( .D(n8173), .E(n221), .CK(clk), .Q(
        \registers[974][3] ) );
  EDFFX1 \registers_reg[974][2]  ( .D(n8125), .E(n221), .CK(clk), .Q(
        \registers[974][2] ) );
  EDFFX1 \registers_reg[974][1]  ( .D(n8069), .E(n221), .CK(clk), .Q(
        \registers[974][1] ) );
  EDFFX1 \registers_reg[974][0]  ( .D(n8008), .E(n221), .CK(clk), .Q(
        \registers[974][0] ) );
  EDFFX1 \registers_reg[970][7]  ( .D(n8394), .E(n217), .CK(clk), .Q(
        \registers[970][7] ) );
  EDFFX1 \registers_reg[970][6]  ( .D(n8336), .E(n217), .CK(clk), .Q(
        \registers[970][6] ) );
  EDFFX1 \registers_reg[970][5]  ( .D(n8278), .E(n217), .CK(clk), .Q(
        \registers[970][5] ) );
  EDFFX1 \registers_reg[970][4]  ( .D(n8220), .E(n217), .CK(clk), .Q(
        \registers[970][4] ) );
  EDFFX1 \registers_reg[970][3]  ( .D(n8174), .E(n217), .CK(clk), .Q(
        \registers[970][3] ) );
  EDFFX1 \registers_reg[970][2]  ( .D(n8123), .E(n217), .CK(clk), .Q(
        \registers[970][2] ) );
  EDFFX1 \registers_reg[970][1]  ( .D(n8067), .E(n217), .CK(clk), .Q(
        \registers[970][1] ) );
  EDFFX1 \registers_reg[970][0]  ( .D(n8009), .E(n217), .CK(clk), .Q(
        \registers[970][0] ) );
  EDFFX1 \registers_reg[966][7]  ( .D(n8392), .E(n378), .CK(clk), .Q(
        \registers[966][7] ) );
  EDFFX1 \registers_reg[966][6]  ( .D(n8334), .E(n378), .CK(clk), .Q(
        \registers[966][6] ) );
  EDFFX1 \registers_reg[966][5]  ( .D(n8276), .E(n378), .CK(clk), .Q(
        \registers[966][5] ) );
  EDFFX1 \registers_reg[966][4]  ( .D(n8218), .E(n378), .CK(clk), .Q(
        \registers[966][4] ) );
  EDFFX1 \registers_reg[966][3]  ( .D(n8175), .E(n378), .CK(clk), .Q(
        \registers[966][3] ) );
  EDFFX1 \registers_reg[966][2]  ( .D(n8124), .E(n378), .CK(clk), .Q(
        \registers[966][2] ) );
  EDFFX1 \registers_reg[966][1]  ( .D(n8068), .E(n378), .CK(clk), .Q(
        \registers[966][1] ) );
  EDFFX1 \registers_reg[966][0]  ( .D(n8007), .E(n378), .CK(clk), .Q(
        \registers[966][0] ) );
  EDFFX1 \registers_reg[962][7]  ( .D(n8393), .E(n374), .CK(clk), .Q(
        \registers[962][7] ) );
  EDFFX1 \registers_reg[962][6]  ( .D(n8335), .E(n374), .CK(clk), .Q(
        \registers[962][6] ) );
  EDFFX1 \registers_reg[962][5]  ( .D(n8277), .E(n374), .CK(clk), .Q(
        \registers[962][5] ) );
  EDFFX1 \registers_reg[962][4]  ( .D(n8219), .E(n374), .CK(clk), .Q(
        \registers[962][4] ) );
  EDFFX1 \registers_reg[962][3]  ( .D(n8173), .E(n374), .CK(clk), .Q(
        \registers[962][3] ) );
  EDFFX1 \registers_reg[962][2]  ( .D(n8125), .E(n374), .CK(clk), .Q(
        \registers[962][2] ) );
  EDFFX1 \registers_reg[962][1]  ( .D(n8069), .E(n374), .CK(clk), .Q(
        \registers[962][1] ) );
  EDFFX1 \registers_reg[962][0]  ( .D(n8008), .E(n374), .CK(clk), .Q(
        \registers[962][0] ) );
  EDFFX1 \registers_reg[958][7]  ( .D(n8394), .E(n908), .CK(clk), .Q(
        \registers[958][7] ) );
  EDFFX1 \registers_reg[958][6]  ( .D(n8336), .E(n908), .CK(clk), .Q(
        \registers[958][6] ) );
  EDFFX1 \registers_reg[958][5]  ( .D(n8278), .E(n908), .CK(clk), .Q(
        \registers[958][5] ) );
  EDFFX1 \registers_reg[958][4]  ( .D(n8220), .E(n908), .CK(clk), .Q(
        \registers[958][4] ) );
  EDFFX1 \registers_reg[958][3]  ( .D(n8174), .E(n908), .CK(clk), .Q(
        \registers[958][3] ) );
  EDFFX1 \registers_reg[958][2]  ( .D(n8123), .E(n908), .CK(clk), .Q(
        \registers[958][2] ) );
  EDFFX1 \registers_reg[958][1]  ( .D(n8067), .E(n908), .CK(clk), .Q(
        \registers[958][1] ) );
  EDFFX1 \registers_reg[958][0]  ( .D(n8009), .E(n908), .CK(clk), .Q(
        \registers[958][0] ) );
  EDFFX1 \registers_reg[954][7]  ( .D(n8393), .E(n904), .CK(clk), .Q(
        \registers[954][7] ) );
  EDFFX1 \registers_reg[954][6]  ( .D(n8335), .E(n904), .CK(clk), .Q(
        \registers[954][6] ) );
  EDFFX1 \registers_reg[954][5]  ( .D(n8277), .E(n904), .CK(clk), .Q(
        \registers[954][5] ) );
  EDFFX1 \registers_reg[954][4]  ( .D(n8219), .E(n904), .CK(clk), .Q(
        \registers[954][4] ) );
  EDFFX1 \registers_reg[954][3]  ( .D(n8173), .E(n904), .CK(clk), .Q(
        \registers[954][3] ) );
  EDFFX1 \registers_reg[954][2]  ( .D(n8125), .E(n904), .CK(clk), .Q(
        \registers[954][2] ) );
  EDFFX1 \registers_reg[954][1]  ( .D(n8069), .E(n904), .CK(clk), .Q(
        \registers[954][1] ) );
  EDFFX1 \registers_reg[954][0]  ( .D(n8008), .E(n904), .CK(clk), .Q(
        \registers[954][0] ) );
  EDFFX1 \registers_reg[950][7]  ( .D(n8394), .E(n900), .CK(clk), .Q(
        \registers[950][7] ) );
  EDFFX1 \registers_reg[950][6]  ( .D(n8336), .E(n900), .CK(clk), .Q(
        \registers[950][6] ) );
  EDFFX1 \registers_reg[950][5]  ( .D(n8278), .E(n900), .CK(clk), .Q(
        \registers[950][5] ) );
  EDFFX1 \registers_reg[950][4]  ( .D(n8220), .E(n900), .CK(clk), .Q(
        \registers[950][4] ) );
  EDFFX1 \registers_reg[950][3]  ( .D(n8174), .E(n900), .CK(clk), .Q(
        \registers[950][3] ) );
  EDFFX1 \registers_reg[950][2]  ( .D(n8123), .E(n900), .CK(clk), .Q(
        \registers[950][2] ) );
  EDFFX1 \registers_reg[950][1]  ( .D(n8067), .E(n900), .CK(clk), .Q(
        \registers[950][1] ) );
  EDFFX1 \registers_reg[950][0]  ( .D(n8009), .E(n900), .CK(clk), .Q(
        \registers[950][0] ) );
  EDFFX1 \registers_reg[946][7]  ( .D(n8392), .E(n213), .CK(clk), .Q(
        \registers[946][7] ) );
  EDFFX1 \registers_reg[946][6]  ( .D(n8334), .E(n213), .CK(clk), .Q(
        \registers[946][6] ) );
  EDFFX1 \registers_reg[946][5]  ( .D(n8276), .E(n213), .CK(clk), .Q(
        \registers[946][5] ) );
  EDFFX1 \registers_reg[946][4]  ( .D(n8218), .E(n213), .CK(clk), .Q(
        \registers[946][4] ) );
  EDFFX1 \registers_reg[946][3]  ( .D(n8175), .E(n213), .CK(clk), .Q(
        \registers[946][3] ) );
  EDFFX1 \registers_reg[946][2]  ( .D(n8124), .E(n213), .CK(clk), .Q(
        \registers[946][2] ) );
  EDFFX1 \registers_reg[946][1]  ( .D(n8068), .E(n213), .CK(clk), .Q(
        \registers[946][1] ) );
  EDFFX1 \registers_reg[946][0]  ( .D(n8007), .E(n213), .CK(clk), .Q(
        \registers[946][0] ) );
  EDFFX1 \registers_reg[942][7]  ( .D(n8393), .E(n209), .CK(clk), .Q(
        \registers[942][7] ) );
  EDFFX1 \registers_reg[942][6]  ( .D(n8335), .E(n209), .CK(clk), .Q(
        \registers[942][6] ) );
  EDFFX1 \registers_reg[942][5]  ( .D(n8277), .E(n209), .CK(clk), .Q(
        \registers[942][5] ) );
  EDFFX1 \registers_reg[942][4]  ( .D(n8219), .E(n209), .CK(clk), .Q(
        \registers[942][4] ) );
  EDFFX1 \registers_reg[942][3]  ( .D(n8170), .E(n209), .CK(clk), .Q(
        \registers[942][3] ) );
  EDFFX1 \registers_reg[942][2]  ( .D(n8125), .E(n209), .CK(clk), .Q(
        \registers[942][2] ) );
  EDFFX1 \registers_reg[942][1]  ( .D(n8069), .E(n209), .CK(clk), .Q(
        \registers[942][1] ) );
  EDFFX1 \registers_reg[942][0]  ( .D(n8008), .E(n209), .CK(clk), .Q(
        \registers[942][0] ) );
  EDFFX1 \registers_reg[938][7]  ( .D(n8394), .E(n205), .CK(clk), .Q(
        \registers[938][7] ) );
  EDFFX1 \registers_reg[938][6]  ( .D(n8336), .E(n205), .CK(clk), .Q(
        \registers[938][6] ) );
  EDFFX1 \registers_reg[938][5]  ( .D(n8278), .E(n205), .CK(clk), .Q(
        \registers[938][5] ) );
  EDFFX1 \registers_reg[938][4]  ( .D(n8220), .E(n205), .CK(clk), .Q(
        \registers[938][4] ) );
  EDFFX1 \registers_reg[938][3]  ( .D(n8171), .E(n205), .CK(clk), .Q(
        \registers[938][3] ) );
  EDFFX1 \registers_reg[938][2]  ( .D(n8123), .E(n205), .CK(clk), .Q(
        \registers[938][2] ) );
  EDFFX1 \registers_reg[938][1]  ( .D(n8067), .E(n205), .CK(clk), .Q(
        \registers[938][1] ) );
  EDFFX1 \registers_reg[938][0]  ( .D(n8009), .E(n205), .CK(clk), .Q(
        \registers[938][0] ) );
  EDFFX1 \registers_reg[934][7]  ( .D(n8392), .E(n371), .CK(clk), .Q(
        \registers[934][7] ) );
  EDFFX1 \registers_reg[934][6]  ( .D(n8334), .E(n371), .CK(clk), .Q(
        \registers[934][6] ) );
  EDFFX1 \registers_reg[934][5]  ( .D(n8276), .E(n371), .CK(clk), .Q(
        \registers[934][5] ) );
  EDFFX1 \registers_reg[934][4]  ( .D(n8218), .E(n371), .CK(clk), .Q(
        \registers[934][4] ) );
  EDFFX1 \registers_reg[934][3]  ( .D(n8172), .E(n371), .CK(clk), .Q(
        \registers[934][3] ) );
  EDFFX1 \registers_reg[934][2]  ( .D(n8121), .E(n371), .CK(clk), .Q(
        \registers[934][2] ) );
  EDFFX1 \registers_reg[934][1]  ( .D(n8065), .E(n371), .CK(clk), .Q(
        \registers[934][1] ) );
  EDFFX1 \registers_reg[934][0]  ( .D(n8004), .E(n371), .CK(clk), .Q(
        \registers[934][0] ) );
  EDFFX1 \registers_reg[930][7]  ( .D(n8393), .E(n367), .CK(clk), .Q(
        \registers[930][7] ) );
  EDFFX1 \registers_reg[930][6]  ( .D(n8335), .E(n367), .CK(clk), .Q(
        \registers[930][6] ) );
  EDFFX1 \registers_reg[930][5]  ( .D(n8277), .E(n367), .CK(clk), .Q(
        \registers[930][5] ) );
  EDFFX1 \registers_reg[930][4]  ( .D(n8219), .E(n367), .CK(clk), .Q(
        \registers[930][4] ) );
  EDFFX1 \registers_reg[930][3]  ( .D(n8170), .E(n367), .CK(clk), .Q(
        \registers[930][3] ) );
  EDFFX1 \registers_reg[930][2]  ( .D(n8122), .E(n367), .CK(clk), .Q(
        \registers[930][2] ) );
  EDFFX1 \registers_reg[930][1]  ( .D(n8066), .E(n367), .CK(clk), .Q(
        \registers[930][1] ) );
  EDFFX1 \registers_reg[930][0]  ( .D(n8005), .E(n367), .CK(clk), .Q(
        \registers[930][0] ) );
  EDFFX1 \registers_reg[926][7]  ( .D(n8389), .E(n896), .CK(clk), .Q(
        \registers[926][7] ) );
  EDFFX1 \registers_reg[926][6]  ( .D(n8331), .E(n896), .CK(clk), .Q(
        \registers[926][6] ) );
  EDFFX1 \registers_reg[926][5]  ( .D(n8273), .E(n896), .CK(clk), .Q(
        \registers[926][5] ) );
  EDFFX1 \registers_reg[926][4]  ( .D(n8215), .E(n896), .CK(clk), .Q(
        \registers[926][4] ) );
  EDFFX1 \registers_reg[926][3]  ( .D(n8171), .E(n896), .CK(clk), .Q(
        \registers[926][3] ) );
  EDFFX1 \registers_reg[926][2]  ( .D(n8120), .E(n896), .CK(clk), .Q(
        \registers[926][2] ) );
  EDFFX1 \registers_reg[926][1]  ( .D(n8064), .E(n896), .CK(clk), .Q(
        \registers[926][1] ) );
  EDFFX1 \registers_reg[926][0]  ( .D(n8006), .E(n896), .CK(clk), .Q(
        \registers[926][0] ) );
  EDFFX1 \registers_reg[922][7]  ( .D(n8390), .E(n892), .CK(clk), .Q(
        \registers[922][7] ) );
  EDFFX1 \registers_reg[922][6]  ( .D(n8332), .E(n892), .CK(clk), .Q(
        \registers[922][6] ) );
  EDFFX1 \registers_reg[922][5]  ( .D(n8274), .E(n892), .CK(clk), .Q(
        \registers[922][5] ) );
  EDFFX1 \registers_reg[922][4]  ( .D(n8216), .E(n892), .CK(clk), .Q(
        \registers[922][4] ) );
  EDFFX1 \registers_reg[922][3]  ( .D(n8172), .E(n892), .CK(clk), .Q(
        \registers[922][3] ) );
  EDFFX1 \registers_reg[922][2]  ( .D(n8121), .E(n892), .CK(clk), .Q(
        \registers[922][2] ) );
  EDFFX1 \registers_reg[922][1]  ( .D(n8065), .E(n892), .CK(clk), .Q(
        \registers[922][1] ) );
  EDFFX1 \registers_reg[922][0]  ( .D(n8004), .E(n892), .CK(clk), .Q(
        \registers[922][0] ) );
  EDFFX1 \registers_reg[918][7]  ( .D(n8391), .E(n888), .CK(clk), .Q(
        \registers[918][7] ) );
  EDFFX1 \registers_reg[918][6]  ( .D(n8333), .E(n888), .CK(clk), .Q(
        \registers[918][6] ) );
  EDFFX1 \registers_reg[918][5]  ( .D(n8275), .E(n888), .CK(clk), .Q(
        \registers[918][5] ) );
  EDFFX1 \registers_reg[918][4]  ( .D(n8217), .E(n888), .CK(clk), .Q(
        \registers[918][4] ) );
  EDFFX1 \registers_reg[918][3]  ( .D(n8170), .E(n888), .CK(clk), .Q(
        \registers[918][3] ) );
  EDFFX1 \registers_reg[918][2]  ( .D(n8122), .E(n888), .CK(clk), .Q(
        \registers[918][2] ) );
  EDFFX1 \registers_reg[918][1]  ( .D(n8066), .E(n888), .CK(clk), .Q(
        \registers[918][1] ) );
  EDFFX1 \registers_reg[918][0]  ( .D(n8005), .E(n888), .CK(clk), .Q(
        \registers[918][0] ) );
  EDFFX1 \registers_reg[914][7]  ( .D(n8389), .E(n201), .CK(clk), .Q(
        \registers[914][7] ) );
  EDFFX1 \registers_reg[914][6]  ( .D(n8331), .E(n201), .CK(clk), .Q(
        \registers[914][6] ) );
  EDFFX1 \registers_reg[914][5]  ( .D(n8273), .E(n201), .CK(clk), .Q(
        \registers[914][5] ) );
  EDFFX1 \registers_reg[914][4]  ( .D(n8215), .E(n201), .CK(clk), .Q(
        \registers[914][4] ) );
  EDFFX1 \registers_reg[914][3]  ( .D(n8171), .E(n201), .CK(clk), .Q(
        \registers[914][3] ) );
  EDFFX1 \registers_reg[914][2]  ( .D(n8120), .E(n201), .CK(clk), .Q(
        \registers[914][2] ) );
  EDFFX1 \registers_reg[914][1]  ( .D(n8064), .E(n201), .CK(clk), .Q(
        \registers[914][1] ) );
  EDFFX1 \registers_reg[914][0]  ( .D(n8006), .E(n201), .CK(clk), .Q(
        \registers[914][0] ) );
  EDFFX1 \registers_reg[910][7]  ( .D(n8390), .E(n197), .CK(clk), .Q(
        \registers[910][7] ) );
  EDFFX1 \registers_reg[910][6]  ( .D(n8332), .E(n197), .CK(clk), .Q(
        \registers[910][6] ) );
  EDFFX1 \registers_reg[910][5]  ( .D(n8274), .E(n197), .CK(clk), .Q(
        \registers[910][5] ) );
  EDFFX1 \registers_reg[910][4]  ( .D(n8216), .E(n197), .CK(clk), .Q(
        \registers[910][4] ) );
  EDFFX1 \registers_reg[910][3]  ( .D(n8172), .E(n197), .CK(clk), .Q(
        \registers[910][3] ) );
  EDFFX1 \registers_reg[910][2]  ( .D(n8121), .E(n197), .CK(clk), .Q(
        \registers[910][2] ) );
  EDFFX1 \registers_reg[910][1]  ( .D(n8065), .E(n197), .CK(clk), .Q(
        \registers[910][1] ) );
  EDFFX1 \registers_reg[910][0]  ( .D(n8004), .E(n197), .CK(clk), .Q(
        \registers[910][0] ) );
  EDFFX1 \registers_reg[906][7]  ( .D(n8391), .E(n193), .CK(clk), .Q(
        \registers[906][7] ) );
  EDFFX1 \registers_reg[906][6]  ( .D(n8333), .E(n193), .CK(clk), .Q(
        \registers[906][6] ) );
  EDFFX1 \registers_reg[906][5]  ( .D(n8275), .E(n193), .CK(clk), .Q(
        \registers[906][5] ) );
  EDFFX1 \registers_reg[906][4]  ( .D(n8217), .E(n193), .CK(clk), .Q(
        \registers[906][4] ) );
  EDFFX1 \registers_reg[906][3]  ( .D(n8170), .E(n193), .CK(clk), .Q(
        \registers[906][3] ) );
  EDFFX1 \registers_reg[906][2]  ( .D(n8122), .E(n193), .CK(clk), .Q(
        \registers[906][2] ) );
  EDFFX1 \registers_reg[906][1]  ( .D(n8066), .E(n193), .CK(clk), .Q(
        \registers[906][1] ) );
  EDFFX1 \registers_reg[906][0]  ( .D(n8005), .E(n193), .CK(clk), .Q(
        \registers[906][0] ) );
  EDFFX1 \registers_reg[902][7]  ( .D(n8389), .E(n364), .CK(clk), .Q(
        \registers[902][7] ) );
  EDFFX1 \registers_reg[902][6]  ( .D(n8331), .E(n364), .CK(clk), .Q(
        \registers[902][6] ) );
  EDFFX1 \registers_reg[902][5]  ( .D(n8273), .E(n364), .CK(clk), .Q(
        \registers[902][5] ) );
  EDFFX1 \registers_reg[902][4]  ( .D(n8215), .E(n364), .CK(clk), .Q(
        \registers[902][4] ) );
  EDFFX1 \registers_reg[902][3]  ( .D(n8171), .E(n364), .CK(clk), .Q(
        \registers[902][3] ) );
  EDFFX1 \registers_reg[902][2]  ( .D(n8120), .E(n364), .CK(clk), .Q(
        \registers[902][2] ) );
  EDFFX1 \registers_reg[902][1]  ( .D(n8064), .E(n364), .CK(clk), .Q(
        \registers[902][1] ) );
  EDFFX1 \registers_reg[902][0]  ( .D(n8006), .E(n364), .CK(clk), .Q(
        \registers[902][0] ) );
  EDFFX1 \registers_reg[898][7]  ( .D(n8390), .E(n360), .CK(clk), .Q(
        \registers[898][7] ) );
  EDFFX1 \registers_reg[898][6]  ( .D(n8332), .E(n360), .CK(clk), .Q(
        \registers[898][6] ) );
  EDFFX1 \registers_reg[898][5]  ( .D(n8274), .E(n360), .CK(clk), .Q(
        \registers[898][5] ) );
  EDFFX1 \registers_reg[898][4]  ( .D(n8216), .E(n360), .CK(clk), .Q(
        \registers[898][4] ) );
  EDFFX1 \registers_reg[898][3]  ( .D(n8172), .E(n360), .CK(clk), .Q(
        \registers[898][3] ) );
  EDFFX1 \registers_reg[898][2]  ( .D(n8121), .E(n360), .CK(clk), .Q(
        \registers[898][2] ) );
  EDFFX1 \registers_reg[898][1]  ( .D(n8065), .E(n360), .CK(clk), .Q(
        \registers[898][1] ) );
  EDFFX1 \registers_reg[898][0]  ( .D(n8004), .E(n360), .CK(clk), .Q(
        \registers[898][0] ) );
  EDFFX1 \registers_reg[894][7]  ( .D(n8392), .E(n884), .CK(clk), .Q(
        \registers[894][7] ) );
  EDFFX1 \registers_reg[894][6]  ( .D(n8334), .E(n884), .CK(clk), .Q(
        \registers[894][6] ) );
  EDFFX1 \registers_reg[894][5]  ( .D(n8276), .E(n884), .CK(clk), .Q(
        \registers[894][5] ) );
  EDFFX1 \registers_reg[894][4]  ( .D(n8218), .E(n884), .CK(clk), .Q(
        \registers[894][4] ) );
  EDFFX1 \registers_reg[894][3]  ( .D(n8175), .E(n884), .CK(clk), .Q(
        \registers[894][3] ) );
  EDFFX1 \registers_reg[894][2]  ( .D(n8124), .E(n884), .CK(clk), .Q(
        \registers[894][2] ) );
  EDFFX1 \registers_reg[894][1]  ( .D(n8068), .E(n884), .CK(clk), .Q(
        \registers[894][1] ) );
  EDFFX1 \registers_reg[894][0]  ( .D(n8007), .E(n884), .CK(clk), .Q(
        \registers[894][0] ) );
  EDFFX1 \registers_reg[890][7]  ( .D(n8404), .E(n880), .CK(clk), .Q(
        \registers[890][7] ) );
  EDFFX1 \registers_reg[890][6]  ( .D(n8346), .E(n880), .CK(clk), .Q(
        \registers[890][6] ) );
  EDFFX1 \registers_reg[890][5]  ( .D(n8288), .E(n880), .CK(clk), .Q(
        \registers[890][5] ) );
  EDFFX1 \registers_reg[890][4]  ( .D(n8230), .E(n880), .CK(clk), .Q(
        \registers[890][4] ) );
  EDFFX1 \registers_reg[890][3]  ( .D(n8182), .E(n880), .CK(clk), .Q(
        \registers[890][3] ) );
  EDFFX1 \registers_reg[890][2]  ( .D(n8137), .E(n880), .CK(clk), .Q(
        \registers[890][2] ) );
  EDFFX1 \registers_reg[890][1]  ( .D(n8081), .E(n880), .CK(clk), .Q(
        \registers[890][1] ) );
  EDFFX1 \registers_reg[890][0]  ( .D(n8020), .E(n880), .CK(clk), .Q(
        \registers[890][0] ) );
  EDFFX1 \registers_reg[886][7]  ( .D(n8405), .E(n876), .CK(clk), .Q(
        \registers[886][7] ) );
  EDFFX1 \registers_reg[886][6]  ( .D(n8347), .E(n876), .CK(clk), .Q(
        \registers[886][6] ) );
  EDFFX1 \registers_reg[886][5]  ( .D(n8289), .E(n876), .CK(clk), .Q(
        \registers[886][5] ) );
  EDFFX1 \registers_reg[886][4]  ( .D(n8231), .E(n876), .CK(clk), .Q(
        \registers[886][4] ) );
  EDFFX1 \registers_reg[886][3]  ( .D(n8183), .E(n876), .CK(clk), .Q(
        \registers[886][3] ) );
  EDFFX1 \registers_reg[886][2]  ( .D(n8135), .E(n876), .CK(clk), .Q(
        \registers[886][2] ) );
  EDFFX1 \registers_reg[886][1]  ( .D(n8079), .E(n876), .CK(clk), .Q(
        \registers[886][1] ) );
  EDFFX1 \registers_reg[886][0]  ( .D(n8021), .E(n876), .CK(clk), .Q(
        \registers[886][0] ) );
  EDFFX1 \registers_reg[882][7]  ( .D(n8406), .E(n189), .CK(clk), .Q(
        \registers[882][7] ) );
  EDFFX1 \registers_reg[882][6]  ( .D(n8348), .E(n189), .CK(clk), .Q(
        \registers[882][6] ) );
  EDFFX1 \registers_reg[882][5]  ( .D(n8290), .E(n189), .CK(clk), .Q(
        \registers[882][5] ) );
  EDFFX1 \registers_reg[882][4]  ( .D(n8232), .E(n189), .CK(clk), .Q(
        \registers[882][4] ) );
  EDFFX1 \registers_reg[882][3]  ( .D(n8184), .E(n189), .CK(clk), .Q(
        \registers[882][3] ) );
  EDFFX1 \registers_reg[882][2]  ( .D(n8133), .E(n189), .CK(clk), .Q(
        \registers[882][2] ) );
  EDFFX1 \registers_reg[882][1]  ( .D(n8077), .E(n189), .CK(clk), .Q(
        \registers[882][1] ) );
  EDFFX1 \registers_reg[882][0]  ( .D(n8016), .E(n189), .CK(clk), .Q(
        \registers[882][0] ) );
  EDFFX1 \registers_reg[878][7]  ( .D(n8404), .E(n185), .CK(clk), .Q(
        \registers[878][7] ) );
  EDFFX1 \registers_reg[878][6]  ( .D(n8346), .E(n185), .CK(clk), .Q(
        \registers[878][6] ) );
  EDFFX1 \registers_reg[878][5]  ( .D(n8288), .E(n185), .CK(clk), .Q(
        \registers[878][5] ) );
  EDFFX1 \registers_reg[878][4]  ( .D(n8230), .E(n185), .CK(clk), .Q(
        \registers[878][4] ) );
  EDFFX1 \registers_reg[878][3]  ( .D(n8182), .E(n185), .CK(clk), .Q(
        \registers[878][3] ) );
  EDFFX1 \registers_reg[878][2]  ( .D(n8134), .E(n185), .CK(clk), .Q(
        \registers[878][2] ) );
  EDFFX1 \registers_reg[878][1]  ( .D(n8078), .E(n185), .CK(clk), .Q(
        \registers[878][1] ) );
  EDFFX1 \registers_reg[878][0]  ( .D(n8017), .E(n185), .CK(clk), .Q(
        \registers[878][0] ) );
  EDFFX1 \registers_reg[874][7]  ( .D(n8405), .E(n181), .CK(clk), .Q(
        \registers[874][7] ) );
  EDFFX1 \registers_reg[874][6]  ( .D(n8347), .E(n181), .CK(clk), .Q(
        \registers[874][6] ) );
  EDFFX1 \registers_reg[874][5]  ( .D(n8289), .E(n181), .CK(clk), .Q(
        \registers[874][5] ) );
  EDFFX1 \registers_reg[874][4]  ( .D(n8231), .E(n181), .CK(clk), .Q(
        \registers[874][4] ) );
  EDFFX1 \registers_reg[874][3]  ( .D(n8180), .E(n181), .CK(clk), .Q(
        \registers[874][3] ) );
  EDFFX1 \registers_reg[874][2]  ( .D(n8132), .E(n181), .CK(clk), .Q(
        \registers[874][2] ) );
  EDFFX1 \registers_reg[874][1]  ( .D(n8076), .E(n181), .CK(clk), .Q(
        \registers[874][1] ) );
  EDFFX1 \registers_reg[874][0]  ( .D(n8018), .E(n181), .CK(clk), .Q(
        \registers[874][0] ) );
  EDFFX1 \registers_reg[870][7]  ( .D(n8401), .E(n357), .CK(clk), .Q(
        \registers[870][7] ) );
  EDFFX1 \registers_reg[870][6]  ( .D(n8343), .E(n357), .CK(clk), .Q(
        \registers[870][6] ) );
  EDFFX1 \registers_reg[870][5]  ( .D(n8285), .E(n357), .CK(clk), .Q(
        \registers[870][5] ) );
  EDFFX1 \registers_reg[870][4]  ( .D(n8227), .E(n357), .CK(clk), .Q(
        \registers[870][4] ) );
  EDFFX1 \registers_reg[870][3]  ( .D(n8181), .E(n357), .CK(clk), .Q(
        \registers[870][3] ) );
  EDFFX1 \registers_reg[870][2]  ( .D(n8133), .E(n357), .CK(clk), .Q(
        \registers[870][2] ) );
  EDFFX1 \registers_reg[870][1]  ( .D(n8077), .E(n357), .CK(clk), .Q(
        \registers[870][1] ) );
  EDFFX1 \registers_reg[870][0]  ( .D(n8016), .E(n357), .CK(clk), .Q(
        \registers[870][0] ) );
  EDFFX1 \registers_reg[866][7]  ( .D(n8402), .E(n353), .CK(clk), .Q(
        \registers[866][7] ) );
  EDFFX1 \registers_reg[866][6]  ( .D(n8344), .E(n353), .CK(clk), .Q(
        \registers[866][6] ) );
  EDFFX1 \registers_reg[866][5]  ( .D(n8286), .E(n353), .CK(clk), .Q(
        \registers[866][5] ) );
  EDFFX1 \registers_reg[866][4]  ( .D(n8228), .E(n353), .CK(clk), .Q(
        \registers[866][4] ) );
  EDFFX1 \registers_reg[866][3]  ( .D(n8179), .E(n353), .CK(clk), .Q(
        \registers[866][3] ) );
  EDFFX1 \registers_reg[866][2]  ( .D(n8134), .E(n353), .CK(clk), .Q(
        \registers[866][2] ) );
  EDFFX1 \registers_reg[866][1]  ( .D(n8078), .E(n353), .CK(clk), .Q(
        \registers[866][1] ) );
  EDFFX1 \registers_reg[866][0]  ( .D(n8017), .E(n353), .CK(clk), .Q(
        \registers[866][0] ) );
  EDFFX1 \registers_reg[862][7]  ( .D(n8403), .E(n872), .CK(clk), .Q(
        \registers[862][7] ) );
  EDFFX1 \registers_reg[862][6]  ( .D(n8345), .E(n872), .CK(clk), .Q(
        \registers[862][6] ) );
  EDFFX1 \registers_reg[862][5]  ( .D(n8287), .E(n872), .CK(clk), .Q(
        \registers[862][5] ) );
  EDFFX1 \registers_reg[862][4]  ( .D(n8229), .E(n872), .CK(clk), .Q(
        \registers[862][4] ) );
  EDFFX1 \registers_reg[862][3]  ( .D(n8180), .E(n872), .CK(clk), .Q(
        \registers[862][3] ) );
  EDFFX1 \registers_reg[862][2]  ( .D(n8132), .E(n872), .CK(clk), .Q(
        \registers[862][2] ) );
  EDFFX1 \registers_reg[862][1]  ( .D(n8076), .E(n872), .CK(clk), .Q(
        \registers[862][1] ) );
  EDFFX1 \registers_reg[862][0]  ( .D(n8018), .E(n872), .CK(clk), .Q(
        \registers[862][0] ) );
  EDFFX1 \registers_reg[858][7]  ( .D(n8401), .E(n868), .CK(clk), .Q(
        \registers[858][7] ) );
  EDFFX1 \registers_reg[858][6]  ( .D(n8343), .E(n868), .CK(clk), .Q(
        \registers[858][6] ) );
  EDFFX1 \registers_reg[858][5]  ( .D(n8285), .E(n868), .CK(clk), .Q(
        \registers[858][5] ) );
  EDFFX1 \registers_reg[858][4]  ( .D(n8227), .E(n868), .CK(clk), .Q(
        \registers[858][4] ) );
  EDFFX1 \registers_reg[858][3]  ( .D(n8181), .E(n868), .CK(clk), .Q(
        \registers[858][3] ) );
  EDFFX1 \registers_reg[858][2]  ( .D(n8133), .E(n868), .CK(clk), .Q(
        \registers[858][2] ) );
  EDFFX1 \registers_reg[858][1]  ( .D(n8077), .E(n868), .CK(clk), .Q(
        \registers[858][1] ) );
  EDFFX1 \registers_reg[858][0]  ( .D(n8016), .E(n868), .CK(clk), .Q(
        \registers[858][0] ) );
  EDFFX1 \registers_reg[854][7]  ( .D(n8402), .E(n864), .CK(clk), .Q(
        \registers[854][7] ) );
  EDFFX1 \registers_reg[854][6]  ( .D(n8344), .E(n864), .CK(clk), .Q(
        \registers[854][6] ) );
  EDFFX1 \registers_reg[854][5]  ( .D(n8286), .E(n864), .CK(clk), .Q(
        \registers[854][5] ) );
  EDFFX1 \registers_reg[854][4]  ( .D(n8228), .E(n864), .CK(clk), .Q(
        \registers[854][4] ) );
  EDFFX1 \registers_reg[854][3]  ( .D(n8179), .E(n864), .CK(clk), .Q(
        \registers[854][3] ) );
  EDFFX1 \registers_reg[854][2]  ( .D(n8134), .E(n864), .CK(clk), .Q(
        \registers[854][2] ) );
  EDFFX1 \registers_reg[854][1]  ( .D(n8078), .E(n864), .CK(clk), .Q(
        \registers[854][1] ) );
  EDFFX1 \registers_reg[854][0]  ( .D(n8017), .E(n864), .CK(clk), .Q(
        \registers[854][0] ) );
  EDFFX1 \registers_reg[850][7]  ( .D(n8403), .E(n177), .CK(clk), .Q(
        \registers[850][7] ) );
  EDFFX1 \registers_reg[850][6]  ( .D(n8345), .E(n177), .CK(clk), .Q(
        \registers[850][6] ) );
  EDFFX1 \registers_reg[850][5]  ( .D(n8287), .E(n177), .CK(clk), .Q(
        \registers[850][5] ) );
  EDFFX1 \registers_reg[850][4]  ( .D(n8229), .E(n177), .CK(clk), .Q(
        \registers[850][4] ) );
  EDFFX1 \registers_reg[850][3]  ( .D(n8180), .E(n177), .CK(clk), .Q(
        \registers[850][3] ) );
  EDFFX1 \registers_reg[850][2]  ( .D(n8132), .E(n177), .CK(clk), .Q(
        \registers[850][2] ) );
  EDFFX1 \registers_reg[850][1]  ( .D(n8076), .E(n177), .CK(clk), .Q(
        \registers[850][1] ) );
  EDFFX1 \registers_reg[850][0]  ( .D(n8018), .E(n177), .CK(clk), .Q(
        \registers[850][0] ) );
  EDFFX1 \registers_reg[846][7]  ( .D(n8401), .E(n173), .CK(clk), .Q(
        \registers[846][7] ) );
  EDFFX1 \registers_reg[846][6]  ( .D(n8343), .E(n173), .CK(clk), .Q(
        \registers[846][6] ) );
  EDFFX1 \registers_reg[846][5]  ( .D(n8285), .E(n173), .CK(clk), .Q(
        \registers[846][5] ) );
  EDFFX1 \registers_reg[846][4]  ( .D(n8227), .E(n173), .CK(clk), .Q(
        \registers[846][4] ) );
  EDFFX1 \registers_reg[846][3]  ( .D(n8181), .E(n173), .CK(clk), .Q(
        \registers[846][3] ) );
  EDFFX1 \registers_reg[846][2]  ( .D(n8133), .E(n173), .CK(clk), .Q(
        \registers[846][2] ) );
  EDFFX1 \registers_reg[846][1]  ( .D(n8077), .E(n173), .CK(clk), .Q(
        \registers[846][1] ) );
  EDFFX1 \registers_reg[846][0]  ( .D(n8016), .E(n173), .CK(clk), .Q(
        \registers[846][0] ) );
  EDFFX1 \registers_reg[842][7]  ( .D(n8402), .E(n169), .CK(clk), .Q(
        \registers[842][7] ) );
  EDFFX1 \registers_reg[842][6]  ( .D(n8344), .E(n169), .CK(clk), .Q(
        \registers[842][6] ) );
  EDFFX1 \registers_reg[842][5]  ( .D(n8286), .E(n169), .CK(clk), .Q(
        \registers[842][5] ) );
  EDFFX1 \registers_reg[842][4]  ( .D(n8228), .E(n169), .CK(clk), .Q(
        \registers[842][4] ) );
  EDFFX1 \registers_reg[842][3]  ( .D(n8179), .E(n169), .CK(clk), .Q(
        \registers[842][3] ) );
  EDFFX1 \registers_reg[842][2]  ( .D(n8134), .E(n169), .CK(clk), .Q(
        \registers[842][2] ) );
  EDFFX1 \registers_reg[842][1]  ( .D(n8078), .E(n169), .CK(clk), .Q(
        \registers[842][1] ) );
  EDFFX1 \registers_reg[842][0]  ( .D(n8017), .E(n169), .CK(clk), .Q(
        \registers[842][0] ) );
  EDFFX1 \registers_reg[838][7]  ( .D(n8403), .E(n350), .CK(clk), .Q(
        \registers[838][7] ) );
  EDFFX1 \registers_reg[838][6]  ( .D(n8345), .E(n350), .CK(clk), .Q(
        \registers[838][6] ) );
  EDFFX1 \registers_reg[838][5]  ( .D(n8287), .E(n350), .CK(clk), .Q(
        \registers[838][5] ) );
  EDFFX1 \registers_reg[838][4]  ( .D(n8229), .E(n350), .CK(clk), .Q(
        \registers[838][4] ) );
  EDFFX1 \registers_reg[838][3]  ( .D(n8180), .E(n350), .CK(clk), .Q(
        \registers[838][3] ) );
  EDFFX1 \registers_reg[838][2]  ( .D(n8132), .E(n350), .CK(clk), .Q(
        \registers[838][2] ) );
  EDFFX1 \registers_reg[838][1]  ( .D(n8076), .E(n350), .CK(clk), .Q(
        \registers[838][1] ) );
  EDFFX1 \registers_reg[838][0]  ( .D(n8018), .E(n350), .CK(clk), .Q(
        \registers[838][0] ) );
  EDFFX1 \registers_reg[834][7]  ( .D(n8401), .E(n346), .CK(clk), .Q(
        \registers[834][7] ) );
  EDFFX1 \registers_reg[834][6]  ( .D(n8343), .E(n346), .CK(clk), .Q(
        \registers[834][6] ) );
  EDFFX1 \registers_reg[834][5]  ( .D(n8285), .E(n346), .CK(clk), .Q(
        \registers[834][5] ) );
  EDFFX1 \registers_reg[834][4]  ( .D(n8227), .E(n346), .CK(clk), .Q(
        \registers[834][4] ) );
  EDFFX1 \registers_reg[834][3]  ( .D(n8181), .E(n346), .CK(clk), .Q(
        \registers[834][3] ) );
  EDFFX1 \registers_reg[834][2]  ( .D(n8133), .E(n346), .CK(clk), .Q(
        \registers[834][2] ) );
  EDFFX1 \registers_reg[834][1]  ( .D(n8077), .E(n346), .CK(clk), .Q(
        \registers[834][1] ) );
  EDFFX1 \registers_reg[834][0]  ( .D(n8016), .E(n346), .CK(clk), .Q(
        \registers[834][0] ) );
  EDFFX1 \registers_reg[830][7]  ( .D(n8403), .E(n860), .CK(clk), .Q(
        \registers[830][7] ) );
  EDFFX1 \registers_reg[830][6]  ( .D(n8345), .E(n860), .CK(clk), .Q(
        \registers[830][6] ) );
  EDFFX1 \registers_reg[830][5]  ( .D(n8287), .E(n860), .CK(clk), .Q(
        \registers[830][5] ) );
  EDFFX1 \registers_reg[830][4]  ( .D(n8229), .E(n860), .CK(clk), .Q(
        \registers[830][4] ) );
  EDFFX1 \registers_reg[830][3]  ( .D(n8180), .E(n860), .CK(clk), .Q(
        \registers[830][3] ) );
  EDFFX1 \registers_reg[830][2]  ( .D(n8129), .E(n860), .CK(clk), .Q(
        \registers[830][2] ) );
  EDFFX1 \registers_reg[830][1]  ( .D(n8073), .E(n860), .CK(clk), .Q(
        \registers[830][1] ) );
  EDFFX1 \registers_reg[830][0]  ( .D(n8015), .E(n860), .CK(clk), .Q(
        \registers[830][0] ) );
  EDFFX1 \registers_reg[826][7]  ( .D(n8401), .E(n856), .CK(clk), .Q(
        \registers[826][7] ) );
  EDFFX1 \registers_reg[826][6]  ( .D(n8343), .E(n856), .CK(clk), .Q(
        \registers[826][6] ) );
  EDFFX1 \registers_reg[826][5]  ( .D(n8285), .E(n856), .CK(clk), .Q(
        \registers[826][5] ) );
  EDFFX1 \registers_reg[826][4]  ( .D(n8227), .E(n856), .CK(clk), .Q(
        \registers[826][4] ) );
  EDFFX1 \registers_reg[826][3]  ( .D(n8181), .E(n856), .CK(clk), .Q(
        \registers[826][3] ) );
  EDFFX1 \registers_reg[826][2]  ( .D(n8130), .E(n856), .CK(clk), .Q(
        \registers[826][2] ) );
  EDFFX1 \registers_reg[826][1]  ( .D(n8074), .E(n856), .CK(clk), .Q(
        \registers[826][1] ) );
  EDFFX1 \registers_reg[826][0]  ( .D(n8013), .E(n856), .CK(clk), .Q(
        \registers[826][0] ) );
  EDFFX1 \registers_reg[822][7]  ( .D(n8400), .E(n852), .CK(clk), .Q(
        \registers[822][7] ) );
  EDFFX1 \registers_reg[822][6]  ( .D(n8342), .E(n852), .CK(clk), .Q(
        \registers[822][6] ) );
  EDFFX1 \registers_reg[822][5]  ( .D(n8284), .E(n852), .CK(clk), .Q(
        \registers[822][5] ) );
  EDFFX1 \registers_reg[822][4]  ( .D(n8226), .E(n852), .CK(clk), .Q(
        \registers[822][4] ) );
  EDFFX1 \registers_reg[822][3]  ( .D(n8179), .E(n852), .CK(clk), .Q(
        \registers[822][3] ) );
  EDFFX1 \registers_reg[822][2]  ( .D(n8131), .E(n852), .CK(clk), .Q(
        \registers[822][2] ) );
  EDFFX1 \registers_reg[822][1]  ( .D(n8075), .E(n852), .CK(clk), .Q(
        \registers[822][1] ) );
  EDFFX1 \registers_reg[822][0]  ( .D(n8014), .E(n852), .CK(clk), .Q(
        \registers[822][0] ) );
  EDFFX1 \registers_reg[818][7]  ( .D(n8398), .E(n165), .CK(clk), .Q(
        \registers[818][7] ) );
  EDFFX1 \registers_reg[818][6]  ( .D(n8340), .E(n165), .CK(clk), .Q(
        \registers[818][6] ) );
  EDFFX1 \registers_reg[818][5]  ( .D(n8282), .E(n165), .CK(clk), .Q(
        \registers[818][5] ) );
  EDFFX1 \registers_reg[818][4]  ( .D(n8224), .E(n165), .CK(clk), .Q(
        \registers[818][4] ) );
  EDFFX1 \registers_reg[818][3]  ( .D(n8180), .E(n165), .CK(clk), .Q(
        \registers[818][3] ) );
  EDFFX1 \registers_reg[818][2]  ( .D(n8129), .E(n165), .CK(clk), .Q(
        \registers[818][2] ) );
  EDFFX1 \registers_reg[818][1]  ( .D(n8073), .E(n165), .CK(clk), .Q(
        \registers[818][1] ) );
  EDFFX1 \registers_reg[818][0]  ( .D(n8015), .E(n165), .CK(clk), .Q(
        \registers[818][0] ) );
  EDFFX1 \registers_reg[814][7]  ( .D(n8399), .E(n161), .CK(clk), .Q(
        \registers[814][7] ) );
  EDFFX1 \registers_reg[814][6]  ( .D(n8341), .E(n161), .CK(clk), .Q(
        \registers[814][6] ) );
  EDFFX1 \registers_reg[814][5]  ( .D(n8283), .E(n161), .CK(clk), .Q(
        \registers[814][5] ) );
  EDFFX1 \registers_reg[814][4]  ( .D(n8225), .E(n161), .CK(clk), .Q(
        \registers[814][4] ) );
  EDFFX1 \registers_reg[814][3]  ( .D(n8181), .E(n161), .CK(clk), .Q(
        \registers[814][3] ) );
  EDFFX1 \registers_reg[814][2]  ( .D(n8130), .E(n161), .CK(clk), .Q(
        \registers[814][2] ) );
  EDFFX1 \registers_reg[814][1]  ( .D(n8074), .E(n161), .CK(clk), .Q(
        \registers[814][1] ) );
  EDFFX1 \registers_reg[814][0]  ( .D(n8013), .E(n161), .CK(clk), .Q(
        \registers[814][0] ) );
  EDFFX1 \registers_reg[810][7]  ( .D(n8400), .E(n157), .CK(clk), .Q(
        \registers[810][7] ) );
  EDFFX1 \registers_reg[810][6]  ( .D(n8342), .E(n157), .CK(clk), .Q(
        \registers[810][6] ) );
  EDFFX1 \registers_reg[810][5]  ( .D(n8284), .E(n157), .CK(clk), .Q(
        \registers[810][5] ) );
  EDFFX1 \registers_reg[810][4]  ( .D(n8226), .E(n157), .CK(clk), .Q(
        \registers[810][4] ) );
  EDFFX1 \registers_reg[810][3]  ( .D(n8176), .E(n157), .CK(clk), .Q(
        \registers[810][3] ) );
  EDFFX1 \registers_reg[810][2]  ( .D(n8131), .E(n157), .CK(clk), .Q(
        \registers[810][2] ) );
  EDFFX1 \registers_reg[810][1]  ( .D(n8075), .E(n157), .CK(clk), .Q(
        \registers[810][1] ) );
  EDFFX1 \registers_reg[810][0]  ( .D(n8014), .E(n157), .CK(clk), .Q(
        \registers[810][0] ) );
  EDFFX1 \registers_reg[806][7]  ( .D(n8398), .E(n328), .CK(clk), .Q(
        \registers[806][7] ) );
  EDFFX1 \registers_reg[806][6]  ( .D(n8340), .E(n328), .CK(clk), .Q(
        \registers[806][6] ) );
  EDFFX1 \registers_reg[806][5]  ( .D(n8282), .E(n328), .CK(clk), .Q(
        \registers[806][5] ) );
  EDFFX1 \registers_reg[806][4]  ( .D(n8224), .E(n328), .CK(clk), .Q(
        \registers[806][4] ) );
  EDFFX1 \registers_reg[806][3]  ( .D(n8177), .E(n328), .CK(clk), .Q(
        \registers[806][3] ) );
  EDFFX1 \registers_reg[806][2]  ( .D(n8129), .E(n328), .CK(clk), .Q(
        \registers[806][2] ) );
  EDFFX1 \registers_reg[806][1]  ( .D(n8073), .E(n328), .CK(clk), .Q(
        \registers[806][1] ) );
  EDFFX1 \registers_reg[806][0]  ( .D(n8015), .E(n328), .CK(clk), .Q(
        \registers[806][0] ) );
  EDFFX1 \registers_reg[802][7]  ( .D(n8399), .E(n324), .CK(clk), .Q(
        \registers[802][7] ) );
  EDFFX1 \registers_reg[802][6]  ( .D(n8341), .E(n324), .CK(clk), .Q(
        \registers[802][6] ) );
  EDFFX1 \registers_reg[802][5]  ( .D(n8283), .E(n324), .CK(clk), .Q(
        \registers[802][5] ) );
  EDFFX1 \registers_reg[802][4]  ( .D(n8225), .E(n324), .CK(clk), .Q(
        \registers[802][4] ) );
  EDFFX1 \registers_reg[802][3]  ( .D(n8178), .E(n324), .CK(clk), .Q(
        \registers[802][3] ) );
  EDFFX1 \registers_reg[802][2]  ( .D(n8130), .E(n324), .CK(clk), .Q(
        \registers[802][2] ) );
  EDFFX1 \registers_reg[802][1]  ( .D(n8074), .E(n324), .CK(clk), .Q(
        \registers[802][1] ) );
  EDFFX1 \registers_reg[802][0]  ( .D(n8013), .E(n324), .CK(clk), .Q(
        \registers[802][0] ) );
  EDFFX1 \registers_reg[798][7]  ( .D(n8400), .E(n848), .CK(clk), .Q(
        \registers[798][7] ) );
  EDFFX1 \registers_reg[798][6]  ( .D(n8342), .E(n848), .CK(clk), .Q(
        \registers[798][6] ) );
  EDFFX1 \registers_reg[798][5]  ( .D(n8284), .E(n848), .CK(clk), .Q(
        \registers[798][5] ) );
  EDFFX1 \registers_reg[798][4]  ( .D(n8226), .E(n848), .CK(clk), .Q(
        \registers[798][4] ) );
  EDFFX1 \registers_reg[798][3]  ( .D(n8176), .E(n848), .CK(clk), .Q(
        \registers[798][3] ) );
  EDFFX1 \registers_reg[798][2]  ( .D(n8131), .E(n848), .CK(clk), .Q(
        \registers[798][2] ) );
  EDFFX1 \registers_reg[798][1]  ( .D(n8075), .E(n848), .CK(clk), .Q(
        \registers[798][1] ) );
  EDFFX1 \registers_reg[798][0]  ( .D(n8014), .E(n848), .CK(clk), .Q(
        \registers[798][0] ) );
  EDFFX1 \registers_reg[794][7]  ( .D(n8398), .E(n844), .CK(clk), .Q(
        \registers[794][7] ) );
  EDFFX1 \registers_reg[794][6]  ( .D(n8340), .E(n844), .CK(clk), .Q(
        \registers[794][6] ) );
  EDFFX1 \registers_reg[794][5]  ( .D(n8282), .E(n844), .CK(clk), .Q(
        \registers[794][5] ) );
  EDFFX1 \registers_reg[794][4]  ( .D(n8224), .E(n844), .CK(clk), .Q(
        \registers[794][4] ) );
  EDFFX1 \registers_reg[794][3]  ( .D(n8177), .E(n844), .CK(clk), .Q(
        \registers[794][3] ) );
  EDFFX1 \registers_reg[794][2]  ( .D(n8129), .E(n844), .CK(clk), .Q(
        \registers[794][2] ) );
  EDFFX1 \registers_reg[794][1]  ( .D(n8073), .E(n844), .CK(clk), .Q(
        \registers[794][1] ) );
  EDFFX1 \registers_reg[794][0]  ( .D(n8015), .E(n844), .CK(clk), .Q(
        \registers[794][0] ) );
  EDFFX1 \registers_reg[790][7]  ( .D(n8399), .E(n840), .CK(clk), .Q(
        \registers[790][7] ) );
  EDFFX1 \registers_reg[790][6]  ( .D(n8341), .E(n840), .CK(clk), .Q(
        \registers[790][6] ) );
  EDFFX1 \registers_reg[790][5]  ( .D(n8283), .E(n840), .CK(clk), .Q(
        \registers[790][5] ) );
  EDFFX1 \registers_reg[790][4]  ( .D(n8225), .E(n840), .CK(clk), .Q(
        \registers[790][4] ) );
  EDFFX1 \registers_reg[790][3]  ( .D(n8178), .E(n840), .CK(clk), .Q(
        \registers[790][3] ) );
  EDFFX1 \registers_reg[790][2]  ( .D(n8130), .E(n840), .CK(clk), .Q(
        \registers[790][2] ) );
  EDFFX1 \registers_reg[790][1]  ( .D(n8074), .E(n840), .CK(clk), .Q(
        \registers[790][1] ) );
  EDFFX1 \registers_reg[790][0]  ( .D(n8013), .E(n840), .CK(clk), .Q(
        \registers[790][0] ) );
  EDFFX1 \registers_reg[786][7]  ( .D(n8400), .E(n153), .CK(clk), .Q(
        \registers[786][7] ) );
  EDFFX1 \registers_reg[786][6]  ( .D(n8342), .E(n153), .CK(clk), .Q(
        \registers[786][6] ) );
  EDFFX1 \registers_reg[786][5]  ( .D(n8284), .E(n153), .CK(clk), .Q(
        \registers[786][5] ) );
  EDFFX1 \registers_reg[786][4]  ( .D(n8226), .E(n153), .CK(clk), .Q(
        \registers[786][4] ) );
  EDFFX1 \registers_reg[786][3]  ( .D(n8176), .E(n153), .CK(clk), .Q(
        \registers[786][3] ) );
  EDFFX1 \registers_reg[786][2]  ( .D(n8131), .E(n153), .CK(clk), .Q(
        \registers[786][2] ) );
  EDFFX1 \registers_reg[786][1]  ( .D(n8075), .E(n153), .CK(clk), .Q(
        \registers[786][1] ) );
  EDFFX1 \registers_reg[786][0]  ( .D(n8014), .E(n153), .CK(clk), .Q(
        \registers[786][0] ) );
  EDFFX1 \registers_reg[782][7]  ( .D(n8398), .E(n149), .CK(clk), .Q(
        \registers[782][7] ) );
  EDFFX1 \registers_reg[782][6]  ( .D(n8340), .E(n149), .CK(clk), .Q(
        \registers[782][6] ) );
  EDFFX1 \registers_reg[782][5]  ( .D(n8282), .E(n149), .CK(clk), .Q(
        \registers[782][5] ) );
  EDFFX1 \registers_reg[782][4]  ( .D(n8224), .E(n149), .CK(clk), .Q(
        \registers[782][4] ) );
  EDFFX1 \registers_reg[782][3]  ( .D(n8177), .E(n149), .CK(clk), .Q(
        \registers[782][3] ) );
  EDFFX1 \registers_reg[782][2]  ( .D(n8126), .E(n149), .CK(clk), .Q(
        \registers[782][2] ) );
  EDFFX1 \registers_reg[782][1]  ( .D(n8070), .E(n149), .CK(clk), .Q(
        \registers[782][1] ) );
  EDFFX1 \registers_reg[782][0]  ( .D(n8015), .E(n149), .CK(clk), .Q(
        \registers[782][0] ) );
  EDFFX1 \registers_reg[778][7]  ( .D(n8399), .E(n145), .CK(clk), .Q(
        \registers[778][7] ) );
  EDFFX1 \registers_reg[778][6]  ( .D(n8341), .E(n145), .CK(clk), .Q(
        \registers[778][6] ) );
  EDFFX1 \registers_reg[778][5]  ( .D(n8283), .E(n145), .CK(clk), .Q(
        \registers[778][5] ) );
  EDFFX1 \registers_reg[778][4]  ( .D(n8225), .E(n145), .CK(clk), .Q(
        \registers[778][4] ) );
  EDFFX1 \registers_reg[778][3]  ( .D(n8178), .E(n145), .CK(clk), .Q(
        \registers[778][3] ) );
  EDFFX1 \registers_reg[778][2]  ( .D(n8127), .E(n145), .CK(clk), .Q(
        \registers[778][2] ) );
  EDFFX1 \registers_reg[778][1]  ( .D(n8071), .E(n145), .CK(clk), .Q(
        \registers[778][1] ) );
  EDFFX1 \registers_reg[778][0]  ( .D(n8010), .E(n145), .CK(clk), .Q(
        \registers[778][0] ) );
  EDFFX1 \registers_reg[774][7]  ( .D(n8395), .E(n321), .CK(clk), .Q(
        \registers[774][7] ) );
  EDFFX1 \registers_reg[774][6]  ( .D(n8337), .E(n321), .CK(clk), .Q(
        \registers[774][6] ) );
  EDFFX1 \registers_reg[774][5]  ( .D(n8279), .E(n321), .CK(clk), .Q(
        \registers[774][5] ) );
  EDFFX1 \registers_reg[774][4]  ( .D(n8221), .E(n321), .CK(clk), .Q(
        \registers[774][4] ) );
  EDFFX1 \registers_reg[774][3]  ( .D(n8176), .E(n321), .CK(clk), .Q(
        \registers[774][3] ) );
  EDFFX1 \registers_reg[774][2]  ( .D(n8128), .E(n321), .CK(clk), .Q(
        \registers[774][2] ) );
  EDFFX1 \registers_reg[774][1]  ( .D(n8072), .E(n321), .CK(clk), .Q(
        \registers[774][1] ) );
  EDFFX1 \registers_reg[774][0]  ( .D(n8011), .E(n321), .CK(clk), .Q(
        \registers[774][0] ) );
  EDFFX1 \registers_reg[770][7]  ( .D(n8396), .E(n317), .CK(clk), .Q(
        \registers[770][7] ) );
  EDFFX1 \registers_reg[770][6]  ( .D(n8338), .E(n317), .CK(clk), .Q(
        \registers[770][6] ) );
  EDFFX1 \registers_reg[770][5]  ( .D(n8280), .E(n317), .CK(clk), .Q(
        \registers[770][5] ) );
  EDFFX1 \registers_reg[770][4]  ( .D(n8222), .E(n317), .CK(clk), .Q(
        \registers[770][4] ) );
  EDFFX1 \registers_reg[770][3]  ( .D(n8177), .E(n317), .CK(clk), .Q(
        \registers[770][3] ) );
  EDFFX1 \registers_reg[770][2]  ( .D(n8126), .E(n317), .CK(clk), .Q(
        \registers[770][2] ) );
  EDFFX1 \registers_reg[770][1]  ( .D(n8070), .E(n317), .CK(clk), .Q(
        \registers[770][1] ) );
  EDFFX1 \registers_reg[770][0]  ( .D(n8012), .E(n317), .CK(clk), .Q(
        \registers[770][0] ) );
  EDFFX1 \registers_reg[766][7]  ( .D(n8382), .E(n836), .CK(clk), .Q(
        \registers[766][7] ) );
  EDFFX1 \registers_reg[766][6]  ( .D(n8324), .E(n836), .CK(clk), .Q(
        \registers[766][6] ) );
  EDFFX1 \registers_reg[766][5]  ( .D(n8266), .E(n836), .CK(clk), .Q(
        \registers[766][5] ) );
  EDFFX1 \registers_reg[766][4]  ( .D(n8208), .E(n836), .CK(clk), .Q(
        \registers[766][4] ) );
  EDFFX1 \registers_reg[766][3]  ( .D(n8166), .E(n836), .CK(clk), .Q(
        \registers[766][3] ) );
  EDFFX1 \registers_reg[766][2]  ( .D(n8112), .E(n836), .CK(clk), .Q(
        \registers[766][2] ) );
  EDFFX1 \registers_reg[766][1]  ( .D(n8056), .E(n836), .CK(clk), .Q(
        \registers[766][1] ) );
  EDFFX1 \registers_reg[766][0]  ( .D(n7996), .E(n836), .CK(clk), .Q(
        \registers[766][0] ) );
  EDFFX1 \registers_reg[762][7]  ( .D(n8383), .E(n832), .CK(clk), .Q(
        \registers[762][7] ) );
  EDFFX1 \registers_reg[762][6]  ( .D(n8325), .E(n832), .CK(clk), .Q(
        \registers[762][6] ) );
  EDFFX1 \registers_reg[762][5]  ( .D(n8267), .E(n832), .CK(clk), .Q(
        \registers[762][5] ) );
  EDFFX1 \registers_reg[762][4]  ( .D(n8209), .E(n832), .CK(clk), .Q(
        \registers[762][4] ) );
  EDFFX1 \registers_reg[762][3]  ( .D(n8164), .E(n832), .CK(clk), .Q(
        \registers[762][3] ) );
  EDFFX1 \registers_reg[762][2]  ( .D(n8113), .E(n832), .CK(clk), .Q(
        \registers[762][2] ) );
  EDFFX1 \registers_reg[762][1]  ( .D(n8057), .E(n832), .CK(clk), .Q(
        \registers[762][1] ) );
  EDFFX1 \registers_reg[762][0]  ( .D(n7997), .E(n832), .CK(clk), .Q(
        \registers[762][0] ) );
  EDFFX1 \registers_reg[758][7]  ( .D(n8381), .E(n828), .CK(clk), .Q(
        \registers[758][7] ) );
  EDFFX1 \registers_reg[758][6]  ( .D(n8323), .E(n828), .CK(clk), .Q(
        \registers[758][6] ) );
  EDFFX1 \registers_reg[758][5]  ( .D(n8265), .E(n828), .CK(clk), .Q(
        \registers[758][5] ) );
  EDFFX1 \registers_reg[758][4]  ( .D(n8207), .E(n828), .CK(clk), .Q(
        \registers[758][4] ) );
  EDFFX1 \registers_reg[758][3]  ( .D(n8165), .E(n828), .CK(clk), .Q(
        \registers[758][3] ) );
  EDFFX1 \registers_reg[758][2]  ( .D(n8111), .E(n828), .CK(clk), .Q(
        \registers[758][2] ) );
  EDFFX1 \registers_reg[758][1]  ( .D(n8055), .E(n828), .CK(clk), .Q(
        \registers[758][1] ) );
  EDFFX1 \registers_reg[758][0]  ( .D(n8670), .E(n828), .CK(clk), .Q(
        \registers[758][0] ) );
  EDFFX1 \registers_reg[754][7]  ( .D(n8382), .E(n141), .CK(clk), .Q(
        \registers[754][7] ) );
  EDFFX1 \registers_reg[754][6]  ( .D(n8324), .E(n141), .CK(clk), .Q(
        \registers[754][6] ) );
  EDFFX1 \registers_reg[754][5]  ( .D(n8266), .E(n141), .CK(clk), .Q(
        \registers[754][5] ) );
  EDFFX1 \registers_reg[754][4]  ( .D(n8208), .E(n141), .CK(clk), .Q(
        \registers[754][4] ) );
  EDFFX1 \registers_reg[754][3]  ( .D(n8166), .E(n141), .CK(clk), .Q(
        \registers[754][3] ) );
  EDFFX1 \registers_reg[754][2]  ( .D(n8112), .E(n141), .CK(clk), .Q(
        \registers[754][2] ) );
  EDFFX1 \registers_reg[754][1]  ( .D(n8056), .E(n141), .CK(clk), .Q(
        \registers[754][1] ) );
  EDFFX1 \registers_reg[754][0]  ( .D(n7996), .E(n141), .CK(clk), .Q(
        \registers[754][0] ) );
  EDFFX1 \registers_reg[750][7]  ( .D(n8383), .E(n137), .CK(clk), .Q(
        \registers[750][7] ) );
  EDFFX1 \registers_reg[750][6]  ( .D(n8325), .E(n137), .CK(clk), .Q(
        \registers[750][6] ) );
  EDFFX1 \registers_reg[750][5]  ( .D(n8267), .E(n137), .CK(clk), .Q(
        \registers[750][5] ) );
  EDFFX1 \registers_reg[750][4]  ( .D(n8209), .E(n137), .CK(clk), .Q(
        \registers[750][4] ) );
  EDFFX1 \registers_reg[750][3]  ( .D(n8188), .E(n137), .CK(clk), .Q(
        \registers[750][3] ) );
  EDFFX1 \registers_reg[750][2]  ( .D(n8113), .E(n137), .CK(clk), .Q(
        \registers[750][2] ) );
  EDFFX1 \registers_reg[750][1]  ( .D(n8057), .E(n137), .CK(clk), .Q(
        \registers[750][1] ) );
  EDFFX1 \registers_reg[750][0]  ( .D(n7997), .E(n137), .CK(clk), .Q(
        \registers[750][0] ) );
  EDFFX1 \registers_reg[746][7]  ( .D(n8381), .E(n133), .CK(clk), .Q(
        \registers[746][7] ) );
  EDFFX1 \registers_reg[746][6]  ( .D(n8323), .E(n133), .CK(clk), .Q(
        \registers[746][6] ) );
  EDFFX1 \registers_reg[746][5]  ( .D(n8265), .E(n133), .CK(clk), .Q(
        \registers[746][5] ) );
  EDFFX1 \registers_reg[746][4]  ( .D(n8207), .E(n133), .CK(clk), .Q(
        \registers[746][4] ) );
  EDFFX1 \registers_reg[746][3]  ( .D(n8162), .E(n133), .CK(clk), .Q(
        \registers[746][3] ) );
  EDFFX1 \registers_reg[746][2]  ( .D(n8111), .E(n133), .CK(clk), .Q(
        \registers[746][2] ) );
  EDFFX1 \registers_reg[746][1]  ( .D(n8055), .E(n133), .CK(clk), .Q(
        \registers[746][1] ) );
  EDFFX1 \registers_reg[746][0]  ( .D(n8673), .E(n133), .CK(clk), .Q(
        \registers[746][0] ) );
  EDFFX1 \registers_reg[742][7]  ( .D(n8382), .E(n314), .CK(clk), .Q(
        \registers[742][7] ) );
  EDFFX1 \registers_reg[742][6]  ( .D(n8324), .E(n314), .CK(clk), .Q(
        \registers[742][6] ) );
  EDFFX1 \registers_reg[742][5]  ( .D(n8266), .E(n314), .CK(clk), .Q(
        \registers[742][5] ) );
  EDFFX1 \registers_reg[742][4]  ( .D(n8208), .E(n314), .CK(clk), .Q(
        \registers[742][4] ) );
  EDFFX1 \registers_reg[742][3]  ( .D(n8163), .E(n314), .CK(clk), .Q(
        \registers[742][3] ) );
  EDFFX1 \registers_reg[742][2]  ( .D(n8112), .E(n314), .CK(clk), .Q(
        \registers[742][2] ) );
  EDFFX1 \registers_reg[742][1]  ( .D(n8056), .E(n314), .CK(clk), .Q(
        \registers[742][1] ) );
  EDFFX1 \registers_reg[742][0]  ( .D(n7996), .E(n314), .CK(clk), .Q(
        \registers[742][0] ) );
  EDFFX1 \registers_reg[738][7]  ( .D(n8383), .E(n310), .CK(clk), .Q(
        \registers[738][7] ) );
  EDFFX1 \registers_reg[738][6]  ( .D(n8325), .E(n310), .CK(clk), .Q(
        \registers[738][6] ) );
  EDFFX1 \registers_reg[738][5]  ( .D(n8267), .E(n310), .CK(clk), .Q(
        \registers[738][5] ) );
  EDFFX1 \registers_reg[738][4]  ( .D(n8209), .E(n310), .CK(clk), .Q(
        \registers[738][4] ) );
  EDFFX1 \registers_reg[738][3]  ( .D(n8189), .E(n310), .CK(clk), .Q(
        \registers[738][3] ) );
  EDFFX1 \registers_reg[738][2]  ( .D(n8113), .E(n310), .CK(clk), .Q(
        \registers[738][2] ) );
  EDFFX1 \registers_reg[738][1]  ( .D(n8057), .E(n310), .CK(clk), .Q(
        \registers[738][1] ) );
  EDFFX1 \registers_reg[738][0]  ( .D(n7997), .E(n310), .CK(clk), .Q(
        \registers[738][0] ) );
  EDFFX1 \registers_reg[734][7]  ( .D(n8381), .E(n824), .CK(clk), .Q(
        \registers[734][7] ) );
  EDFFX1 \registers_reg[734][6]  ( .D(n8323), .E(n824), .CK(clk), .Q(
        \registers[734][6] ) );
  EDFFX1 \registers_reg[734][5]  ( .D(n8265), .E(n824), .CK(clk), .Q(
        \registers[734][5] ) );
  EDFFX1 \registers_reg[734][4]  ( .D(n8207), .E(n824), .CK(clk), .Q(
        \registers[734][4] ) );
  EDFFX1 \registers_reg[734][3]  ( .D(n8162), .E(n824), .CK(clk), .Q(
        \registers[734][3] ) );
  EDFFX1 \registers_reg[734][2]  ( .D(n8111), .E(n824), .CK(clk), .Q(
        \registers[734][2] ) );
  EDFFX1 \registers_reg[734][1]  ( .D(n8055), .E(n824), .CK(clk), .Q(
        \registers[734][1] ) );
  EDFFX1 \registers_reg[734][0]  ( .D(n8672), .E(n824), .CK(clk), .Q(
        \registers[734][0] ) );
  EDFFX1 \registers_reg[730][7]  ( .D(n8382), .E(n820), .CK(clk), .Q(
        \registers[730][7] ) );
  EDFFX1 \registers_reg[730][6]  ( .D(n8324), .E(n820), .CK(clk), .Q(
        \registers[730][6] ) );
  EDFFX1 \registers_reg[730][5]  ( .D(n8266), .E(n820), .CK(clk), .Q(
        \registers[730][5] ) );
  EDFFX1 \registers_reg[730][4]  ( .D(n8208), .E(n820), .CK(clk), .Q(
        \registers[730][4] ) );
  EDFFX1 \registers_reg[730][3]  ( .D(n8163), .E(n820), .CK(clk), .Q(
        \registers[730][3] ) );
  EDFFX1 \registers_reg[730][2]  ( .D(n8109), .E(n820), .CK(clk), .Q(
        \registers[730][2] ) );
  EDFFX1 \registers_reg[730][1]  ( .D(n8053), .E(n820), .CK(clk), .Q(
        \registers[730][1] ) );
  EDFFX1 \registers_reg[730][0]  ( .D(n7995), .E(n820), .CK(clk), .Q(
        \registers[730][0] ) );
  EDFFX1 \registers_reg[726][7]  ( .D(n8378), .E(n816), .CK(clk), .Q(
        \registers[726][7] ) );
  EDFFX1 \registers_reg[726][6]  ( .D(n8320), .E(n816), .CK(clk), .Q(
        \registers[726][6] ) );
  EDFFX1 \registers_reg[726][5]  ( .D(n8262), .E(n816), .CK(clk), .Q(
        \registers[726][5] ) );
  EDFFX1 \registers_reg[726][4]  ( .D(n8204), .E(n816), .CK(clk), .Q(
        \registers[726][4] ) );
  EDFFX1 \registers_reg[726][3]  ( .D(n8190), .E(n816), .CK(clk), .Q(
        \registers[726][3] ) );
  EDFFX1 \registers_reg[726][2]  ( .D(n8110), .E(n816), .CK(clk), .Q(
        \registers[726][2] ) );
  EDFFX1 \registers_reg[726][1]  ( .D(n8054), .E(n816), .CK(clk), .Q(
        \registers[726][1] ) );
  EDFFX1 \registers_reg[726][0]  ( .D(n8026), .E(n816), .CK(clk), .Q(
        \registers[726][0] ) );
  EDFFX1 \registers_reg[722][7]  ( .D(n8379), .E(n129), .CK(clk), .Q(
        \registers[722][7] ) );
  EDFFX1 \registers_reg[722][6]  ( .D(n8321), .E(n129), .CK(clk), .Q(
        \registers[722][6] ) );
  EDFFX1 \registers_reg[722][5]  ( .D(n8263), .E(n129), .CK(clk), .Q(
        \registers[722][5] ) );
  EDFFX1 \registers_reg[722][4]  ( .D(n8205), .E(n129), .CK(clk), .Q(
        \registers[722][4] ) );
  EDFFX1 \registers_reg[722][3]  ( .D(n8162), .E(n129), .CK(clk), .Q(
        \registers[722][3] ) );
  EDFFX1 \registers_reg[722][2]  ( .D(n8108), .E(n129), .CK(clk), .Q(
        \registers[722][2] ) );
  EDFFX1 \registers_reg[722][1]  ( .D(n8052), .E(n129), .CK(clk), .Q(
        \registers[722][1] ) );
  EDFFX1 \registers_reg[722][0]  ( .D(n8034), .E(n129), .CK(clk), .Q(
        \registers[722][0] ) );
  EDFFX1 \registers_reg[718][7]  ( .D(n8380), .E(n125), .CK(clk), .Q(
        \registers[718][7] ) );
  EDFFX1 \registers_reg[718][6]  ( .D(n8322), .E(n125), .CK(clk), .Q(
        \registers[718][6] ) );
  EDFFX1 \registers_reg[718][5]  ( .D(n8264), .E(n125), .CK(clk), .Q(
        \registers[718][5] ) );
  EDFFX1 \registers_reg[718][4]  ( .D(n8206), .E(n125), .CK(clk), .Q(
        \registers[718][4] ) );
  EDFFX1 \registers_reg[718][3]  ( .D(n8163), .E(n125), .CK(clk), .Q(
        \registers[718][3] ) );
  EDFFX1 \registers_reg[718][2]  ( .D(n8109), .E(n125), .CK(clk), .Q(
        \registers[718][2] ) );
  EDFFX1 \registers_reg[718][1]  ( .D(n8053), .E(n125), .CK(clk), .Q(
        \registers[718][1] ) );
  EDFFX1 \registers_reg[718][0]  ( .D(n7995), .E(n125), .CK(clk), .Q(
        \registers[718][0] ) );
  EDFFX1 \registers_reg[714][7]  ( .D(n8378), .E(n121), .CK(clk), .Q(
        \registers[714][7] ) );
  EDFFX1 \registers_reg[714][6]  ( .D(n8320), .E(n121), .CK(clk), .Q(
        \registers[714][6] ) );
  EDFFX1 \registers_reg[714][5]  ( .D(n8262), .E(n121), .CK(clk), .Q(
        \registers[714][5] ) );
  EDFFX1 \registers_reg[714][4]  ( .D(n8204), .E(n121), .CK(clk), .Q(
        \registers[714][4] ) );
  EDFFX1 \registers_reg[714][3]  ( .D(n8185), .E(n121), .CK(clk), .Q(
        \registers[714][3] ) );
  EDFFX1 \registers_reg[714][2]  ( .D(n8110), .E(n121), .CK(clk), .Q(
        \registers[714][2] ) );
  EDFFX1 \registers_reg[714][1]  ( .D(n8054), .E(n121), .CK(clk), .Q(
        \registers[714][1] ) );
  EDFFX1 \registers_reg[714][0]  ( .D(n8022), .E(n121), .CK(clk), .Q(
        \registers[714][0] ) );
  EDFFX1 \registers_reg[710][7]  ( .D(n8379), .E(n307), .CK(clk), .Q(
        \registers[710][7] ) );
  EDFFX1 \registers_reg[710][6]  ( .D(n8321), .E(n307), .CK(clk), .Q(
        \registers[710][6] ) );
  EDFFX1 \registers_reg[710][5]  ( .D(n8263), .E(n307), .CK(clk), .Q(
        \registers[710][5] ) );
  EDFFX1 \registers_reg[710][4]  ( .D(n8205), .E(n307), .CK(clk), .Q(
        \registers[710][4] ) );
  EDFFX1 \registers_reg[710][3]  ( .D(n8162), .E(n307), .CK(clk), .Q(
        \registers[710][3] ) );
  EDFFX1 \registers_reg[710][2]  ( .D(n8108), .E(n307), .CK(clk), .Q(
        \registers[710][2] ) );
  EDFFX1 \registers_reg[710][1]  ( .D(n8052), .E(n307), .CK(clk), .Q(
        \registers[710][1] ) );
  EDFFX1 \registers_reg[710][0]  ( .D(n8035), .E(n307), .CK(clk), .Q(
        \registers[710][0] ) );
  EDFFX1 \registers_reg[706][7]  ( .D(n8380), .E(n303), .CK(clk), .Q(
        \registers[706][7] ) );
  EDFFX1 \registers_reg[706][6]  ( .D(n8322), .E(n303), .CK(clk), .Q(
        \registers[706][6] ) );
  EDFFX1 \registers_reg[706][5]  ( .D(n8264), .E(n303), .CK(clk), .Q(
        \registers[706][5] ) );
  EDFFX1 \registers_reg[706][4]  ( .D(n8206), .E(n303), .CK(clk), .Q(
        \registers[706][4] ) );
  EDFFX1 \registers_reg[706][3]  ( .D(n8163), .E(n303), .CK(clk), .Q(
        \registers[706][3] ) );
  EDFFX1 \registers_reg[706][2]  ( .D(n8109), .E(n303), .CK(clk), .Q(
        \registers[706][2] ) );
  EDFFX1 \registers_reg[706][1]  ( .D(n8053), .E(n303), .CK(clk), .Q(
        \registers[706][1] ) );
  EDFFX1 \registers_reg[706][0]  ( .D(n7995), .E(n303), .CK(clk), .Q(
        \registers[706][0] ) );
  EDFFX1 \registers_reg[702][7]  ( .D(n8379), .E(n812), .CK(clk), .Q(
        \registers[702][7] ) );
  EDFFX1 \registers_reg[702][6]  ( .D(n8321), .E(n812), .CK(clk), .Q(
        \registers[702][6] ) );
  EDFFX1 \registers_reg[702][5]  ( .D(n8263), .E(n812), .CK(clk), .Q(
        \registers[702][5] ) );
  EDFFX1 \registers_reg[702][4]  ( .D(n8205), .E(n812), .CK(clk), .Q(
        \registers[702][4] ) );
  EDFFX1 \registers_reg[702][3]  ( .D(n8162), .E(n812), .CK(clk), .Q(
        \registers[702][3] ) );
  EDFFX1 \registers_reg[702][2]  ( .D(n8108), .E(n812), .CK(clk), .Q(
        \registers[702][2] ) );
  EDFFX1 \registers_reg[702][1]  ( .D(n8052), .E(n812), .CK(clk), .Q(
        \registers[702][1] ) );
  EDFFX1 \registers_reg[702][0]  ( .D(n8036), .E(n812), .CK(clk), .Q(
        \registers[702][0] ) );
  EDFFX1 \registers_reg[698][7]  ( .D(n8380), .E(n808), .CK(clk), .Q(
        \registers[698][7] ) );
  EDFFX1 \registers_reg[698][6]  ( .D(n8322), .E(n808), .CK(clk), .Q(
        \registers[698][6] ) );
  EDFFX1 \registers_reg[698][5]  ( .D(n8264), .E(n808), .CK(clk), .Q(
        \registers[698][5] ) );
  EDFFX1 \registers_reg[698][4]  ( .D(n8206), .E(n808), .CK(clk), .Q(
        \registers[698][4] ) );
  EDFFX1 \registers_reg[698][3]  ( .D(n8163), .E(n808), .CK(clk), .Q(
        \registers[698][3] ) );
  EDFFX1 \registers_reg[698][2]  ( .D(n8109), .E(n808), .CK(clk), .Q(
        \registers[698][2] ) );
  EDFFX1 \registers_reg[698][1]  ( .D(n8053), .E(n808), .CK(clk), .Q(
        \registers[698][1] ) );
  EDFFX1 \registers_reg[698][0]  ( .D(n7995), .E(n808), .CK(clk), .Q(
        \registers[698][0] ) );
  EDFFX1 \registers_reg[694][7]  ( .D(n8378), .E(n804), .CK(clk), .Q(
        \registers[694][7] ) );
  EDFFX1 \registers_reg[694][6]  ( .D(n8320), .E(n804), .CK(clk), .Q(
        \registers[694][6] ) );
  EDFFX1 \registers_reg[694][5]  ( .D(n8262), .E(n804), .CK(clk), .Q(
        \registers[694][5] ) );
  EDFFX1 \registers_reg[694][4]  ( .D(n8204), .E(n804), .CK(clk), .Q(
        \registers[694][4] ) );
  EDFFX1 \registers_reg[694][3]  ( .D(n8186), .E(n804), .CK(clk), .Q(
        \registers[694][3] ) );
  EDFFX1 \registers_reg[694][2]  ( .D(n8110), .E(n804), .CK(clk), .Q(
        \registers[694][2] ) );
  EDFFX1 \registers_reg[694][1]  ( .D(n8054), .E(n804), .CK(clk), .Q(
        \registers[694][1] ) );
  EDFFX1 \registers_reg[694][0]  ( .D(n8023), .E(n804), .CK(clk), .Q(
        \registers[694][0] ) );
  EDFFX1 \registers_reg[690][7]  ( .D(n8379), .E(n117), .CK(clk), .Q(
        \registers[690][7] ) );
  EDFFX1 \registers_reg[690][6]  ( .D(n8321), .E(n117), .CK(clk), .Q(
        \registers[690][6] ) );
  EDFFX1 \registers_reg[690][5]  ( .D(n8263), .E(n117), .CK(clk), .Q(
        \registers[690][5] ) );
  EDFFX1 \registers_reg[690][4]  ( .D(n8205), .E(n117), .CK(clk), .Q(
        \registers[690][4] ) );
  EDFFX1 \registers_reg[690][3]  ( .D(n8161), .E(n117), .CK(clk), .Q(
        \registers[690][3] ) );
  EDFFX1 \registers_reg[690][2]  ( .D(n8108), .E(n117), .CK(clk), .Q(
        \registers[690][2] ) );
  EDFFX1 \registers_reg[690][1]  ( .D(n8052), .E(n117), .CK(clk), .Q(
        \registers[690][1] ) );
  EDFFX1 \registers_reg[690][0]  ( .D(n8046), .E(n117), .CK(clk), .Q(
        \registers[690][0] ) );
  EDFFX1 \registers_reg[686][7]  ( .D(n8380), .E(n113), .CK(clk), .Q(
        \registers[686][7] ) );
  EDFFX1 \registers_reg[686][6]  ( .D(n8322), .E(n113), .CK(clk), .Q(
        \registers[686][6] ) );
  EDFFX1 \registers_reg[686][5]  ( .D(n8264), .E(n113), .CK(clk), .Q(
        \registers[686][5] ) );
  EDFFX1 \registers_reg[686][4]  ( .D(n8206), .E(n113), .CK(clk), .Q(
        \registers[686][4] ) );
  EDFFX1 \registers_reg[686][3]  ( .D(n8161), .E(n113), .CK(clk), .Q(
        \registers[686][3] ) );
  EDFFX1 \registers_reg[686][2]  ( .D(n8109), .E(n113), .CK(clk), .Q(
        \registers[686][2] ) );
  EDFFX1 \registers_reg[686][1]  ( .D(n8053), .E(n113), .CK(clk), .Q(
        \registers[686][1] ) );
  EDFFX1 \registers_reg[686][0]  ( .D(n7995), .E(n113), .CK(clk), .Q(
        \registers[686][0] ) );
  EDFFX1 \registers_reg[682][7]  ( .D(n8378), .E(n109), .CK(clk), .Q(
        \registers[682][7] ) );
  EDFFX1 \registers_reg[682][6]  ( .D(n8320), .E(n109), .CK(clk), .Q(
        \registers[682][6] ) );
  EDFFX1 \registers_reg[682][5]  ( .D(n8262), .E(n109), .CK(clk), .Q(
        \registers[682][5] ) );
  EDFFX1 \registers_reg[682][4]  ( .D(n8204), .E(n109), .CK(clk), .Q(
        \registers[682][4] ) );
  EDFFX1 \registers_reg[682][3]  ( .D(n8161), .E(n109), .CK(clk), .Q(
        \registers[682][3] ) );
  EDFFX1 \registers_reg[682][2]  ( .D(n8110), .E(n109), .CK(clk), .Q(
        \registers[682][2] ) );
  EDFFX1 \registers_reg[682][1]  ( .D(n8054), .E(n109), .CK(clk), .Q(
        \registers[682][1] ) );
  EDFFX1 \registers_reg[682][0]  ( .D(n8024), .E(n109), .CK(clk), .Q(
        \registers[682][0] ) );
  EDFFX1 \registers_reg[678][7]  ( .D(n8377), .E(n300), .CK(clk), .Q(
        \registers[678][7] ) );
  EDFFX1 \registers_reg[678][6]  ( .D(n8319), .E(n300), .CK(clk), .Q(
        \registers[678][6] ) );
  EDFFX1 \registers_reg[678][5]  ( .D(n8261), .E(n300), .CK(clk), .Q(
        \registers[678][5] ) );
  EDFFX1 \registers_reg[678][4]  ( .D(n8203), .E(n300), .CK(clk), .Q(
        \registers[678][4] ) );
  EDFFX1 \registers_reg[678][3]  ( .D(n8161), .E(n300), .CK(clk), .Q(
        \registers[678][3] ) );
  EDFFX1 \registers_reg[678][2]  ( .D(n8105), .E(n300), .CK(clk), .Q(
        \registers[678][2] ) );
  EDFFX1 \registers_reg[678][1]  ( .D(n8049), .E(n300), .CK(clk), .Q(
        \registers[678][1] ) );
  EDFFX1 \registers_reg[678][0]  ( .D(n7994), .E(n300), .CK(clk), .Q(
        \registers[678][0] ) );
  EDFFX1 \registers_reg[674][7]  ( .D(n8377), .E(n296), .CK(clk), .Q(
        \registers[674][7] ) );
  EDFFX1 \registers_reg[674][6]  ( .D(n8319), .E(n296), .CK(clk), .Q(
        \registers[674][6] ) );
  EDFFX1 \registers_reg[674][5]  ( .D(n8261), .E(n296), .CK(clk), .Q(
        \registers[674][5] ) );
  EDFFX1 \registers_reg[674][4]  ( .D(n8203), .E(n296), .CK(clk), .Q(
        \registers[674][4] ) );
  EDFFX1 \registers_reg[674][3]  ( .D(n8184), .E(n296), .CK(clk), .Q(
        \registers[674][3] ) );
  EDFFX1 \registers_reg[674][2]  ( .D(n8106), .E(n296), .CK(clk), .Q(
        \registers[674][2] ) );
  EDFFX1 \registers_reg[674][1]  ( .D(n8050), .E(n296), .CK(clk), .Q(
        \registers[674][1] ) );
  EDFFX1 \registers_reg[674][0]  ( .D(n7994), .E(n296), .CK(clk), .Q(
        \registers[674][0] ) );
  EDFFX1 \registers_reg[670][7]  ( .D(n8377), .E(n800), .CK(clk), .Q(
        \registers[670][7] ) );
  EDFFX1 \registers_reg[670][6]  ( .D(n8319), .E(n800), .CK(clk), .Q(
        \registers[670][6] ) );
  EDFFX1 \registers_reg[670][5]  ( .D(n8261), .E(n800), .CK(clk), .Q(
        \registers[670][5] ) );
  EDFFX1 \registers_reg[670][4]  ( .D(n8203), .E(n800), .CK(clk), .Q(
        \registers[670][4] ) );
  EDFFX1 \registers_reg[670][3]  ( .D(n8182), .E(n800), .CK(clk), .Q(
        \registers[670][3] ) );
  EDFFX1 \registers_reg[670][2]  ( .D(n8107), .E(n800), .CK(clk), .Q(
        \registers[670][2] ) );
  EDFFX1 \registers_reg[670][1]  ( .D(n8051), .E(n800), .CK(clk), .Q(
        \registers[670][1] ) );
  EDFFX1 \registers_reg[670][0]  ( .D(n7994), .E(n800), .CK(clk), .Q(
        \registers[670][0] ) );
  EDFFX1 \registers_reg[666][7]  ( .D(n8398), .E(n796), .CK(clk), .Q(
        \registers[666][7] ) );
  EDFFX1 \registers_reg[666][6]  ( .D(n8340), .E(n796), .CK(clk), .Q(
        \registers[666][6] ) );
  EDFFX1 \registers_reg[666][5]  ( .D(n8282), .E(n796), .CK(clk), .Q(
        \registers[666][5] ) );
  EDFFX1 \registers_reg[666][4]  ( .D(n8224), .E(n796), .CK(clk), .Q(
        \registers[666][4] ) );
  EDFFX1 \registers_reg[666][3]  ( .D(n8183), .E(n796), .CK(clk), .Q(
        \registers[666][3] ) );
  EDFFX1 \registers_reg[666][2]  ( .D(n8105), .E(n796), .CK(clk), .Q(
        \registers[666][2] ) );
  EDFFX1 \registers_reg[666][1]  ( .D(n8049), .E(n796), .CK(clk), .Q(
        \registers[666][1] ) );
  EDFFX1 \registers_reg[666][0]  ( .D(n8688), .E(n796), .CK(clk), .Q(
        \registers[666][0] ) );
  EDFFX1 \registers_reg[662][7]  ( .D(n8399), .E(n792), .CK(clk), .Q(
        \registers[662][7] ) );
  EDFFX1 \registers_reg[662][6]  ( .D(n8341), .E(n792), .CK(clk), .Q(
        \registers[662][6] ) );
  EDFFX1 \registers_reg[662][5]  ( .D(n8283), .E(n792), .CK(clk), .Q(
        \registers[662][5] ) );
  EDFFX1 \registers_reg[662][4]  ( .D(n8225), .E(n792), .CK(clk), .Q(
        \registers[662][4] ) );
  EDFFX1 \registers_reg[662][3]  ( .D(n8184), .E(n792), .CK(clk), .Q(
        \registers[662][3] ) );
  EDFFX1 \registers_reg[662][2]  ( .D(n8106), .E(n792), .CK(clk), .Q(
        \registers[662][2] ) );
  EDFFX1 \registers_reg[662][1]  ( .D(n8050), .E(n792), .CK(clk), .Q(
        \registers[662][1] ) );
  EDFFX1 \registers_reg[662][0]  ( .D(n8033), .E(n792), .CK(clk), .Q(
        \registers[662][0] ) );
  EDFFX1 \registers_reg[658][7]  ( .D(n8392), .E(n105), .CK(clk), .Q(
        \registers[658][7] ) );
  EDFFX1 \registers_reg[658][6]  ( .D(n8334), .E(n105), .CK(clk), .Q(
        \registers[658][6] ) );
  EDFFX1 \registers_reg[658][5]  ( .D(n8276), .E(n105), .CK(clk), .Q(
        \registers[658][5] ) );
  EDFFX1 \registers_reg[658][4]  ( .D(n8218), .E(n105), .CK(clk), .Q(
        \registers[658][4] ) );
  EDFFX1 \registers_reg[658][3]  ( .D(n8182), .E(n105), .CK(clk), .Q(
        \registers[658][3] ) );
  EDFFX1 \registers_reg[658][2]  ( .D(n8107), .E(n105), .CK(clk), .Q(
        \registers[658][2] ) );
  EDFFX1 \registers_reg[658][1]  ( .D(n8051), .E(n105), .CK(clk), .Q(
        \registers[658][1] ) );
  EDFFX1 \registers_reg[658][0]  ( .D(data_in[0]), .E(n105), .CK(clk), .Q(
        \registers[658][0] ) );
  EDFFX1 \registers_reg[654][7]  ( .D(n8393), .E(n101), .CK(clk), .Q(
        \registers[654][7] ) );
  EDFFX1 \registers_reg[654][6]  ( .D(n8335), .E(n101), .CK(clk), .Q(
        \registers[654][6] ) );
  EDFFX1 \registers_reg[654][5]  ( .D(n8277), .E(n101), .CK(clk), .Q(
        \registers[654][5] ) );
  EDFFX1 \registers_reg[654][4]  ( .D(n8219), .E(n101), .CK(clk), .Q(
        \registers[654][4] ) );
  EDFFX1 \registers_reg[654][3]  ( .D(n8183), .E(n101), .CK(clk), .Q(
        \registers[654][3] ) );
  EDFFX1 \registers_reg[654][2]  ( .D(n8105), .E(n101), .CK(clk), .Q(
        \registers[654][2] ) );
  EDFFX1 \registers_reg[654][1]  ( .D(n8049), .E(n101), .CK(clk), .Q(
        \registers[654][1] ) );
  EDFFX1 \registers_reg[654][0]  ( .D(n8663), .E(n101), .CK(clk), .Q(
        \registers[654][0] ) );
  EDFFX1 \registers_reg[650][7]  ( .D(n8389), .E(n97), .CK(clk), .Q(
        \registers[650][7] ) );
  EDFFX1 \registers_reg[650][6]  ( .D(n8331), .E(n97), .CK(clk), .Q(
        \registers[650][6] ) );
  EDFFX1 \registers_reg[650][5]  ( .D(n8273), .E(n97), .CK(clk), .Q(
        \registers[650][5] ) );
  EDFFX1 \registers_reg[650][4]  ( .D(n8215), .E(n97), .CK(clk), .Q(
        \registers[650][4] ) );
  EDFFX1 \registers_reg[650][3]  ( .D(n8753), .E(n97), .CK(clk), .Q(
        \registers[650][3] ) );
  EDFFX1 \registers_reg[650][2]  ( .D(n8106), .E(n97), .CK(clk), .Q(
        \registers[650][2] ) );
  EDFFX1 \registers_reg[650][1]  ( .D(n8050), .E(n97), .CK(clk), .Q(
        \registers[650][1] ) );
  EDFFX1 \registers_reg[650][0]  ( .D(n8001), .E(n97), .CK(clk), .Q(
        \registers[650][0] ) );
  EDFFX1 \registers_reg[646][7]  ( .D(n8390), .E(n293), .CK(clk), .Q(
        \registers[646][7] ) );
  EDFFX1 \registers_reg[646][6]  ( .D(n8332), .E(n293), .CK(clk), .Q(
        \registers[646][6] ) );
  EDFFX1 \registers_reg[646][5]  ( .D(n8274), .E(n293), .CK(clk), .Q(
        \registers[646][5] ) );
  EDFFX1 \registers_reg[646][4]  ( .D(n8216), .E(n293), .CK(clk), .Q(
        \registers[646][4] ) );
  EDFFX1 \registers_reg[646][3]  ( .D(n8170), .E(n293), .CK(clk), .Q(
        \registers[646][3] ) );
  EDFFX1 \registers_reg[646][2]  ( .D(n8107), .E(n293), .CK(clk), .Q(
        \registers[646][2] ) );
  EDFFX1 \registers_reg[646][1]  ( .D(n8051), .E(n293), .CK(clk), .Q(
        \registers[646][1] ) );
  EDFFX1 \registers_reg[646][0]  ( .D(n8002), .E(n293), .CK(clk), .Q(
        \registers[646][0] ) );
  EDFFX1 \registers_reg[642][7]  ( .D(n8386), .E(n289), .CK(clk), .Q(
        \registers[642][7] ) );
  EDFFX1 \registers_reg[642][6]  ( .D(n8328), .E(n289), .CK(clk), .Q(
        \registers[642][6] ) );
  EDFFX1 \registers_reg[642][5]  ( .D(n8270), .E(n289), .CK(clk), .Q(
        \registers[642][5] ) );
  EDFFX1 \registers_reg[642][4]  ( .D(n8212), .E(n289), .CK(clk), .Q(
        \registers[642][4] ) );
  EDFFX1 \registers_reg[642][3]  ( .D(n8171), .E(n289), .CK(clk), .Q(
        \registers[642][3] ) );
  EDFFX1 \registers_reg[642][2]  ( .D(n8105), .E(n289), .CK(clk), .Q(
        \registers[642][2] ) );
  EDFFX1 \registers_reg[642][1]  ( .D(n8049), .E(n289), .CK(clk), .Q(
        \registers[642][1] ) );
  EDFFX1 \registers_reg[642][0]  ( .D(n8003), .E(n289), .CK(clk), .Q(
        \registers[642][0] ) );
  EDFFX1 \registers_reg[638][7]  ( .D(n8390), .E(n788), .CK(clk), .Q(
        \registers[638][7] ) );
  EDFFX1 \registers_reg[638][6]  ( .D(n8332), .E(n788), .CK(clk), .Q(
        \registers[638][6] ) );
  EDFFX1 \registers_reg[638][5]  ( .D(n8274), .E(n788), .CK(clk), .Q(
        \registers[638][5] ) );
  EDFFX1 \registers_reg[638][4]  ( .D(n8216), .E(n788), .CK(clk), .Q(
        \registers[638][4] ) );
  EDFFX1 \registers_reg[638][3]  ( .D(n8172), .E(n788), .CK(clk), .Q(
        \registers[638][3] ) );
  EDFFX1 \registers_reg[638][2]  ( .D(n8121), .E(n788), .CK(clk), .Q(
        \registers[638][2] ) );
  EDFFX1 \registers_reg[638][1]  ( .D(n8065), .E(n788), .CK(clk), .Q(
        \registers[638][1] ) );
  EDFFX1 \registers_reg[638][0]  ( .D(n8006), .E(n788), .CK(clk), .Q(
        \registers[638][0] ) );
  EDFFX1 \registers_reg[634][7]  ( .D(n8391), .E(n784), .CK(clk), .Q(
        \registers[634][7] ) );
  EDFFX1 \registers_reg[634][6]  ( .D(n8333), .E(n784), .CK(clk), .Q(
        \registers[634][6] ) );
  EDFFX1 \registers_reg[634][5]  ( .D(n8275), .E(n784), .CK(clk), .Q(
        \registers[634][5] ) );
  EDFFX1 \registers_reg[634][4]  ( .D(n8217), .E(n784), .CK(clk), .Q(
        \registers[634][4] ) );
  EDFFX1 \registers_reg[634][3]  ( .D(n8170), .E(n784), .CK(clk), .Q(
        \registers[634][3] ) );
  EDFFX1 \registers_reg[634][2]  ( .D(n8122), .E(n784), .CK(clk), .Q(
        \registers[634][2] ) );
  EDFFX1 \registers_reg[634][1]  ( .D(n8066), .E(n784), .CK(clk), .Q(
        \registers[634][1] ) );
  EDFFX1 \registers_reg[634][0]  ( .D(n8004), .E(n784), .CK(clk), .Q(
        \registers[634][0] ) );
  EDFFX1 \registers_reg[630][7]  ( .D(n8389), .E(n780), .CK(clk), .Q(
        \registers[630][7] ) );
  EDFFX1 \registers_reg[630][6]  ( .D(n8331), .E(n780), .CK(clk), .Q(
        \registers[630][6] ) );
  EDFFX1 \registers_reg[630][5]  ( .D(n8273), .E(n780), .CK(clk), .Q(
        \registers[630][5] ) );
  EDFFX1 \registers_reg[630][4]  ( .D(n8215), .E(n780), .CK(clk), .Q(
        \registers[630][4] ) );
  EDFFX1 \registers_reg[630][3]  ( .D(n8171), .E(n780), .CK(clk), .Q(
        \registers[630][3] ) );
  EDFFX1 \registers_reg[630][2]  ( .D(n8117), .E(n780), .CK(clk), .Q(
        \registers[630][2] ) );
  EDFFX1 \registers_reg[630][1]  ( .D(n8061), .E(n780), .CK(clk), .Q(
        \registers[630][1] ) );
  EDFFX1 \registers_reg[630][0]  ( .D(n8005), .E(n780), .CK(clk), .Q(
        \registers[630][0] ) );
  EDFFX1 \registers_reg[626][7]  ( .D(n8390), .E(n93), .CK(clk), .Q(
        \registers[626][7] ) );
  EDFFX1 \registers_reg[626][6]  ( .D(n8332), .E(n93), .CK(clk), .Q(
        \registers[626][6] ) );
  EDFFX1 \registers_reg[626][5]  ( .D(n8274), .E(n93), .CK(clk), .Q(
        \registers[626][5] ) );
  EDFFX1 \registers_reg[626][4]  ( .D(n8216), .E(n93), .CK(clk), .Q(
        \registers[626][4] ) );
  EDFFX1 \registers_reg[626][3]  ( .D(n8172), .E(n93), .CK(clk), .Q(
        \registers[626][3] ) );
  EDFFX1 \registers_reg[626][2]  ( .D(n8118), .E(n93), .CK(clk), .Q(
        \registers[626][2] ) );
  EDFFX1 \registers_reg[626][1]  ( .D(n8062), .E(n93), .CK(clk), .Q(
        \registers[626][1] ) );
  EDFFX1 \registers_reg[626][0]  ( .D(n8003), .E(n93), .CK(clk), .Q(
        \registers[626][0] ) );
  EDFFX1 \registers_reg[622][7]  ( .D(n8386), .E(n89), .CK(clk), .Q(
        \registers[622][7] ) );
  EDFFX1 \registers_reg[622][6]  ( .D(n8328), .E(n89), .CK(clk), .Q(
        \registers[622][6] ) );
  EDFFX1 \registers_reg[622][5]  ( .D(n8270), .E(n89), .CK(clk), .Q(
        \registers[622][5] ) );
  EDFFX1 \registers_reg[622][4]  ( .D(n8212), .E(n89), .CK(clk), .Q(
        \registers[622][4] ) );
  EDFFX1 \registers_reg[622][3]  ( .D(n8167), .E(n89), .CK(clk), .Q(
        \registers[622][3] ) );
  EDFFX1 \registers_reg[622][2]  ( .D(n8119), .E(n89), .CK(clk), .Q(
        \registers[622][2] ) );
  EDFFX1 \registers_reg[622][1]  ( .D(n8063), .E(n89), .CK(clk), .Q(
        \registers[622][1] ) );
  EDFFX1 \registers_reg[622][0]  ( .D(n8001), .E(n89), .CK(clk), .Q(
        \registers[622][0] ) );
  EDFFX1 \registers_reg[618][7]  ( .D(n8387), .E(n85), .CK(clk), .Q(
        \registers[618][7] ) );
  EDFFX1 \registers_reg[618][6]  ( .D(n8329), .E(n85), .CK(clk), .Q(
        \registers[618][6] ) );
  EDFFX1 \registers_reg[618][5]  ( .D(n8271), .E(n85), .CK(clk), .Q(
        \registers[618][5] ) );
  EDFFX1 \registers_reg[618][4]  ( .D(n8213), .E(n85), .CK(clk), .Q(
        \registers[618][4] ) );
  EDFFX1 \registers_reg[618][3]  ( .D(n8168), .E(n85), .CK(clk), .Q(
        \registers[618][3] ) );
  EDFFX1 \registers_reg[618][2]  ( .D(n8117), .E(n85), .CK(clk), .Q(
        \registers[618][2] ) );
  EDFFX1 \registers_reg[618][1]  ( .D(n8061), .E(n85), .CK(clk), .Q(
        \registers[618][1] ) );
  EDFFX1 \registers_reg[618][0]  ( .D(n8002), .E(n85), .CK(clk), .Q(
        \registers[618][0] ) );
  EDFFX1 \registers_reg[614][7]  ( .D(n8388), .E(n286), .CK(clk), .Q(
        \registers[614][7] ) );
  EDFFX1 \registers_reg[614][6]  ( .D(n8330), .E(n286), .CK(clk), .Q(
        \registers[614][6] ) );
  EDFFX1 \registers_reg[614][5]  ( .D(n8272), .E(n286), .CK(clk), .Q(
        \registers[614][5] ) );
  EDFFX1 \registers_reg[614][4]  ( .D(n8214), .E(n286), .CK(clk), .Q(
        \registers[614][4] ) );
  EDFFX1 \registers_reg[614][3]  ( .D(n8169), .E(n286), .CK(clk), .Q(
        \registers[614][3] ) );
  EDFFX1 \registers_reg[614][2]  ( .D(n8118), .E(n286), .CK(clk), .Q(
        \registers[614][2] ) );
  EDFFX1 \registers_reg[614][1]  ( .D(n8062), .E(n286), .CK(clk), .Q(
        \registers[614][1] ) );
  EDFFX1 \registers_reg[614][0]  ( .D(n8003), .E(n286), .CK(clk), .Q(
        \registers[614][0] ) );
  EDFFX1 \registers_reg[610][7]  ( .D(n8386), .E(n282), .CK(clk), .Q(
        \registers[610][7] ) );
  EDFFX1 \registers_reg[610][6]  ( .D(n8328), .E(n282), .CK(clk), .Q(
        \registers[610][6] ) );
  EDFFX1 \registers_reg[610][5]  ( .D(n8270), .E(n282), .CK(clk), .Q(
        \registers[610][5] ) );
  EDFFX1 \registers_reg[610][4]  ( .D(n8212), .E(n282), .CK(clk), .Q(
        \registers[610][4] ) );
  EDFFX1 \registers_reg[610][3]  ( .D(n8167), .E(n282), .CK(clk), .Q(
        \registers[610][3] ) );
  EDFFX1 \registers_reg[610][2]  ( .D(n8119), .E(n282), .CK(clk), .Q(
        \registers[610][2] ) );
  EDFFX1 \registers_reg[610][1]  ( .D(n8063), .E(n282), .CK(clk), .Q(
        \registers[610][1] ) );
  EDFFX1 \registers_reg[610][0]  ( .D(n8001), .E(n282), .CK(clk), .Q(
        \registers[610][0] ) );
  EDFFX1 \registers_reg[606][7]  ( .D(n8387), .E(n776), .CK(clk), .Q(
        \registers[606][7] ) );
  EDFFX1 \registers_reg[606][6]  ( .D(n8329), .E(n776), .CK(clk), .Q(
        \registers[606][6] ) );
  EDFFX1 \registers_reg[606][5]  ( .D(n8271), .E(n776), .CK(clk), .Q(
        \registers[606][5] ) );
  EDFFX1 \registers_reg[606][4]  ( .D(n8213), .E(n776), .CK(clk), .Q(
        \registers[606][4] ) );
  EDFFX1 \registers_reg[606][3]  ( .D(n8168), .E(n776), .CK(clk), .Q(
        \registers[606][3] ) );
  EDFFX1 \registers_reg[606][2]  ( .D(n8117), .E(n776), .CK(clk), .Q(
        \registers[606][2] ) );
  EDFFX1 \registers_reg[606][1]  ( .D(n8061), .E(n776), .CK(clk), .Q(
        \registers[606][1] ) );
  EDFFX1 \registers_reg[606][0]  ( .D(n8002), .E(n776), .CK(clk), .Q(
        \registers[606][0] ) );
  EDFFX1 \registers_reg[602][7]  ( .D(n8388), .E(n772), .CK(clk), .Q(
        \registers[602][7] ) );
  EDFFX1 \registers_reg[602][6]  ( .D(n8330), .E(n772), .CK(clk), .Q(
        \registers[602][6] ) );
  EDFFX1 \registers_reg[602][5]  ( .D(n8272), .E(n772), .CK(clk), .Q(
        \registers[602][5] ) );
  EDFFX1 \registers_reg[602][4]  ( .D(n8214), .E(n772), .CK(clk), .Q(
        \registers[602][4] ) );
  EDFFX1 \registers_reg[602][3]  ( .D(n8169), .E(n772), .CK(clk), .Q(
        \registers[602][3] ) );
  EDFFX1 \registers_reg[602][2]  ( .D(n8118), .E(n772), .CK(clk), .Q(
        \registers[602][2] ) );
  EDFFX1 \registers_reg[602][1]  ( .D(n8062), .E(n772), .CK(clk), .Q(
        \registers[602][1] ) );
  EDFFX1 \registers_reg[602][0]  ( .D(n8003), .E(n772), .CK(clk), .Q(
        \registers[602][0] ) );
  EDFFX1 \registers_reg[598][7]  ( .D(n8386), .E(n768), .CK(clk), .Q(
        \registers[598][7] ) );
  EDFFX1 \registers_reg[598][6]  ( .D(n8328), .E(n768), .CK(clk), .Q(
        \registers[598][6] ) );
  EDFFX1 \registers_reg[598][5]  ( .D(n8270), .E(n768), .CK(clk), .Q(
        \registers[598][5] ) );
  EDFFX1 \registers_reg[598][4]  ( .D(n8212), .E(n768), .CK(clk), .Q(
        \registers[598][4] ) );
  EDFFX1 \registers_reg[598][3]  ( .D(n8167), .E(n768), .CK(clk), .Q(
        \registers[598][3] ) );
  EDFFX1 \registers_reg[598][2]  ( .D(n8119), .E(n768), .CK(clk), .Q(
        \registers[598][2] ) );
  EDFFX1 \registers_reg[598][1]  ( .D(n8063), .E(n768), .CK(clk), .Q(
        \registers[598][1] ) );
  EDFFX1 \registers_reg[598][0]  ( .D(n8001), .E(n768), .CK(clk), .Q(
        \registers[598][0] ) );
  EDFFX1 \registers_reg[594][7]  ( .D(n8387), .E(n81), .CK(clk), .Q(
        \registers[594][7] ) );
  EDFFX1 \registers_reg[594][6]  ( .D(n8329), .E(n81), .CK(clk), .Q(
        \registers[594][6] ) );
  EDFFX1 \registers_reg[594][5]  ( .D(n8271), .E(n81), .CK(clk), .Q(
        \registers[594][5] ) );
  EDFFX1 \registers_reg[594][4]  ( .D(n8213), .E(n81), .CK(clk), .Q(
        \registers[594][4] ) );
  EDFFX1 \registers_reg[594][3]  ( .D(n8168), .E(n81), .CK(clk), .Q(
        \registers[594][3] ) );
  EDFFX1 \registers_reg[594][2]  ( .D(n8117), .E(n81), .CK(clk), .Q(
        \registers[594][2] ) );
  EDFFX1 \registers_reg[594][1]  ( .D(n8061), .E(n81), .CK(clk), .Q(
        \registers[594][1] ) );
  EDFFX1 \registers_reg[594][0]  ( .D(n8002), .E(n81), .CK(clk), .Q(
        \registers[594][0] ) );
  EDFFX1 \registers_reg[590][7]  ( .D(n8388), .E(n77), .CK(clk), .Q(
        \registers[590][7] ) );
  EDFFX1 \registers_reg[590][6]  ( .D(n8330), .E(n77), .CK(clk), .Q(
        \registers[590][6] ) );
  EDFFX1 \registers_reg[590][5]  ( .D(n8272), .E(n77), .CK(clk), .Q(
        \registers[590][5] ) );
  EDFFX1 \registers_reg[590][4]  ( .D(n8214), .E(n77), .CK(clk), .Q(
        \registers[590][4] ) );
  EDFFX1 \registers_reg[590][3]  ( .D(n8169), .E(n77), .CK(clk), .Q(
        \registers[590][3] ) );
  EDFFX1 \registers_reg[590][2]  ( .D(n8118), .E(n77), .CK(clk), .Q(
        \registers[590][2] ) );
  EDFFX1 \registers_reg[590][1]  ( .D(n8062), .E(n77), .CK(clk), .Q(
        \registers[590][1] ) );
  EDFFX1 \registers_reg[590][0]  ( .D(n8003), .E(n77), .CK(clk), .Q(
        \registers[590][0] ) );
  EDFFX1 \registers_reg[586][7]  ( .D(n8386), .E(n73), .CK(clk), .Q(
        \registers[586][7] ) );
  EDFFX1 \registers_reg[586][6]  ( .D(n8328), .E(n73), .CK(clk), .Q(
        \registers[586][6] ) );
  EDFFX1 \registers_reg[586][5]  ( .D(n8270), .E(n73), .CK(clk), .Q(
        \registers[586][5] ) );
  EDFFX1 \registers_reg[586][4]  ( .D(n8212), .E(n73), .CK(clk), .Q(
        \registers[586][4] ) );
  EDFFX1 \registers_reg[586][3]  ( .D(n8167), .E(n73), .CK(clk), .Q(
        \registers[586][3] ) );
  EDFFX1 \registers_reg[586][2]  ( .D(n8119), .E(n73), .CK(clk), .Q(
        \registers[586][2] ) );
  EDFFX1 \registers_reg[586][1]  ( .D(n8063), .E(n73), .CK(clk), .Q(
        \registers[586][1] ) );
  EDFFX1 \registers_reg[586][0]  ( .D(n8001), .E(n73), .CK(clk), .Q(
        \registers[586][0] ) );
  EDFFX1 \registers_reg[582][7]  ( .D(n8387), .E(n279), .CK(clk), .Q(
        \registers[582][7] ) );
  EDFFX1 \registers_reg[582][6]  ( .D(n8329), .E(n279), .CK(clk), .Q(
        \registers[582][6] ) );
  EDFFX1 \registers_reg[582][5]  ( .D(n8271), .E(n279), .CK(clk), .Q(
        \registers[582][5] ) );
  EDFFX1 \registers_reg[582][4]  ( .D(n8213), .E(n279), .CK(clk), .Q(
        \registers[582][4] ) );
  EDFFX1 \registers_reg[582][3]  ( .D(n8168), .E(n279), .CK(clk), .Q(
        \registers[582][3] ) );
  EDFFX1 \registers_reg[582][2]  ( .D(n8117), .E(n279), .CK(clk), .Q(
        \registers[582][2] ) );
  EDFFX1 \registers_reg[582][1]  ( .D(n8061), .E(n279), .CK(clk), .Q(
        \registers[582][1] ) );
  EDFFX1 \registers_reg[582][0]  ( .D(n8002), .E(n279), .CK(clk), .Q(
        \registers[582][0] ) );
  EDFFX1 \registers_reg[578][7]  ( .D(n8388), .E(n275), .CK(clk), .Q(
        \registers[578][7] ) );
  EDFFX1 \registers_reg[578][6]  ( .D(n8330), .E(n275), .CK(clk), .Q(
        \registers[578][6] ) );
  EDFFX1 \registers_reg[578][5]  ( .D(n8272), .E(n275), .CK(clk), .Q(
        \registers[578][5] ) );
  EDFFX1 \registers_reg[578][4]  ( .D(n8214), .E(n275), .CK(clk), .Q(
        \registers[578][4] ) );
  EDFFX1 \registers_reg[578][3]  ( .D(n8169), .E(n275), .CK(clk), .Q(
        \registers[578][3] ) );
  EDFFX1 \registers_reg[578][2]  ( .D(n8115), .E(n275), .CK(clk), .Q(
        \registers[578][2] ) );
  EDFFX1 \registers_reg[578][1]  ( .D(n8059), .E(n275), .CK(clk), .Q(
        \registers[578][1] ) );
  EDFFX1 \registers_reg[578][0]  ( .D(n8003), .E(n275), .CK(clk), .Q(
        \registers[578][0] ) );
  EDFFX1 \registers_reg[574][7]  ( .D(n8385), .E(n764), .CK(clk), .Q(
        \registers[574][7] ) );
  EDFFX1 \registers_reg[574][6]  ( .D(n8327), .E(n764), .CK(clk), .Q(
        \registers[574][6] ) );
  EDFFX1 \registers_reg[574][5]  ( .D(n8269), .E(n764), .CK(clk), .Q(
        \registers[574][5] ) );
  EDFFX1 \registers_reg[574][4]  ( .D(n8211), .E(n764), .CK(clk), .Q(
        \registers[574][4] ) );
  EDFFX1 \registers_reg[574][3]  ( .D(n8168), .E(n764), .CK(clk), .Q(
        \registers[574][3] ) );
  EDFFX1 \registers_reg[574][2]  ( .D(n8114), .E(n764), .CK(clk), .Q(
        \registers[574][2] ) );
  EDFFX1 \registers_reg[574][1]  ( .D(n8058), .E(n764), .CK(clk), .Q(
        \registers[574][1] ) );
  EDFFX1 \registers_reg[574][0]  ( .D(n7999), .E(n764), .CK(clk), .Q(
        \registers[574][0] ) );
  EDFFX1 \registers_reg[570][7]  ( .D(n8384), .E(n760), .CK(clk), .Q(
        \registers[570][7] ) );
  EDFFX1 \registers_reg[570][6]  ( .D(n8326), .E(n760), .CK(clk), .Q(
        \registers[570][6] ) );
  EDFFX1 \registers_reg[570][5]  ( .D(n8268), .E(n760), .CK(clk), .Q(
        \registers[570][5] ) );
  EDFFX1 \registers_reg[570][4]  ( .D(n8210), .E(n760), .CK(clk), .Q(
        \registers[570][4] ) );
  EDFFX1 \registers_reg[570][3]  ( .D(n8169), .E(n760), .CK(clk), .Q(
        \registers[570][3] ) );
  EDFFX1 \registers_reg[570][2]  ( .D(n8115), .E(n760), .CK(clk), .Q(
        \registers[570][2] ) );
  EDFFX1 \registers_reg[570][1]  ( .D(n8059), .E(n760), .CK(clk), .Q(
        \registers[570][1] ) );
  EDFFX1 \registers_reg[570][0]  ( .D(n8000), .E(n760), .CK(clk), .Q(
        \registers[570][0] ) );
  EDFFX1 \registers_reg[566][7]  ( .D(n8404), .E(n756), .CK(clk), .Q(
        \registers[566][7] ) );
  EDFFX1 \registers_reg[566][6]  ( .D(n8346), .E(n756), .CK(clk), .Q(
        \registers[566][6] ) );
  EDFFX1 \registers_reg[566][5]  ( .D(n8288), .E(n756), .CK(clk), .Q(
        \registers[566][5] ) );
  EDFFX1 \registers_reg[566][4]  ( .D(n8230), .E(n756), .CK(clk), .Q(
        \registers[566][4] ) );
  EDFFX1 \registers_reg[566][3]  ( .D(n8167), .E(n756), .CK(clk), .Q(
        \registers[566][3] ) );
  EDFFX1 \registers_reg[566][2]  ( .D(n8116), .E(n756), .CK(clk), .Q(
        \registers[566][2] ) );
  EDFFX1 \registers_reg[566][1]  ( .D(n8060), .E(n756), .CK(clk), .Q(
        \registers[566][1] ) );
  EDFFX1 \registers_reg[566][0]  ( .D(n7998), .E(n756), .CK(clk), .Q(
        \registers[566][0] ) );
  EDFFX1 \registers_reg[562][7]  ( .D(n8385), .E(n69), .CK(clk), .Q(
        \registers[562][7] ) );
  EDFFX1 \registers_reg[562][6]  ( .D(n8327), .E(n69), .CK(clk), .Q(
        \registers[562][6] ) );
  EDFFX1 \registers_reg[562][5]  ( .D(n8269), .E(n69), .CK(clk), .Q(
        \registers[562][5] ) );
  EDFFX1 \registers_reg[562][4]  ( .D(n8211), .E(n69), .CK(clk), .Q(
        \registers[562][4] ) );
  EDFFX1 \registers_reg[562][3]  ( .D(n8165), .E(n69), .CK(clk), .Q(
        \registers[562][3] ) );
  EDFFX1 \registers_reg[562][2]  ( .D(n8114), .E(n69), .CK(clk), .Q(
        \registers[562][2] ) );
  EDFFX1 \registers_reg[562][1]  ( .D(n8058), .E(n69), .CK(clk), .Q(
        \registers[562][1] ) );
  EDFFX1 \registers_reg[562][0]  ( .D(n7999), .E(n69), .CK(clk), .Q(
        \registers[562][0] ) );
  EDFFX1 \registers_reg[558][7]  ( .D(n8384), .E(n65), .CK(clk), .Q(
        \registers[558][7] ) );
  EDFFX1 \registers_reg[558][6]  ( .D(n8326), .E(n65), .CK(clk), .Q(
        \registers[558][6] ) );
  EDFFX1 \registers_reg[558][5]  ( .D(n8268), .E(n65), .CK(clk), .Q(
        \registers[558][5] ) );
  EDFFX1 \registers_reg[558][4]  ( .D(n8210), .E(n65), .CK(clk), .Q(
        \registers[558][4] ) );
  EDFFX1 \registers_reg[558][3]  ( .D(n8166), .E(n65), .CK(clk), .Q(
        \registers[558][3] ) );
  EDFFX1 \registers_reg[558][2]  ( .D(n8115), .E(n65), .CK(clk), .Q(
        \registers[558][2] ) );
  EDFFX1 \registers_reg[558][1]  ( .D(n8059), .E(n65), .CK(clk), .Q(
        \registers[558][1] ) );
  EDFFX1 \registers_reg[558][0]  ( .D(n8000), .E(n65), .CK(clk), .Q(
        \registers[558][0] ) );
  EDFFX1 \registers_reg[554][7]  ( .D(n8424), .E(n61), .CK(clk), .Q(
        \registers[554][7] ) );
  EDFFX1 \registers_reg[554][6]  ( .D(n8366), .E(n61), .CK(clk), .Q(
        \registers[554][6] ) );
  EDFFX1 \registers_reg[554][5]  ( .D(n8308), .E(n61), .CK(clk), .Q(
        \registers[554][5] ) );
  EDFFX1 \registers_reg[554][4]  ( .D(n8250), .E(n61), .CK(clk), .Q(
        \registers[554][4] ) );
  EDFFX1 \registers_reg[554][3]  ( .D(n8164), .E(n61), .CK(clk), .Q(
        \registers[554][3] ) );
  EDFFX1 \registers_reg[554][2]  ( .D(n8116), .E(n61), .CK(clk), .Q(
        \registers[554][2] ) );
  EDFFX1 \registers_reg[554][1]  ( .D(n8060), .E(n61), .CK(clk), .Q(
        \registers[554][1] ) );
  EDFFX1 \registers_reg[554][0]  ( .D(n7998), .E(n61), .CK(clk), .Q(
        \registers[554][0] ) );
  EDFFX1 \registers_reg[550][7]  ( .D(n8385), .E(n272), .CK(clk), .Q(
        \registers[550][7] ) );
  EDFFX1 \registers_reg[550][6]  ( .D(n8327), .E(n272), .CK(clk), .Q(
        \registers[550][6] ) );
  EDFFX1 \registers_reg[550][5]  ( .D(n8269), .E(n272), .CK(clk), .Q(
        \registers[550][5] ) );
  EDFFX1 \registers_reg[550][4]  ( .D(n8211), .E(n272), .CK(clk), .Q(
        \registers[550][4] ) );
  EDFFX1 \registers_reg[550][3]  ( .D(n8165), .E(n272), .CK(clk), .Q(
        \registers[550][3] ) );
  EDFFX1 \registers_reg[550][2]  ( .D(n8114), .E(n272), .CK(clk), .Q(
        \registers[550][2] ) );
  EDFFX1 \registers_reg[550][1]  ( .D(n8058), .E(n272), .CK(clk), .Q(
        \registers[550][1] ) );
  EDFFX1 \registers_reg[550][0]  ( .D(n7999), .E(n272), .CK(clk), .Q(
        \registers[550][0] ) );
  EDFFX1 \registers_reg[546][7]  ( .D(n8384), .E(n268), .CK(clk), .Q(
        \registers[546][7] ) );
  EDFFX1 \registers_reg[546][6]  ( .D(n8326), .E(n268), .CK(clk), .Q(
        \registers[546][6] ) );
  EDFFX1 \registers_reg[546][5]  ( .D(n8268), .E(n268), .CK(clk), .Q(
        \registers[546][5] ) );
  EDFFX1 \registers_reg[546][4]  ( .D(n8210), .E(n268), .CK(clk), .Q(
        \registers[546][4] ) );
  EDFFX1 \registers_reg[546][3]  ( .D(n8166), .E(n268), .CK(clk), .Q(
        \registers[546][3] ) );
  EDFFX1 \registers_reg[546][2]  ( .D(n8115), .E(n268), .CK(clk), .Q(
        \registers[546][2] ) );
  EDFFX1 \registers_reg[546][1]  ( .D(n8059), .E(n268), .CK(clk), .Q(
        \registers[546][1] ) );
  EDFFX1 \registers_reg[546][0]  ( .D(n8000), .E(n268), .CK(clk), .Q(
        \registers[546][0] ) );
  EDFFX1 \registers_reg[542][7]  ( .D(n8421), .E(n752), .CK(clk), .Q(
        \registers[542][7] ) );
  EDFFX1 \registers_reg[542][6]  ( .D(n8363), .E(n752), .CK(clk), .Q(
        \registers[542][6] ) );
  EDFFX1 \registers_reg[542][5]  ( .D(n8305), .E(n752), .CK(clk), .Q(
        \registers[542][5] ) );
  EDFFX1 \registers_reg[542][4]  ( .D(n8247), .E(n752), .CK(clk), .Q(
        \registers[542][4] ) );
  EDFFX1 \registers_reg[542][3]  ( .D(n8164), .E(n752), .CK(clk), .Q(
        \registers[542][3] ) );
  EDFFX1 \registers_reg[542][2]  ( .D(n8116), .E(n752), .CK(clk), .Q(
        \registers[542][2] ) );
  EDFFX1 \registers_reg[542][1]  ( .D(n8060), .E(n752), .CK(clk), .Q(
        \registers[542][1] ) );
  EDFFX1 \registers_reg[542][0]  ( .D(n7998), .E(n752), .CK(clk), .Q(
        \registers[542][0] ) );
  EDFFX1 \registers_reg[538][7]  ( .D(n8385), .E(n748), .CK(clk), .Q(
        \registers[538][7] ) );
  EDFFX1 \registers_reg[538][6]  ( .D(n8327), .E(n748), .CK(clk), .Q(
        \registers[538][6] ) );
  EDFFX1 \registers_reg[538][5]  ( .D(n8269), .E(n748), .CK(clk), .Q(
        \registers[538][5] ) );
  EDFFX1 \registers_reg[538][4]  ( .D(n8211), .E(n748), .CK(clk), .Q(
        \registers[538][4] ) );
  EDFFX1 \registers_reg[538][3]  ( .D(n8165), .E(n748), .CK(clk), .Q(
        \registers[538][3] ) );
  EDFFX1 \registers_reg[538][2]  ( .D(n8114), .E(n748), .CK(clk), .Q(
        \registers[538][2] ) );
  EDFFX1 \registers_reg[538][1]  ( .D(n8058), .E(n748), .CK(clk), .Q(
        \registers[538][1] ) );
  EDFFX1 \registers_reg[538][0]  ( .D(n7999), .E(n748), .CK(clk), .Q(
        \registers[538][0] ) );
  EDFFX1 \registers_reg[534][7]  ( .D(n8384), .E(n744), .CK(clk), .Q(
        \registers[534][7] ) );
  EDFFX1 \registers_reg[534][6]  ( .D(n8326), .E(n744), .CK(clk), .Q(
        \registers[534][6] ) );
  EDFFX1 \registers_reg[534][5]  ( .D(n8268), .E(n744), .CK(clk), .Q(
        \registers[534][5] ) );
  EDFFX1 \registers_reg[534][4]  ( .D(n8210), .E(n744), .CK(clk), .Q(
        \registers[534][4] ) );
  EDFFX1 \registers_reg[534][3]  ( .D(n8166), .E(n744), .CK(clk), .Q(
        \registers[534][3] ) );
  EDFFX1 \registers_reg[534][2]  ( .D(n8115), .E(n744), .CK(clk), .Q(
        \registers[534][2] ) );
  EDFFX1 \registers_reg[534][1]  ( .D(n8059), .E(n744), .CK(clk), .Q(
        \registers[534][1] ) );
  EDFFX1 \registers_reg[534][0]  ( .D(n8000), .E(n744), .CK(clk), .Q(
        \registers[534][0] ) );
  EDFFX1 \registers_reg[530][7]  ( .D(n8424), .E(n57), .CK(clk), .Q(
        \registers[530][7] ) );
  EDFFX1 \registers_reg[530][6]  ( .D(n8366), .E(n57), .CK(clk), .Q(
        \registers[530][6] ) );
  EDFFX1 \registers_reg[530][5]  ( .D(n8308), .E(n57), .CK(clk), .Q(
        \registers[530][5] ) );
  EDFFX1 \registers_reg[530][4]  ( .D(n8250), .E(n57), .CK(clk), .Q(
        \registers[530][4] ) );
  EDFFX1 \registers_reg[530][3]  ( .D(n8164), .E(n57), .CK(clk), .Q(
        \registers[530][3] ) );
  EDFFX1 \registers_reg[530][2]  ( .D(n8116), .E(n57), .CK(clk), .Q(
        \registers[530][2] ) );
  EDFFX1 \registers_reg[530][1]  ( .D(n8060), .E(n57), .CK(clk), .Q(
        \registers[530][1] ) );
  EDFFX1 \registers_reg[530][0]  ( .D(n7998), .E(n57), .CK(clk), .Q(
        \registers[530][0] ) );
  EDFFX1 \registers_reg[526][7]  ( .D(n8381), .E(n52), .CK(clk), .Q(
        \registers[526][7] ) );
  EDFFX1 \registers_reg[526][6]  ( .D(n8323), .E(n52), .CK(clk), .Q(
        \registers[526][6] ) );
  EDFFX1 \registers_reg[526][5]  ( .D(n8265), .E(n52), .CK(clk), .Q(
        \registers[526][5] ) );
  EDFFX1 \registers_reg[526][4]  ( .D(n8207), .E(n52), .CK(clk), .Q(
        \registers[526][4] ) );
  EDFFX1 \registers_reg[526][3]  ( .D(n8165), .E(n52), .CK(clk), .Q(
        \registers[526][3] ) );
  EDFFX1 \registers_reg[526][2]  ( .D(n8111), .E(n52), .CK(clk), .Q(
        \registers[526][2] ) );
  EDFFX1 \registers_reg[526][1]  ( .D(n8055), .E(n52), .CK(clk), .Q(
        \registers[526][1] ) );
  EDFFX1 \registers_reg[526][0]  ( .D(n7997), .E(n52), .CK(clk), .Q(
        \registers[526][0] ) );
  EDFFX1 \registers_reg[522][7]  ( .D(n8382), .E(n48), .CK(clk), .Q(
        \registers[522][7] ) );
  EDFFX1 \registers_reg[522][6]  ( .D(n8324), .E(n48), .CK(clk), .Q(
        \registers[522][6] ) );
  EDFFX1 \registers_reg[522][5]  ( .D(n8266), .E(n48), .CK(clk), .Q(
        \registers[522][5] ) );
  EDFFX1 \registers_reg[522][4]  ( .D(n8208), .E(n48), .CK(clk), .Q(
        \registers[522][4] ) );
  EDFFX1 \registers_reg[522][3]  ( .D(n8166), .E(n48), .CK(clk), .Q(
        \registers[522][3] ) );
  EDFFX1 \registers_reg[522][2]  ( .D(n8112), .E(n48), .CK(clk), .Q(
        \registers[522][2] ) );
  EDFFX1 \registers_reg[522][1]  ( .D(n8056), .E(n48), .CK(clk), .Q(
        \registers[522][1] ) );
  EDFFX1 \registers_reg[522][0]  ( .D(n8675), .E(n48), .CK(clk), .Q(
        \registers[522][0] ) );
  EDFFX1 \registers_reg[518][7]  ( .D(n8383), .E(n265), .CK(clk), .Q(
        \registers[518][7] ) );
  EDFFX1 \registers_reg[518][6]  ( .D(n8325), .E(n265), .CK(clk), .Q(
        \registers[518][6] ) );
  EDFFX1 \registers_reg[518][5]  ( .D(n8267), .E(n265), .CK(clk), .Q(
        \registers[518][5] ) );
  EDFFX1 \registers_reg[518][4]  ( .D(n8209), .E(n265), .CK(clk), .Q(
        \registers[518][4] ) );
  EDFFX1 \registers_reg[518][3]  ( .D(n8164), .E(n265), .CK(clk), .Q(
        \registers[518][3] ) );
  EDFFX1 \registers_reg[518][2]  ( .D(n8113), .E(n265), .CK(clk), .Q(
        \registers[518][2] ) );
  EDFFX1 \registers_reg[518][1]  ( .D(n8057), .E(n265), .CK(clk), .Q(
        \registers[518][1] ) );
  EDFFX1 \registers_reg[518][0]  ( .D(n7996), .E(n265), .CK(clk), .Q(
        \registers[518][0] ) );
  EDFFX1 \registers_reg[514][7]  ( .D(n8381), .E(n261), .CK(clk), .Q(
        \registers[514][7] ) );
  EDFFX1 \registers_reg[514][6]  ( .D(n8323), .E(n261), .CK(clk), .Q(
        \registers[514][6] ) );
  EDFFX1 \registers_reg[514][5]  ( .D(n8265), .E(n261), .CK(clk), .Q(
        \registers[514][5] ) );
  EDFFX1 \registers_reg[514][4]  ( .D(n8207), .E(n261), .CK(clk), .Q(
        \registers[514][4] ) );
  EDFFX1 \registers_reg[514][3]  ( .D(n8165), .E(n261), .CK(clk), .Q(
        \registers[514][3] ) );
  EDFFX1 \registers_reg[514][2]  ( .D(n8111), .E(n261), .CK(clk), .Q(
        \registers[514][2] ) );
  EDFFX1 \registers_reg[514][1]  ( .D(n8055), .E(n261), .CK(clk), .Q(
        \registers[514][1] ) );
  EDFFX1 \registers_reg[514][0]  ( .D(n7997), .E(n261), .CK(clk), .Q(
        \registers[514][0] ) );
  EDFFX1 \registers_reg[510][7]  ( .D(n8429), .E(n740), .CK(clk), .Q(
        \registers[510][7] ) );
  EDFFX1 \registers_reg[510][6]  ( .D(n8371), .E(n740), .CK(clk), .Q(
        \registers[510][6] ) );
  EDFFX1 \registers_reg[510][5]  ( .D(n8313), .E(n740), .CK(clk), .Q(
        \registers[510][5] ) );
  EDFFX1 \registers_reg[510][4]  ( .D(n8255), .E(n740), .CK(clk), .Q(
        \registers[510][4] ) );
  EDFFX1 \registers_reg[510][3]  ( .D(n8200), .E(n740), .CK(clk), .Q(
        \registers[510][3] ) );
  EDFFX1 \registers_reg[510][2]  ( .D(n8157), .E(n740), .CK(clk), .Q(
        \registers[510][2] ) );
  EDFFX1 \registers_reg[510][1]  ( .D(n8101), .E(n740), .CK(clk), .Q(
        \registers[510][1] ) );
  EDFFX1 \registers_reg[510][0]  ( .D(n8041), .E(n740), .CK(clk), .Q(
        \registers[510][0] ) );
  EDFFX1 \registers_reg[506][7]  ( .D(n8425), .E(n736), .CK(clk), .Q(
        \registers[506][7] ) );
  EDFFX1 \registers_reg[506][6]  ( .D(n8367), .E(n736), .CK(clk), .Q(
        \registers[506][6] ) );
  EDFFX1 \registers_reg[506][5]  ( .D(n8309), .E(n736), .CK(clk), .Q(
        \registers[506][5] ) );
  EDFFX1 \registers_reg[506][4]  ( .D(n8251), .E(n736), .CK(clk), .Q(
        \registers[506][4] ) );
  EDFFX1 \registers_reg[506][3]  ( .D(n8201), .E(n736), .CK(clk), .Q(
        \registers[506][3] ) );
  EDFFX1 \registers_reg[506][2]  ( .D(n8155), .E(n736), .CK(clk), .Q(
        \registers[506][2] ) );
  EDFFX1 \registers_reg[506][1]  ( .D(n8099), .E(n736), .CK(clk), .Q(
        \registers[506][1] ) );
  EDFFX1 \registers_reg[506][0]  ( .D(n8042), .E(n736), .CK(clk), .Q(
        \registers[506][0] ) );
  EDFFX1 \registers_reg[502][7]  ( .D(n8426), .E(n732), .CK(clk), .Q(
        \registers[502][7] ) );
  EDFFX1 \registers_reg[502][6]  ( .D(n8368), .E(n732), .CK(clk), .Q(
        \registers[502][6] ) );
  EDFFX1 \registers_reg[502][5]  ( .D(n8310), .E(n732), .CK(clk), .Q(
        \registers[502][5] ) );
  EDFFX1 \registers_reg[502][4]  ( .D(n8252), .E(n732), .CK(clk), .Q(
        \registers[502][4] ) );
  EDFFX1 \registers_reg[502][3]  ( .D(n8202), .E(n732), .CK(clk), .Q(
        \registers[502][3] ) );
  EDFFX1 \registers_reg[502][2]  ( .D(n8156), .E(n732), .CK(clk), .Q(
        \registers[502][2] ) );
  EDFFX1 \registers_reg[502][1]  ( .D(n8100), .E(n732), .CK(clk), .Q(
        \registers[502][1] ) );
  EDFFX1 \registers_reg[502][0]  ( .D(n8040), .E(n732), .CK(clk), .Q(
        \registers[502][0] ) );
  EDFFX1 \registers_reg[498][7]  ( .D(n8427), .E(n44), .CK(clk), .Q(
        \registers[498][7] ) );
  EDFFX1 \registers_reg[498][6]  ( .D(n8369), .E(n44), .CK(clk), .Q(
        \registers[498][6] ) );
  EDFFX1 \registers_reg[498][5]  ( .D(n8311), .E(n44), .CK(clk), .Q(
        \registers[498][5] ) );
  EDFFX1 \registers_reg[498][4]  ( .D(n8253), .E(n44), .CK(clk), .Q(
        \registers[498][4] ) );
  EDFFX1 \registers_reg[498][3]  ( .D(n8200), .E(n44), .CK(clk), .Q(
        \registers[498][3] ) );
  EDFFX1 \registers_reg[498][2]  ( .D(n8157), .E(n44), .CK(clk), .Q(
        \registers[498][2] ) );
  EDFFX1 \registers_reg[498][1]  ( .D(n8101), .E(n44), .CK(clk), .Q(
        \registers[498][1] ) );
  EDFFX1 \registers_reg[498][0]  ( .D(n8041), .E(n44), .CK(clk), .Q(
        \registers[498][0] ) );
  EDFFX1 \registers_reg[494][7]  ( .D(n8425), .E(n40), .CK(clk), .Q(
        \registers[494][7] ) );
  EDFFX1 \registers_reg[494][6]  ( .D(n8367), .E(n40), .CK(clk), .Q(
        \registers[494][6] ) );
  EDFFX1 \registers_reg[494][5]  ( .D(n8309), .E(n40), .CK(clk), .Q(
        \registers[494][5] ) );
  EDFFX1 \registers_reg[494][4]  ( .D(n8251), .E(n40), .CK(clk), .Q(
        \registers[494][4] ) );
  EDFFX1 \registers_reg[494][3]  ( .D(n8201), .E(n40), .CK(clk), .Q(
        \registers[494][3] ) );
  EDFFX1 \registers_reg[494][2]  ( .D(n8155), .E(n40), .CK(clk), .Q(
        \registers[494][2] ) );
  EDFFX1 \registers_reg[494][1]  ( .D(n8099), .E(n40), .CK(clk), .Q(
        \registers[494][1] ) );
  EDFFX1 \registers_reg[494][0]  ( .D(n8042), .E(n40), .CK(clk), .Q(
        \registers[494][0] ) );
  EDFFX1 \registers_reg[490][7]  ( .D(n8426), .E(n36), .CK(clk), .Q(
        \registers[490][7] ) );
  EDFFX1 \registers_reg[490][6]  ( .D(n8368), .E(n36), .CK(clk), .Q(
        \registers[490][6] ) );
  EDFFX1 \registers_reg[490][5]  ( .D(n8310), .E(n36), .CK(clk), .Q(
        \registers[490][5] ) );
  EDFFX1 \registers_reg[490][4]  ( .D(n8252), .E(n36), .CK(clk), .Q(
        \registers[490][4] ) );
  EDFFX1 \registers_reg[490][3]  ( .D(n8202), .E(n36), .CK(clk), .Q(
        \registers[490][3] ) );
  EDFFX1 \registers_reg[490][2]  ( .D(n8156), .E(n36), .CK(clk), .Q(
        \registers[490][2] ) );
  EDFFX1 \registers_reg[490][1]  ( .D(n8100), .E(n36), .CK(clk), .Q(
        \registers[490][1] ) );
  EDFFX1 \registers_reg[490][0]  ( .D(n8040), .E(n36), .CK(clk), .Q(
        \registers[490][0] ) );
  EDFFX1 \registers_reg[486][7]  ( .D(n8427), .E(n258), .CK(clk), .Q(
        \registers[486][7] ) );
  EDFFX1 \registers_reg[486][6]  ( .D(n8369), .E(n258), .CK(clk), .Q(
        \registers[486][6] ) );
  EDFFX1 \registers_reg[486][5]  ( .D(n8311), .E(n258), .CK(clk), .Q(
        \registers[486][5] ) );
  EDFFX1 \registers_reg[486][4]  ( .D(n8253), .E(n258), .CK(clk), .Q(
        \registers[486][4] ) );
  EDFFX1 \registers_reg[486][3]  ( .D(n8197), .E(n258), .CK(clk), .Q(
        \registers[486][3] ) );
  EDFFX1 \registers_reg[486][2]  ( .D(n8157), .E(n258), .CK(clk), .Q(
        \registers[486][2] ) );
  EDFFX1 \registers_reg[486][1]  ( .D(n8101), .E(n258), .CK(clk), .Q(
        \registers[486][1] ) );
  EDFFX1 \registers_reg[486][0]  ( .D(n8041), .E(n258), .CK(clk), .Q(
        \registers[486][0] ) );
  EDFFX1 \registers_reg[482][7]  ( .D(n8425), .E(n254), .CK(clk), .Q(
        \registers[482][7] ) );
  EDFFX1 \registers_reg[482][6]  ( .D(n8367), .E(n254), .CK(clk), .Q(
        \registers[482][6] ) );
  EDFFX1 \registers_reg[482][5]  ( .D(n8309), .E(n254), .CK(clk), .Q(
        \registers[482][5] ) );
  EDFFX1 \registers_reg[482][4]  ( .D(n8251), .E(n254), .CK(clk), .Q(
        \registers[482][4] ) );
  EDFFX1 \registers_reg[482][3]  ( .D(n8198), .E(n254), .CK(clk), .Q(
        \registers[482][3] ) );
  EDFFX1 \registers_reg[482][2]  ( .D(n8155), .E(n254), .CK(clk), .Q(
        \registers[482][2] ) );
  EDFFX1 \registers_reg[482][1]  ( .D(n8099), .E(n254), .CK(clk), .Q(
        \registers[482][1] ) );
  EDFFX1 \registers_reg[482][0]  ( .D(n8042), .E(n254), .CK(clk), .Q(
        \registers[482][0] ) );
  EDFFX1 \registers_reg[478][7]  ( .D(n8426), .E(n728), .CK(clk), .Q(
        \registers[478][7] ) );
  EDFFX1 \registers_reg[478][6]  ( .D(n8368), .E(n728), .CK(clk), .Q(
        \registers[478][6] ) );
  EDFFX1 \registers_reg[478][5]  ( .D(n8310), .E(n728), .CK(clk), .Q(
        \registers[478][5] ) );
  EDFFX1 \registers_reg[478][4]  ( .D(n8252), .E(n728), .CK(clk), .Q(
        \registers[478][4] ) );
  EDFFX1 \registers_reg[478][3]  ( .D(n8199), .E(n728), .CK(clk), .Q(
        \registers[478][3] ) );
  EDFFX1 \registers_reg[478][2]  ( .D(n8156), .E(n728), .CK(clk), .Q(
        \registers[478][2] ) );
  EDFFX1 \registers_reg[478][1]  ( .D(n8100), .E(n728), .CK(clk), .Q(
        \registers[478][1] ) );
  EDFFX1 \registers_reg[478][0]  ( .D(n8040), .E(n728), .CK(clk), .Q(
        \registers[478][0] ) );
  EDFFX1 \registers_reg[474][7]  ( .D(n8427), .E(n724), .CK(clk), .Q(
        \registers[474][7] ) );
  EDFFX1 \registers_reg[474][6]  ( .D(n8369), .E(n724), .CK(clk), .Q(
        \registers[474][6] ) );
  EDFFX1 \registers_reg[474][5]  ( .D(n8311), .E(n724), .CK(clk), .Q(
        \registers[474][5] ) );
  EDFFX1 \registers_reg[474][4]  ( .D(n8253), .E(n724), .CK(clk), .Q(
        \registers[474][4] ) );
  EDFFX1 \registers_reg[474][3]  ( .D(n8197), .E(n724), .CK(clk), .Q(
        \registers[474][3] ) );
  EDFFX1 \registers_reg[474][2]  ( .D(n8157), .E(n724), .CK(clk), .Q(
        \registers[474][2] ) );
  EDFFX1 \registers_reg[474][1]  ( .D(n8101), .E(n724), .CK(clk), .Q(
        \registers[474][1] ) );
  EDFFX1 \registers_reg[474][0]  ( .D(n8041), .E(n724), .CK(clk), .Q(
        \registers[474][0] ) );
  EDFFX1 \registers_reg[470][7]  ( .D(n8425), .E(n720), .CK(clk), .Q(
        \registers[470][7] ) );
  EDFFX1 \registers_reg[470][6]  ( .D(n8367), .E(n720), .CK(clk), .Q(
        \registers[470][6] ) );
  EDFFX1 \registers_reg[470][5]  ( .D(n8309), .E(n720), .CK(clk), .Q(
        \registers[470][5] ) );
  EDFFX1 \registers_reg[470][4]  ( .D(n8251), .E(n720), .CK(clk), .Q(
        \registers[470][4] ) );
  EDFFX1 \registers_reg[470][3]  ( .D(n8198), .E(n720), .CK(clk), .Q(
        \registers[470][3] ) );
  EDFFX1 \registers_reg[470][2]  ( .D(n8152), .E(n720), .CK(clk), .Q(
        \registers[470][2] ) );
  EDFFX1 \registers_reg[470][1]  ( .D(n8096), .E(n720), .CK(clk), .Q(
        \registers[470][1] ) );
  EDFFX1 \registers_reg[470][0]  ( .D(n8039), .E(n720), .CK(clk), .Q(
        \registers[470][0] ) );
  EDFFX1 \registers_reg[466][7]  ( .D(n8426), .E(n32), .CK(clk), .Q(
        \registers[466][7] ) );
  EDFFX1 \registers_reg[466][6]  ( .D(n8368), .E(n32), .CK(clk), .Q(
        \registers[466][6] ) );
  EDFFX1 \registers_reg[466][5]  ( .D(n8310), .E(n32), .CK(clk), .Q(
        \registers[466][5] ) );
  EDFFX1 \registers_reg[466][4]  ( .D(n8252), .E(n32), .CK(clk), .Q(
        \registers[466][4] ) );
  EDFFX1 \registers_reg[466][3]  ( .D(n8199), .E(n32), .CK(clk), .Q(
        \registers[466][3] ) );
  EDFFX1 \registers_reg[466][2]  ( .D(n8153), .E(n32), .CK(clk), .Q(
        \registers[466][2] ) );
  EDFFX1 \registers_reg[466][1]  ( .D(n8097), .E(n32), .CK(clk), .Q(
        \registers[466][1] ) );
  EDFFX1 \registers_reg[466][0]  ( .D(n8037), .E(n32), .CK(clk), .Q(
        \registers[466][0] ) );
  EDFFX1 \registers_reg[462][7]  ( .D(n8427), .E(n28), .CK(clk), .Q(
        \registers[462][7] ) );
  EDFFX1 \registers_reg[462][6]  ( .D(n8369), .E(n28), .CK(clk), .Q(
        \registers[462][6] ) );
  EDFFX1 \registers_reg[462][5]  ( .D(n8311), .E(n28), .CK(clk), .Q(
        \registers[462][5] ) );
  EDFFX1 \registers_reg[462][4]  ( .D(n8253), .E(n28), .CK(clk), .Q(
        \registers[462][4] ) );
  EDFFX1 \registers_reg[462][3]  ( .D(n8197), .E(n28), .CK(clk), .Q(
        \registers[462][3] ) );
  EDFFX1 \registers_reg[462][2]  ( .D(n8154), .E(n28), .CK(clk), .Q(
        \registers[462][2] ) );
  EDFFX1 \registers_reg[462][1]  ( .D(n8098), .E(n28), .CK(clk), .Q(
        \registers[462][1] ) );
  EDFFX1 \registers_reg[462][0]  ( .D(n8038), .E(n28), .CK(clk), .Q(
        \registers[462][0] ) );
  EDFFX1 \registers_reg[458][7]  ( .D(n8425), .E(n24), .CK(clk), .Q(
        \registers[458][7] ) );
  EDFFX1 \registers_reg[458][6]  ( .D(n8367), .E(n24), .CK(clk), .Q(
        \registers[458][6] ) );
  EDFFX1 \registers_reg[458][5]  ( .D(n8309), .E(n24), .CK(clk), .Q(
        \registers[458][5] ) );
  EDFFX1 \registers_reg[458][4]  ( .D(n8251), .E(n24), .CK(clk), .Q(
        \registers[458][4] ) );
  EDFFX1 \registers_reg[458][3]  ( .D(n8198), .E(n24), .CK(clk), .Q(
        \registers[458][3] ) );
  EDFFX1 \registers_reg[458][2]  ( .D(n8152), .E(n24), .CK(clk), .Q(
        \registers[458][2] ) );
  EDFFX1 \registers_reg[458][1]  ( .D(n8096), .E(n24), .CK(clk), .Q(
        \registers[458][1] ) );
  EDFFX1 \registers_reg[458][0]  ( .D(n8039), .E(n24), .CK(clk), .Q(
        \registers[458][0] ) );
  EDFFX1 \registers_reg[454][7]  ( .D(n8424), .E(n251), .CK(clk), .Q(
        \registers[454][7] ) );
  EDFFX1 \registers_reg[454][6]  ( .D(n8366), .E(n251), .CK(clk), .Q(
        \registers[454][6] ) );
  EDFFX1 \registers_reg[454][5]  ( .D(n8308), .E(n251), .CK(clk), .Q(
        \registers[454][5] ) );
  EDFFX1 \registers_reg[454][4]  ( .D(n8250), .E(n251), .CK(clk), .Q(
        \registers[454][4] ) );
  EDFFX1 \registers_reg[454][3]  ( .D(n8199), .E(n251), .CK(clk), .Q(
        \registers[454][3] ) );
  EDFFX1 \registers_reg[454][2]  ( .D(n8153), .E(n251), .CK(clk), .Q(
        \registers[454][2] ) );
  EDFFX1 \registers_reg[454][1]  ( .D(n8097), .E(n251), .CK(clk), .Q(
        \registers[454][1] ) );
  EDFFX1 \registers_reg[454][0]  ( .D(n8037), .E(n251), .CK(clk), .Q(
        \registers[454][0] ) );
  EDFFX1 \registers_reg[450][7]  ( .D(n8422), .E(n247), .CK(clk), .Q(
        \registers[450][7] ) );
  EDFFX1 \registers_reg[450][6]  ( .D(n8364), .E(n247), .CK(clk), .Q(
        \registers[450][6] ) );
  EDFFX1 \registers_reg[450][5]  ( .D(n8306), .E(n247), .CK(clk), .Q(
        \registers[450][5] ) );
  EDFFX1 \registers_reg[450][4]  ( .D(n8248), .E(n247), .CK(clk), .Q(
        \registers[450][4] ) );
  EDFFX1 \registers_reg[450][3]  ( .D(n8197), .E(n247), .CK(clk), .Q(
        \registers[450][3] ) );
  EDFFX1 \registers_reg[450][2]  ( .D(n8154), .E(n247), .CK(clk), .Q(
        \registers[450][2] ) );
  EDFFX1 \registers_reg[450][1]  ( .D(n8098), .E(n247), .CK(clk), .Q(
        \registers[450][1] ) );
  EDFFX1 \registers_reg[450][0]  ( .D(n8038), .E(n247), .CK(clk), .Q(
        \registers[450][0] ) );
  EDFFX1 \registers_reg[446][7]  ( .D(n8424), .E(n716), .CK(clk), .Q(
        \registers[446][7] ) );
  EDFFX1 \registers_reg[446][6]  ( .D(n8366), .E(n716), .CK(clk), .Q(
        \registers[446][6] ) );
  EDFFX1 \registers_reg[446][5]  ( .D(n8308), .E(n716), .CK(clk), .Q(
        \registers[446][5] ) );
  EDFFX1 \registers_reg[446][4]  ( .D(n8250), .E(n716), .CK(clk), .Q(
        \registers[446][4] ) );
  EDFFX1 \registers_reg[446][3]  ( .D(n8199), .E(n716), .CK(clk), .Q(
        \registers[446][3] ) );
  EDFFX1 \registers_reg[446][2]  ( .D(n8153), .E(n716), .CK(clk), .Q(
        \registers[446][2] ) );
  EDFFX1 \registers_reg[446][1]  ( .D(n8097), .E(n716), .CK(clk), .Q(
        \registers[446][1] ) );
  EDFFX1 \registers_reg[446][0]  ( .D(n8037), .E(n716), .CK(clk), .Q(
        \registers[446][0] ) );
  EDFFX1 \registers_reg[442][7]  ( .D(n8422), .E(n712), .CK(clk), .Q(
        \registers[442][7] ) );
  EDFFX1 \registers_reg[442][6]  ( .D(n8364), .E(n712), .CK(clk), .Q(
        \registers[442][6] ) );
  EDFFX1 \registers_reg[442][5]  ( .D(n8306), .E(n712), .CK(clk), .Q(
        \registers[442][5] ) );
  EDFFX1 \registers_reg[442][4]  ( .D(n8248), .E(n712), .CK(clk), .Q(
        \registers[442][4] ) );
  EDFFX1 \registers_reg[442][3]  ( .D(n8197), .E(n712), .CK(clk), .Q(
        \registers[442][3] ) );
  EDFFX1 \registers_reg[442][2]  ( .D(n8154), .E(n712), .CK(clk), .Q(
        \registers[442][2] ) );
  EDFFX1 \registers_reg[442][1]  ( .D(n8098), .E(n712), .CK(clk), .Q(
        \registers[442][1] ) );
  EDFFX1 \registers_reg[442][0]  ( .D(n8038), .E(n712), .CK(clk), .Q(
        \registers[442][0] ) );
  EDFFX1 \registers_reg[438][7]  ( .D(n8423), .E(n708), .CK(clk), .Q(
        \registers[438][7] ) );
  EDFFX1 \registers_reg[438][6]  ( .D(n8365), .E(n708), .CK(clk), .Q(
        \registers[438][6] ) );
  EDFFX1 \registers_reg[438][5]  ( .D(n8307), .E(n708), .CK(clk), .Q(
        \registers[438][5] ) );
  EDFFX1 \registers_reg[438][4]  ( .D(n8249), .E(n708), .CK(clk), .Q(
        \registers[438][4] ) );
  EDFFX1 \registers_reg[438][3]  ( .D(n8198), .E(n708), .CK(clk), .Q(
        \registers[438][3] ) );
  EDFFX1 \registers_reg[438][2]  ( .D(n8152), .E(n708), .CK(clk), .Q(
        \registers[438][2] ) );
  EDFFX1 \registers_reg[438][1]  ( .D(n8096), .E(n708), .CK(clk), .Q(
        \registers[438][1] ) );
  EDFFX1 \registers_reg[438][0]  ( .D(n8039), .E(n708), .CK(clk), .Q(
        \registers[438][0] ) );
  EDFFX1 \registers_reg[434][7]  ( .D(n8424), .E(n20), .CK(clk), .Q(
        \registers[434][7] ) );
  EDFFX1 \registers_reg[434][6]  ( .D(n8366), .E(n20), .CK(clk), .Q(
        \registers[434][6] ) );
  EDFFX1 \registers_reg[434][5]  ( .D(n8308), .E(n20), .CK(clk), .Q(
        \registers[434][5] ) );
  EDFFX1 \registers_reg[434][4]  ( .D(n8250), .E(n20), .CK(clk), .Q(
        \registers[434][4] ) );
  EDFFX1 \registers_reg[434][3]  ( .D(n8199), .E(n20), .CK(clk), .Q(
        \registers[434][3] ) );
  EDFFX1 \registers_reg[434][2]  ( .D(n8153), .E(n20), .CK(clk), .Q(
        \registers[434][2] ) );
  EDFFX1 \registers_reg[434][1]  ( .D(n8097), .E(n20), .CK(clk), .Q(
        \registers[434][1] ) );
  EDFFX1 \registers_reg[434][0]  ( .D(n8037), .E(n20), .CK(clk), .Q(
        \registers[434][0] ) );
  EDFFX1 \registers_reg[430][7]  ( .D(n8422), .E(n16), .CK(clk), .Q(
        \registers[430][7] ) );
  EDFFX1 \registers_reg[430][6]  ( .D(n8364), .E(n16), .CK(clk), .Q(
        \registers[430][6] ) );
  EDFFX1 \registers_reg[430][5]  ( .D(n8306), .E(n16), .CK(clk), .Q(
        \registers[430][5] ) );
  EDFFX1 \registers_reg[430][4]  ( .D(n8248), .E(n16), .CK(clk), .Q(
        \registers[430][4] ) );
  EDFFX1 \registers_reg[430][3]  ( .D(n8197), .E(n16), .CK(clk), .Q(
        \registers[430][3] ) );
  EDFFX1 \registers_reg[430][2]  ( .D(n8154), .E(n16), .CK(clk), .Q(
        \registers[430][2] ) );
  EDFFX1 \registers_reg[430][1]  ( .D(n8098), .E(n16), .CK(clk), .Q(
        \registers[430][1] ) );
  EDFFX1 \registers_reg[430][0]  ( .D(n8038), .E(n16), .CK(clk), .Q(
        \registers[430][0] ) );
  EDFFX1 \registers_reg[426][7]  ( .D(n8423), .E(n12), .CK(clk), .Q(
        \registers[426][7] ) );
  EDFFX1 \registers_reg[426][6]  ( .D(n8365), .E(n12), .CK(clk), .Q(
        \registers[426][6] ) );
  EDFFX1 \registers_reg[426][5]  ( .D(n8307), .E(n12), .CK(clk), .Q(
        \registers[426][5] ) );
  EDFFX1 \registers_reg[426][4]  ( .D(n8249), .E(n12), .CK(clk), .Q(
        \registers[426][4] ) );
  EDFFX1 \registers_reg[426][3]  ( .D(n8198), .E(n12), .CK(clk), .Q(
        \registers[426][3] ) );
  EDFFX1 \registers_reg[426][2]  ( .D(n8152), .E(n12), .CK(clk), .Q(
        \registers[426][2] ) );
  EDFFX1 \registers_reg[426][1]  ( .D(n8096), .E(n12), .CK(clk), .Q(
        \registers[426][1] ) );
  EDFFX1 \registers_reg[426][0]  ( .D(n8039), .E(n12), .CK(clk), .Q(
        \registers[426][0] ) );
  EDFFX1 \registers_reg[422][7]  ( .D(n8424), .E(n244), .CK(clk), .Q(
        \registers[422][7] ) );
  EDFFX1 \registers_reg[422][6]  ( .D(n8366), .E(n244), .CK(clk), .Q(
        \registers[422][6] ) );
  EDFFX1 \registers_reg[422][5]  ( .D(n8308), .E(n244), .CK(clk), .Q(
        \registers[422][5] ) );
  EDFFX1 \registers_reg[422][4]  ( .D(n8250), .E(n244), .CK(clk), .Q(
        \registers[422][4] ) );
  EDFFX1 \registers_reg[422][3]  ( .D(n8196), .E(n244), .CK(clk), .Q(
        \registers[422][3] ) );
  EDFFX1 \registers_reg[422][2]  ( .D(n8151), .E(n244), .CK(clk), .Q(
        \registers[422][2] ) );
  EDFFX1 \registers_reg[422][1]  ( .D(n8095), .E(n244), .CK(clk), .Q(
        \registers[422][1] ) );
  EDFFX1 \registers_reg[422][0]  ( .D(n8034), .E(n244), .CK(clk), .Q(
        \registers[422][0] ) );
  EDFFX1 \registers_reg[418][7]  ( .D(n8422), .E(n240), .CK(clk), .Q(
        \registers[418][7] ) );
  EDFFX1 \registers_reg[418][6]  ( .D(n8364), .E(n240), .CK(clk), .Q(
        \registers[418][6] ) );
  EDFFX1 \registers_reg[418][5]  ( .D(n8306), .E(n240), .CK(clk), .Q(
        \registers[418][5] ) );
  EDFFX1 \registers_reg[418][4]  ( .D(n8248), .E(n240), .CK(clk), .Q(
        \registers[418][4] ) );
  EDFFX1 \registers_reg[418][3]  ( .D(n8194), .E(n240), .CK(clk), .Q(
        \registers[418][3] ) );
  EDFFX1 \registers_reg[418][2]  ( .D(n8726), .E(n240), .CK(clk), .Q(
        \registers[418][2] ) );
  EDFFX1 \registers_reg[418][1]  ( .D(n8698), .E(n240), .CK(clk), .Q(
        \registers[418][1] ) );
  EDFFX1 \registers_reg[418][0]  ( .D(n8035), .E(n240), .CK(clk), .Q(
        \registers[418][0] ) );
  EDFFX1 \registers_reg[414][7]  ( .D(n8423), .E(n704), .CK(clk), .Q(
        \registers[414][7] ) );
  EDFFX1 \registers_reg[414][6]  ( .D(n8365), .E(n704), .CK(clk), .Q(
        \registers[414][6] ) );
  EDFFX1 \registers_reg[414][5]  ( .D(n8307), .E(n704), .CK(clk), .Q(
        \registers[414][5] ) );
  EDFFX1 \registers_reg[414][4]  ( .D(n8249), .E(n704), .CK(clk), .Q(
        \registers[414][4] ) );
  EDFFX1 \registers_reg[414][3]  ( .D(n8195), .E(n704), .CK(clk), .Q(
        \registers[414][3] ) );
  EDFFX1 \registers_reg[414][2]  ( .D(n8150), .E(n704), .CK(clk), .Q(
        \registers[414][2] ) );
  EDFFX1 \registers_reg[414][1]  ( .D(n8094), .E(n704), .CK(clk), .Q(
        \registers[414][1] ) );
  EDFFX1 \registers_reg[414][0]  ( .D(n8036), .E(n704), .CK(clk), .Q(
        \registers[414][0] ) );
  EDFFX1 \registers_reg[410][7]  ( .D(n8424), .E(n700), .CK(clk), .Q(
        \registers[410][7] ) );
  EDFFX1 \registers_reg[410][6]  ( .D(n8366), .E(n700), .CK(clk), .Q(
        \registers[410][6] ) );
  EDFFX1 \registers_reg[410][5]  ( .D(n8308), .E(n700), .CK(clk), .Q(
        \registers[410][5] ) );
  EDFFX1 \registers_reg[410][4]  ( .D(n8250), .E(n700), .CK(clk), .Q(
        \registers[410][4] ) );
  EDFFX1 \registers_reg[410][3]  ( .D(n8196), .E(n700), .CK(clk), .Q(
        \registers[410][3] ) );
  EDFFX1 \registers_reg[410][2]  ( .D(n8151), .E(n700), .CK(clk), .Q(
        \registers[410][2] ) );
  EDFFX1 \registers_reg[410][1]  ( .D(n8095), .E(n700), .CK(clk), .Q(
        \registers[410][1] ) );
  EDFFX1 \registers_reg[410][0]  ( .D(n8034), .E(n700), .CK(clk), .Q(
        \registers[410][0] ) );
  EDFFX1 \registers_reg[406][7]  ( .D(n8420), .E(n696), .CK(clk), .Q(
        \registers[406][7] ) );
  EDFFX1 \registers_reg[406][6]  ( .D(n8362), .E(n696), .CK(clk), .Q(
        \registers[406][6] ) );
  EDFFX1 \registers_reg[406][5]  ( .D(n8304), .E(n696), .CK(clk), .Q(
        \registers[406][5] ) );
  EDFFX1 \registers_reg[406][4]  ( .D(n8246), .E(n696), .CK(clk), .Q(
        \registers[406][4] ) );
  EDFFX1 \registers_reg[406][3]  ( .D(n8194), .E(n696), .CK(clk), .Q(
        \registers[406][3] ) );
  EDFFX1 \registers_reg[406][2]  ( .D(n8724), .E(n696), .CK(clk), .Q(
        \registers[406][2] ) );
  EDFFX1 \registers_reg[406][1]  ( .D(n8696), .E(n696), .CK(clk), .Q(
        \registers[406][1] ) );
  EDFFX1 \registers_reg[406][0]  ( .D(n8035), .E(n696), .CK(clk), .Q(
        \registers[406][0] ) );
  EDFFX1 \registers_reg[402][7]  ( .D(n8421), .E(n692), .CK(clk), .Q(
        \registers[402][7] ) );
  EDFFX1 \registers_reg[402][6]  ( .D(n8363), .E(n692), .CK(clk), .Q(
        \registers[402][6] ) );
  EDFFX1 \registers_reg[402][5]  ( .D(n8305), .E(n692), .CK(clk), .Q(
        \registers[402][5] ) );
  EDFFX1 \registers_reg[402][4]  ( .D(n8247), .E(n692), .CK(clk), .Q(
        \registers[402][4] ) );
  EDFFX1 \registers_reg[402][3]  ( .D(n8195), .E(n692), .CK(clk), .Q(
        \registers[402][3] ) );
  EDFFX1 \registers_reg[402][2]  ( .D(n8150), .E(n692), .CK(clk), .Q(
        \registers[402][2] ) );
  EDFFX1 \registers_reg[402][1]  ( .D(n8094), .E(n692), .CK(clk), .Q(
        \registers[402][1] ) );
  EDFFX1 \registers_reg[402][0]  ( .D(n8036), .E(n692), .CK(clk), .Q(
        \registers[402][0] ) );
  EDFFX1 \registers_reg[398][7]  ( .D(n8419), .E(n688), .CK(clk), .Q(
        \registers[398][7] ) );
  EDFFX1 \registers_reg[398][6]  ( .D(n8361), .E(n688), .CK(clk), .Q(
        \registers[398][6] ) );
  EDFFX1 \registers_reg[398][5]  ( .D(n8303), .E(n688), .CK(clk), .Q(
        \registers[398][5] ) );
  EDFFX1 \registers_reg[398][4]  ( .D(n8245), .E(n688), .CK(clk), .Q(
        \registers[398][4] ) );
  EDFFX1 \registers_reg[398][3]  ( .D(n8196), .E(n688), .CK(clk), .Q(
        \registers[398][3] ) );
  EDFFX1 \registers_reg[398][2]  ( .D(n8151), .E(n688), .CK(clk), .Q(
        \registers[398][2] ) );
  EDFFX1 \registers_reg[398][1]  ( .D(n8095), .E(n688), .CK(clk), .Q(
        \registers[398][1] ) );
  EDFFX1 \registers_reg[398][0]  ( .D(n8034), .E(n688), .CK(clk), .Q(
        \registers[398][0] ) );
  EDFFX1 \registers_reg[394][7]  ( .D(n8420), .E(n684), .CK(clk), .Q(
        \registers[394][7] ) );
  EDFFX1 \registers_reg[394][6]  ( .D(n8362), .E(n684), .CK(clk), .Q(
        \registers[394][6] ) );
  EDFFX1 \registers_reg[394][5]  ( .D(n8304), .E(n684), .CK(clk), .Q(
        \registers[394][5] ) );
  EDFFX1 \registers_reg[394][4]  ( .D(n8246), .E(n684), .CK(clk), .Q(
        \registers[394][4] ) );
  EDFFX1 \registers_reg[394][3]  ( .D(n8194), .E(n684), .CK(clk), .Q(
        \registers[394][3] ) );
  EDFFX1 \registers_reg[394][2]  ( .D(n8729), .E(n684), .CK(clk), .Q(
        \registers[394][2] ) );
  EDFFX1 \registers_reg[394][1]  ( .D(n8701), .E(n684), .CK(clk), .Q(
        \registers[394][1] ) );
  EDFFX1 \registers_reg[394][0]  ( .D(n8035), .E(n684), .CK(clk), .Q(
        \registers[394][0] ) );
  EDFFX1 \registers_reg[390][7]  ( .D(n8421), .E(n1000), .CK(clk), .Q(
        \registers[390][7] ) );
  EDFFX1 \registers_reg[390][6]  ( .D(n8363), .E(n1000), .CK(clk), .Q(
        \registers[390][6] ) );
  EDFFX1 \registers_reg[390][5]  ( .D(n8305), .E(n1000), .CK(clk), .Q(
        \registers[390][5] ) );
  EDFFX1 \registers_reg[390][4]  ( .D(n8247), .E(n1000), .CK(clk), .Q(
        \registers[390][4] ) );
  EDFFX1 \registers_reg[390][3]  ( .D(n8195), .E(n1000), .CK(clk), .Q(
        \registers[390][3] ) );
  EDFFX1 \registers_reg[390][2]  ( .D(n8150), .E(n1000), .CK(clk), .Q(
        \registers[390][2] ) );
  EDFFX1 \registers_reg[390][1]  ( .D(n8094), .E(n1000), .CK(clk), .Q(
        \registers[390][1] ) );
  EDFFX1 \registers_reg[390][0]  ( .D(n8036), .E(n1000), .CK(clk), .Q(
        \registers[390][0] ) );
  EDFFX1 \registers_reg[386][7]  ( .D(n8419), .E(n996), .CK(clk), .Q(
        \registers[386][7] ) );
  EDFFX1 \registers_reg[386][6]  ( .D(n8361), .E(n996), .CK(clk), .Q(
        \registers[386][6] ) );
  EDFFX1 \registers_reg[386][5]  ( .D(n8303), .E(n996), .CK(clk), .Q(
        \registers[386][5] ) );
  EDFFX1 \registers_reg[386][4]  ( .D(n8245), .E(n996), .CK(clk), .Q(
        \registers[386][4] ) );
  EDFFX1 \registers_reg[386][3]  ( .D(n8196), .E(n996), .CK(clk), .Q(
        \registers[386][3] ) );
  EDFFX1 \registers_reg[386][2]  ( .D(n8151), .E(n996), .CK(clk), .Q(
        \registers[386][2] ) );
  EDFFX1 \registers_reg[386][1]  ( .D(n8095), .E(n996), .CK(clk), .Q(
        \registers[386][1] ) );
  EDFFX1 \registers_reg[386][0]  ( .D(n8034), .E(n996), .CK(clk), .Q(
        \registers[386][0] ) );
  EDFFX1 \registers_reg[382][7]  ( .D(n8434), .E(n680), .CK(clk), .Q(
        \registers[382][7] ) );
  EDFFX1 \registers_reg[382][6]  ( .D(n8376), .E(n680), .CK(clk), .Q(
        \registers[382][6] ) );
  EDFFX1 \registers_reg[382][5]  ( .D(n8318), .E(n680), .CK(clk), .Q(
        \registers[382][5] ) );
  EDFFX1 \registers_reg[382][4]  ( .D(n8260), .E(n680), .CK(clk), .Q(
        \registers[382][4] ) );
  EDFFX1 \registers_reg[382][3]  ( .D(n8172), .E(n680), .CK(clk), .Q(
        \registers[382][3] ) );
  EDFFX1 \registers_reg[382][2]  ( .D(n8108), .E(n680), .CK(clk), .Q(
        \registers[382][2] ) );
  EDFFX1 \registers_reg[382][1]  ( .D(n8052), .E(n680), .CK(clk), .Q(
        \registers[382][1] ) );
  EDFFX1 \registers_reg[382][0]  ( .D(n8005), .E(n680), .CK(clk), .Q(
        \registers[382][0] ) );
  EDFFX1 \registers_reg[378][7]  ( .D(n8434), .E(n676), .CK(clk), .Q(
        \registers[378][7] ) );
  EDFFX1 \registers_reg[378][6]  ( .D(n8376), .E(n676), .CK(clk), .Q(
        \registers[378][6] ) );
  EDFFX1 \registers_reg[378][5]  ( .D(n8318), .E(n676), .CK(clk), .Q(
        \registers[378][5] ) );
  EDFFX1 \registers_reg[378][4]  ( .D(n8260), .E(n676), .CK(clk), .Q(
        \registers[378][4] ) );
  EDFFX1 \registers_reg[378][3]  ( .D(n8185), .E(n676), .CK(clk), .Q(
        \registers[378][3] ) );
  EDFFX1 \registers_reg[378][2]  ( .D(n8109), .E(n676), .CK(clk), .Q(
        \registers[378][2] ) );
  EDFFX1 \registers_reg[378][1]  ( .D(n8053), .E(n676), .CK(clk), .Q(
        \registers[378][1] ) );
  EDFFX1 \registers_reg[378][0]  ( .D(n8000), .E(n676), .CK(clk), .Q(
        \registers[378][0] ) );
  EDFFX1 \registers_reg[374][7]  ( .D(n8433), .E(n672), .CK(clk), .Q(
        \registers[374][7] ) );
  EDFFX1 \registers_reg[374][6]  ( .D(n8375), .E(n672), .CK(clk), .Q(
        \registers[374][6] ) );
  EDFFX1 \registers_reg[374][5]  ( .D(n8317), .E(n672), .CK(clk), .Q(
        \registers[374][5] ) );
  EDFFX1 \registers_reg[374][4]  ( .D(n8259), .E(n672), .CK(clk), .Q(
        \registers[374][4] ) );
  EDFFX1 \registers_reg[374][3]  ( .D(n8187), .E(n672), .CK(clk), .Q(
        \registers[374][3] ) );
  EDFFX1 \registers_reg[374][2]  ( .D(n8110), .E(n672), .CK(clk), .Q(
        \registers[374][2] ) );
  EDFFX1 \registers_reg[374][1]  ( .D(n8054), .E(n672), .CK(clk), .Q(
        \registers[374][1] ) );
  EDFFX1 \registers_reg[374][0]  ( .D(n8006), .E(n672), .CK(clk), .Q(
        \registers[374][0] ) );
  EDFFX1 \registers_reg[370][7]  ( .D(n8434), .E(n668), .CK(clk), .Q(
        \registers[370][7] ) );
  EDFFX1 \registers_reg[370][6]  ( .D(n8376), .E(n668), .CK(clk), .Q(
        \registers[370][6] ) );
  EDFFX1 \registers_reg[370][5]  ( .D(n8318), .E(n668), .CK(clk), .Q(
        \registers[370][5] ) );
  EDFFX1 \registers_reg[370][4]  ( .D(n8260), .E(n668), .CK(clk), .Q(
        \registers[370][4] ) );
  EDFFX1 \registers_reg[370][3]  ( .D(n8173), .E(n668), .CK(clk), .Q(
        \registers[370][3] ) );
  EDFFX1 \registers_reg[370][2]  ( .D(n8158), .E(n668), .CK(clk), .Q(
        \registers[370][2] ) );
  EDFFX1 \registers_reg[370][1]  ( .D(n8102), .E(n668), .CK(clk), .Q(
        \registers[370][1] ) );
  EDFFX1 \registers_reg[370][0]  ( .D(n8046), .E(n668), .CK(clk), .Q(
        \registers[370][0] ) );
  EDFFX1 \registers_reg[366][7]  ( .D(n8433), .E(n664), .CK(clk), .Q(
        \registers[366][7] ) );
  EDFFX1 \registers_reg[366][6]  ( .D(n8375), .E(n664), .CK(clk), .Q(
        \registers[366][6] ) );
  EDFFX1 \registers_reg[366][5]  ( .D(n8317), .E(n664), .CK(clk), .Q(
        \registers[366][5] ) );
  EDFFX1 \registers_reg[366][4]  ( .D(n8259), .E(n664), .CK(clk), .Q(
        \registers[366][4] ) );
  EDFFX1 \registers_reg[366][3]  ( .D(n8186), .E(n664), .CK(clk), .Q(
        \registers[366][3] ) );
  EDFFX1 \registers_reg[366][2]  ( .D(n8117), .E(n664), .CK(clk), .Q(
        \registers[366][2] ) );
  EDFFX1 \registers_reg[366][1]  ( .D(n8061), .E(n664), .CK(clk), .Q(
        \registers[366][1] ) );
  EDFFX1 \registers_reg[366][0]  ( .D(n8047), .E(n664), .CK(clk), .Q(
        \registers[366][0] ) );
  EDFFX1 \registers_reg[362][7]  ( .D(n8433), .E(n660), .CK(clk), .Q(
        \registers[362][7] ) );
  EDFFX1 \registers_reg[362][6]  ( .D(n8375), .E(n660), .CK(clk), .Q(
        \registers[362][6] ) );
  EDFFX1 \registers_reg[362][5]  ( .D(n8317), .E(n660), .CK(clk), .Q(
        \registers[362][5] ) );
  EDFFX1 \registers_reg[362][4]  ( .D(n8259), .E(n660), .CK(clk), .Q(
        \registers[362][4] ) );
  EDFFX1 \registers_reg[362][3]  ( .D(n8768), .E(n660), .CK(clk), .Q(
        \registers[362][3] ) );
  EDFFX1 \registers_reg[362][2]  ( .D(n8148), .E(n660), .CK(clk), .Q(
        \registers[362][2] ) );
  EDFFX1 \registers_reg[362][1]  ( .D(n8092), .E(n660), .CK(clk), .Q(
        \registers[362][1] ) );
  EDFFX1 \registers_reg[362][0]  ( .D(n8048), .E(n660), .CK(clk), .Q(
        \registers[362][0] ) );
  EDFFX1 \registers_reg[358][7]  ( .D(n8434), .E(n993), .CK(clk), .Q(
        \registers[358][7] ) );
  EDFFX1 \registers_reg[358][6]  ( .D(n8376), .E(n993), .CK(clk), .Q(
        \registers[358][6] ) );
  EDFFX1 \registers_reg[358][5]  ( .D(n8318), .E(n993), .CK(clk), .Q(
        \registers[358][5] ) );
  EDFFX1 \registers_reg[358][4]  ( .D(n8260), .E(n993), .CK(clk), .Q(
        \registers[358][4] ) );
  EDFFX1 \registers_reg[358][3]  ( .D(n8768), .E(n993), .CK(clk), .Q(
        \registers[358][3] ) );
  EDFFX1 \registers_reg[358][2]  ( .D(n8152), .E(n993), .CK(clk), .Q(
        \registers[358][2] ) );
  EDFFX1 \registers_reg[358][1]  ( .D(n8096), .E(n993), .CK(clk), .Q(
        \registers[358][1] ) );
  EDFFX1 \registers_reg[358][0]  ( .D(n8046), .E(n993), .CK(clk), .Q(
        \registers[358][0] ) );
  EDFFX1 \registers_reg[354][7]  ( .D(n8434), .E(n989), .CK(clk), .Q(
        \registers[354][7] ) );
  EDFFX1 \registers_reg[354][6]  ( .D(n8376), .E(n989), .CK(clk), .Q(
        \registers[354][6] ) );
  EDFFX1 \registers_reg[354][5]  ( .D(n8318), .E(n989), .CK(clk), .Q(
        \registers[354][5] ) );
  EDFFX1 \registers_reg[354][4]  ( .D(n8260), .E(n989), .CK(clk), .Q(
        \registers[354][4] ) );
  EDFFX1 \registers_reg[354][3]  ( .D(n8174), .E(n989), .CK(clk), .Q(
        \registers[354][3] ) );
  EDFFX1 \registers_reg[354][2]  ( .D(n8118), .E(n989), .CK(clk), .Q(
        \registers[354][2] ) );
  EDFFX1 \registers_reg[354][1]  ( .D(n8062), .E(n989), .CK(clk), .Q(
        \registers[354][1] ) );
  EDFFX1 \registers_reg[354][0]  ( .D(n8047), .E(n989), .CK(clk), .Q(
        \registers[354][0] ) );
  EDFFX1 \registers_reg[350][7]  ( .D(n8431), .E(n656), .CK(clk), .Q(
        \registers[350][7] ) );
  EDFFX1 \registers_reg[350][6]  ( .D(n8373), .E(n656), .CK(clk), .Q(
        \registers[350][6] ) );
  EDFFX1 \registers_reg[350][5]  ( .D(n8315), .E(n656), .CK(clk), .Q(
        \registers[350][5] ) );
  EDFFX1 \registers_reg[350][4]  ( .D(n8257), .E(n656), .CK(clk), .Q(
        \registers[350][4] ) );
  EDFFX1 \registers_reg[350][3]  ( .D(n8202), .E(n656), .CK(clk), .Q(
        \registers[350][3] ) );
  EDFFX1 \registers_reg[350][2]  ( .D(n8149), .E(n656), .CK(clk), .Q(
        \registers[350][2] ) );
  EDFFX1 \registers_reg[350][1]  ( .D(n8093), .E(n656), .CK(clk), .Q(
        \registers[350][1] ) );
  EDFFX1 \registers_reg[350][0]  ( .D(n8048), .E(n656), .CK(clk), .Q(
        \registers[350][0] ) );
  EDFFX1 \registers_reg[346][7]  ( .D(n8432), .E(n652), .CK(clk), .Q(
        \registers[346][7] ) );
  EDFFX1 \registers_reg[346][6]  ( .D(n8374), .E(n652), .CK(clk), .Q(
        \registers[346][6] ) );
  EDFFX1 \registers_reg[346][5]  ( .D(n8316), .E(n652), .CK(clk), .Q(
        \registers[346][5] ) );
  EDFFX1 \registers_reg[346][4]  ( .D(n8258), .E(n652), .CK(clk), .Q(
        \registers[346][4] ) );
  EDFFX1 \registers_reg[346][3]  ( .D(n8168), .E(n652), .CK(clk), .Q(
        \registers[346][3] ) );
  EDFFX1 \registers_reg[346][2]  ( .D(n8153), .E(n652), .CK(clk), .Q(
        \registers[346][2] ) );
  EDFFX1 \registers_reg[346][1]  ( .D(n8097), .E(n652), .CK(clk), .Q(
        \registers[346][1] ) );
  EDFFX1 \registers_reg[346][0]  ( .D(n8046), .E(n652), .CK(clk), .Q(
        \registers[346][0] ) );
  EDFFX1 \registers_reg[342][7]  ( .D(n8430), .E(n648), .CK(clk), .Q(
        \registers[342][7] ) );
  EDFFX1 \registers_reg[342][6]  ( .D(n8372), .E(n648), .CK(clk), .Q(
        \registers[342][6] ) );
  EDFFX1 \registers_reg[342][5]  ( .D(n8314), .E(n648), .CK(clk), .Q(
        \registers[342][5] ) );
  EDFFX1 \registers_reg[342][4]  ( .D(n8256), .E(n648), .CK(clk), .Q(
        \registers[342][4] ) );
  EDFFX1 \registers_reg[342][3]  ( .D(n8175), .E(n648), .CK(clk), .Q(
        \registers[342][3] ) );
  EDFFX1 \registers_reg[342][2]  ( .D(n8119), .E(n648), .CK(clk), .Q(
        \registers[342][2] ) );
  EDFFX1 \registers_reg[342][1]  ( .D(n8063), .E(n648), .CK(clk), .Q(
        \registers[342][1] ) );
  EDFFX1 \registers_reg[342][0]  ( .D(n8047), .E(n648), .CK(clk), .Q(
        \registers[342][0] ) );
  EDFFX1 \registers_reg[338][7]  ( .D(n8431), .E(n644), .CK(clk), .Q(
        \registers[338][7] ) );
  EDFFX1 \registers_reg[338][6]  ( .D(n8373), .E(n644), .CK(clk), .Q(
        \registers[338][6] ) );
  EDFFX1 \registers_reg[338][5]  ( .D(n8315), .E(n644), .CK(clk), .Q(
        \registers[338][5] ) );
  EDFFX1 \registers_reg[338][4]  ( .D(n8257), .E(n644), .CK(clk), .Q(
        \registers[338][4] ) );
  EDFFX1 \registers_reg[338][3]  ( .D(n8200), .E(n644), .CK(clk), .Q(
        \registers[338][3] ) );
  EDFFX1 \registers_reg[338][2]  ( .D(n8144), .E(n644), .CK(clk), .Q(
        \registers[338][2] ) );
  EDFFX1 \registers_reg[338][1]  ( .D(n8088), .E(n644), .CK(clk), .Q(
        \registers[338][1] ) );
  EDFFX1 \registers_reg[338][0]  ( .D(n8048), .E(n644), .CK(clk), .Q(
        \registers[338][0] ) );
  EDFFX1 \registers_reg[334][7]  ( .D(n8432), .E(n640), .CK(clk), .Q(
        \registers[334][7] ) );
  EDFFX1 \registers_reg[334][6]  ( .D(n8374), .E(n640), .CK(clk), .Q(
        \registers[334][6] ) );
  EDFFX1 \registers_reg[334][5]  ( .D(n8316), .E(n640), .CK(clk), .Q(
        \registers[334][5] ) );
  EDFFX1 \registers_reg[334][4]  ( .D(n8258), .E(n640), .CK(clk), .Q(
        \registers[334][4] ) );
  EDFFX1 \registers_reg[334][3]  ( .D(n8169), .E(n640), .CK(clk), .Q(
        \registers[334][3] ) );
  EDFFX1 \registers_reg[334][2]  ( .D(n8154), .E(n640), .CK(clk), .Q(
        \registers[334][2] ) );
  EDFFX1 \registers_reg[334][1]  ( .D(n8098), .E(n640), .CK(clk), .Q(
        \registers[334][1] ) );
  EDFFX1 \registers_reg[334][0]  ( .D(n8046), .E(n640), .CK(clk), .Q(
        \registers[334][0] ) );
  EDFFX1 \registers_reg[330][7]  ( .D(n8430), .E(n636), .CK(clk), .Q(
        \registers[330][7] ) );
  EDFFX1 \registers_reg[330][6]  ( .D(n8372), .E(n636), .CK(clk), .Q(
        \registers[330][6] ) );
  EDFFX1 \registers_reg[330][5]  ( .D(n8314), .E(n636), .CK(clk), .Q(
        \registers[330][5] ) );
  EDFFX1 \registers_reg[330][4]  ( .D(n8256), .E(n636), .CK(clk), .Q(
        \registers[330][4] ) );
  EDFFX1 \registers_reg[330][3]  ( .D(n8188), .E(n636), .CK(clk), .Q(
        \registers[330][3] ) );
  EDFFX1 \registers_reg[330][2]  ( .D(n8114), .E(n636), .CK(clk), .Q(
        \registers[330][2] ) );
  EDFFX1 \registers_reg[330][1]  ( .D(n8058), .E(n636), .CK(clk), .Q(
        \registers[330][1] ) );
  EDFFX1 \registers_reg[330][0]  ( .D(n8047), .E(n636), .CK(clk), .Q(
        \registers[330][0] ) );
  EDFFX1 \registers_reg[326][7]  ( .D(n8431), .E(n986), .CK(clk), .Q(
        \registers[326][7] ) );
  EDFFX1 \registers_reg[326][6]  ( .D(n8373), .E(n986), .CK(clk), .Q(
        \registers[326][6] ) );
  EDFFX1 \registers_reg[326][5]  ( .D(n8315), .E(n986), .CK(clk), .Q(
        \registers[326][5] ) );
  EDFFX1 \registers_reg[326][4]  ( .D(n8257), .E(n986), .CK(clk), .Q(
        \registers[326][4] ) );
  EDFFX1 \registers_reg[326][3]  ( .D(n8201), .E(n986), .CK(clk), .Q(
        \registers[326][3] ) );
  EDFFX1 \registers_reg[326][2]  ( .D(n8146), .E(n986), .CK(clk), .Q(
        \registers[326][2] ) );
  EDFFX1 \registers_reg[326][1]  ( .D(n8090), .E(n986), .CK(clk), .Q(
        \registers[326][1] ) );
  EDFFX1 \registers_reg[326][0]  ( .D(n8048), .E(n986), .CK(clk), .Q(
        \registers[326][0] ) );
  EDFFX1 \registers_reg[322][7]  ( .D(n8432), .E(n982), .CK(clk), .Q(
        \registers[322][7] ) );
  EDFFX1 \registers_reg[322][6]  ( .D(n8374), .E(n982), .CK(clk), .Q(
        \registers[322][6] ) );
  EDFFX1 \registers_reg[322][5]  ( .D(n8316), .E(n982), .CK(clk), .Q(
        \registers[322][5] ) );
  EDFFX1 \registers_reg[322][4]  ( .D(n8258), .E(n982), .CK(clk), .Q(
        \registers[322][4] ) );
  EDFFX1 \registers_reg[322][3]  ( .D(n8166), .E(n982), .CK(clk), .Q(
        \registers[322][3] ) );
  EDFFX1 \registers_reg[322][2]  ( .D(n8150), .E(n982), .CK(clk), .Q(
        \registers[322][2] ) );
  EDFFX1 \registers_reg[322][1]  ( .D(n8094), .E(n982), .CK(clk), .Q(
        \registers[322][1] ) );
  EDFFX1 \registers_reg[322][0]  ( .D(n8046), .E(n982), .CK(clk), .Q(
        \registers[322][0] ) );
  EDFFX1 \registers_reg[318][7]  ( .D(n8431), .E(n632), .CK(clk), .Q(
        \registers[318][7] ) );
  EDFFX1 \registers_reg[318][6]  ( .D(n8373), .E(n632), .CK(clk), .Q(
        \registers[318][6] ) );
  EDFFX1 \registers_reg[318][5]  ( .D(n8315), .E(n632), .CK(clk), .Q(
        \registers[318][5] ) );
  EDFFX1 \registers_reg[318][4]  ( .D(n8257), .E(n632), .CK(clk), .Q(
        \registers[318][4] ) );
  EDFFX1 \registers_reg[318][3]  ( .D(n8197), .E(n632), .CK(clk), .Q(
        \registers[318][3] ) );
  EDFFX1 \registers_reg[318][2]  ( .D(n8158), .E(n632), .CK(clk), .Q(
        \registers[318][2] ) );
  EDFFX1 \registers_reg[318][1]  ( .D(n8102), .E(n632), .CK(clk), .Q(
        \registers[318][1] ) );
  EDFFX1 \registers_reg[318][0]  ( .D(n8045), .E(n632), .CK(clk), .Q(
        \registers[318][0] ) );
  EDFFX1 \registers_reg[314][7]  ( .D(n8432), .E(n628), .CK(clk), .Q(
        \registers[314][7] ) );
  EDFFX1 \registers_reg[314][6]  ( .D(n8374), .E(n628), .CK(clk), .Q(
        \registers[314][6] ) );
  EDFFX1 \registers_reg[314][5]  ( .D(n8316), .E(n628), .CK(clk), .Q(
        \registers[314][5] ) );
  EDFFX1 \registers_reg[314][4]  ( .D(n8258), .E(n628), .CK(clk), .Q(
        \registers[314][4] ) );
  EDFFX1 \registers_reg[314][3]  ( .D(n8164), .E(n628), .CK(clk), .Q(
        \registers[314][3] ) );
  EDFFX1 \registers_reg[314][2]  ( .D(n8159), .E(n628), .CK(clk), .Q(
        \registers[314][2] ) );
  EDFFX1 \registers_reg[314][1]  ( .D(n8103), .E(n628), .CK(clk), .Q(
        \registers[314][1] ) );
  EDFFX1 \registers_reg[314][0]  ( .D(n8043), .E(n628), .CK(clk), .Q(
        \registers[314][0] ) );
  EDFFX1 \registers_reg[310][7]  ( .D(n8430), .E(n624), .CK(clk), .Q(
        \registers[310][7] ) );
  EDFFX1 \registers_reg[310][6]  ( .D(n8372), .E(n624), .CK(clk), .Q(
        \registers[310][6] ) );
  EDFFX1 \registers_reg[310][5]  ( .D(n8314), .E(n624), .CK(clk), .Q(
        \registers[310][5] ) );
  EDFFX1 \registers_reg[310][4]  ( .D(n8256), .E(n624), .CK(clk), .Q(
        \registers[310][4] ) );
  EDFFX1 \registers_reg[310][3]  ( .D(n8189), .E(n624), .CK(clk), .Q(
        \registers[310][3] ) );
  EDFFX1 \registers_reg[310][2]  ( .D(n8160), .E(n624), .CK(clk), .Q(
        \registers[310][2] ) );
  EDFFX1 \registers_reg[310][1]  ( .D(n8104), .E(n624), .CK(clk), .Q(
        \registers[310][1] ) );
  EDFFX1 \registers_reg[310][0]  ( .D(n8044), .E(n624), .CK(clk), .Q(
        \registers[310][0] ) );
  EDFFX1 \registers_reg[306][7]  ( .D(n8431), .E(n620), .CK(clk), .Q(
        \registers[306][7] ) );
  EDFFX1 \registers_reg[306][6]  ( .D(n8373), .E(n620), .CK(clk), .Q(
        \registers[306][6] ) );
  EDFFX1 \registers_reg[306][5]  ( .D(n8315), .E(n620), .CK(clk), .Q(
        \registers[306][5] ) );
  EDFFX1 \registers_reg[306][4]  ( .D(n8257), .E(n620), .CK(clk), .Q(
        \registers[306][4] ) );
  EDFFX1 \registers_reg[306][3]  ( .D(n8198), .E(n620), .CK(clk), .Q(
        \registers[306][3] ) );
  EDFFX1 \registers_reg[306][2]  ( .D(n8158), .E(n620), .CK(clk), .Q(
        \registers[306][2] ) );
  EDFFX1 \registers_reg[306][1]  ( .D(n8102), .E(n620), .CK(clk), .Q(
        \registers[306][1] ) );
  EDFFX1 \registers_reg[306][0]  ( .D(n8045), .E(n620), .CK(clk), .Q(
        \registers[306][0] ) );
  EDFFX1 \registers_reg[302][7]  ( .D(n8428), .E(n616), .CK(clk), .Q(
        \registers[302][7] ) );
  EDFFX1 \registers_reg[302][6]  ( .D(n8370), .E(n616), .CK(clk), .Q(
        \registers[302][6] ) );
  EDFFX1 \registers_reg[302][5]  ( .D(n8312), .E(n616), .CK(clk), .Q(
        \registers[302][5] ) );
  EDFFX1 \registers_reg[302][4]  ( .D(n8254), .E(n616), .CK(clk), .Q(
        \registers[302][4] ) );
  EDFFX1 \registers_reg[302][3]  ( .D(n8165), .E(n616), .CK(clk), .Q(
        \registers[302][3] ) );
  EDFFX1 \registers_reg[302][2]  ( .D(n8159), .E(n616), .CK(clk), .Q(
        \registers[302][2] ) );
  EDFFX1 \registers_reg[302][1]  ( .D(n8103), .E(n616), .CK(clk), .Q(
        \registers[302][1] ) );
  EDFFX1 \registers_reg[302][0]  ( .D(n8043), .E(n616), .CK(clk), .Q(
        \registers[302][0] ) );
  EDFFX1 \registers_reg[298][7]  ( .D(n8429), .E(n612), .CK(clk), .Q(
        \registers[298][7] ) );
  EDFFX1 \registers_reg[298][6]  ( .D(n8371), .E(n612), .CK(clk), .Q(
        \registers[298][6] ) );
  EDFFX1 \registers_reg[298][5]  ( .D(n8313), .E(n612), .CK(clk), .Q(
        \registers[298][5] ) );
  EDFFX1 \registers_reg[298][4]  ( .D(n8255), .E(n612), .CK(clk), .Q(
        \registers[298][4] ) );
  EDFFX1 \registers_reg[298][3]  ( .D(n8190), .E(n612), .CK(clk), .Q(
        \registers[298][3] ) );
  EDFFX1 \registers_reg[298][2]  ( .D(n8160), .E(n612), .CK(clk), .Q(
        \registers[298][2] ) );
  EDFFX1 \registers_reg[298][1]  ( .D(n8104), .E(n612), .CK(clk), .Q(
        \registers[298][1] ) );
  EDFFX1 \registers_reg[298][0]  ( .D(n8044), .E(n612), .CK(clk), .Q(
        \registers[298][0] ) );
  EDFFX1 \registers_reg[294][7]  ( .D(n8427), .E(n979), .CK(clk), .Q(
        \registers[294][7] ) );
  EDFFX1 \registers_reg[294][6]  ( .D(n8369), .E(n979), .CK(clk), .Q(
        \registers[294][6] ) );
  EDFFX1 \registers_reg[294][5]  ( .D(n8311), .E(n979), .CK(clk), .Q(
        \registers[294][5] ) );
  EDFFX1 \registers_reg[294][4]  ( .D(n8253), .E(n979), .CK(clk), .Q(
        \registers[294][4] ) );
  EDFFX1 \registers_reg[294][3]  ( .D(n8201), .E(n979), .CK(clk), .Q(
        \registers[294][3] ) );
  EDFFX1 \registers_reg[294][2]  ( .D(n8158), .E(n979), .CK(clk), .Q(
        \registers[294][2] ) );
  EDFFX1 \registers_reg[294][1]  ( .D(n8102), .E(n979), .CK(clk), .Q(
        \registers[294][1] ) );
  EDFFX1 \registers_reg[294][0]  ( .D(n8045), .E(n979), .CK(clk), .Q(
        \registers[294][0] ) );
  EDFFX1 \registers_reg[290][7]  ( .D(n8428), .E(n975), .CK(clk), .Q(
        \registers[290][7] ) );
  EDFFX1 \registers_reg[290][6]  ( .D(n8370), .E(n975), .CK(clk), .Q(
        \registers[290][6] ) );
  EDFFX1 \registers_reg[290][5]  ( .D(n8312), .E(n975), .CK(clk), .Q(
        \registers[290][5] ) );
  EDFFX1 \registers_reg[290][4]  ( .D(n8254), .E(n975), .CK(clk), .Q(
        \registers[290][4] ) );
  EDFFX1 \registers_reg[290][3]  ( .D(n8202), .E(n975), .CK(clk), .Q(
        \registers[290][3] ) );
  EDFFX1 \registers_reg[290][2]  ( .D(n8159), .E(n975), .CK(clk), .Q(
        \registers[290][2] ) );
  EDFFX1 \registers_reg[290][1]  ( .D(n8103), .E(n975), .CK(clk), .Q(
        \registers[290][1] ) );
  EDFFX1 \registers_reg[290][0]  ( .D(n8043), .E(n975), .CK(clk), .Q(
        \registers[290][0] ) );
  EDFFX1 \registers_reg[286][7]  ( .D(n8429), .E(n608), .CK(clk), .Q(
        \registers[286][7] ) );
  EDFFX1 \registers_reg[286][6]  ( .D(n8371), .E(n608), .CK(clk), .Q(
        \registers[286][6] ) );
  EDFFX1 \registers_reg[286][5]  ( .D(n8313), .E(n608), .CK(clk), .Q(
        \registers[286][5] ) );
  EDFFX1 \registers_reg[286][4]  ( .D(n8255), .E(n608), .CK(clk), .Q(
        \registers[286][4] ) );
  EDFFX1 \registers_reg[286][3]  ( .D(n8200), .E(n608), .CK(clk), .Q(
        \registers[286][3] ) );
  EDFFX1 \registers_reg[286][2]  ( .D(n8160), .E(n608), .CK(clk), .Q(
        \registers[286][2] ) );
  EDFFX1 \registers_reg[286][1]  ( .D(n8104), .E(n608), .CK(clk), .Q(
        \registers[286][1] ) );
  EDFFX1 \registers_reg[286][0]  ( .D(n8044), .E(n608), .CK(clk), .Q(
        \registers[286][0] ) );
  EDFFX1 \registers_reg[282][7]  ( .D(n8874), .E(n604), .CK(clk), .Q(
        \registers[282][7] ) );
  EDFFX1 \registers_reg[282][6]  ( .D(n8845), .E(n604), .CK(clk), .Q(
        \registers[282][6] ) );
  EDFFX1 \registers_reg[282][5]  ( .D(n8816), .E(n604), .CK(clk), .Q(
        \registers[282][5] ) );
  EDFFX1 \registers_reg[282][4]  ( .D(n8787), .E(n604), .CK(clk), .Q(
        \registers[282][4] ) );
  EDFFX1 \registers_reg[282][3]  ( .D(n8201), .E(n604), .CK(clk), .Q(
        \registers[282][3] ) );
  EDFFX1 \registers_reg[282][2]  ( .D(n8158), .E(n604), .CK(clk), .Q(
        \registers[282][2] ) );
  EDFFX1 \registers_reg[282][1]  ( .D(n8102), .E(n604), .CK(clk), .Q(
        \registers[282][1] ) );
  EDFFX1 \registers_reg[282][0]  ( .D(n8045), .E(n604), .CK(clk), .Q(
        \registers[282][0] ) );
  EDFFX1 \registers_reg[278][7]  ( .D(n8428), .E(n600), .CK(clk), .Q(
        \registers[278][7] ) );
  EDFFX1 \registers_reg[278][6]  ( .D(n8370), .E(n600), .CK(clk), .Q(
        \registers[278][6] ) );
  EDFFX1 \registers_reg[278][5]  ( .D(n8312), .E(n600), .CK(clk), .Q(
        \registers[278][5] ) );
  EDFFX1 \registers_reg[278][4]  ( .D(n8254), .E(n600), .CK(clk), .Q(
        \registers[278][4] ) );
  EDFFX1 \registers_reg[278][3]  ( .D(n8202), .E(n600), .CK(clk), .Q(
        \registers[278][3] ) );
  EDFFX1 \registers_reg[278][2]  ( .D(n8159), .E(n600), .CK(clk), .Q(
        \registers[278][2] ) );
  EDFFX1 \registers_reg[278][1]  ( .D(n8103), .E(n600), .CK(clk), .Q(
        \registers[278][1] ) );
  EDFFX1 \registers_reg[278][0]  ( .D(n8043), .E(n600), .CK(clk), .Q(
        \registers[278][0] ) );
  EDFFX1 \registers_reg[274][7]  ( .D(n8429), .E(n596), .CK(clk), .Q(
        \registers[274][7] ) );
  EDFFX1 \registers_reg[274][6]  ( .D(n8371), .E(n596), .CK(clk), .Q(
        \registers[274][6] ) );
  EDFFX1 \registers_reg[274][5]  ( .D(n8313), .E(n596), .CK(clk), .Q(
        \registers[274][5] ) );
  EDFFX1 \registers_reg[274][4]  ( .D(n8255), .E(n596), .CK(clk), .Q(
        \registers[274][4] ) );
  EDFFX1 \registers_reg[274][3]  ( .D(n8200), .E(n596), .CK(clk), .Q(
        \registers[274][3] ) );
  EDFFX1 \registers_reg[274][2]  ( .D(n8160), .E(n596), .CK(clk), .Q(
        \registers[274][2] ) );
  EDFFX1 \registers_reg[274][1]  ( .D(n8104), .E(n596), .CK(clk), .Q(
        \registers[274][1] ) );
  EDFFX1 \registers_reg[274][0]  ( .D(n8044), .E(n596), .CK(clk), .Q(
        \registers[274][0] ) );
  EDFFX1 \registers_reg[270][7]  ( .D(n8428), .E(n592), .CK(clk), .Q(
        \registers[270][7] ) );
  EDFFX1 \registers_reg[270][6]  ( .D(n8370), .E(n592), .CK(clk), .Q(
        \registers[270][6] ) );
  EDFFX1 \registers_reg[270][5]  ( .D(n8312), .E(n592), .CK(clk), .Q(
        \registers[270][5] ) );
  EDFFX1 \registers_reg[270][4]  ( .D(n8254), .E(n592), .CK(clk), .Q(
        \registers[270][4] ) );
  EDFFX1 \registers_reg[270][3]  ( .D(n8201), .E(n592), .CK(clk), .Q(
        \registers[270][3] ) );
  EDFFX1 \registers_reg[270][2]  ( .D(n8155), .E(n592), .CK(clk), .Q(
        \registers[270][2] ) );
  EDFFX1 \registers_reg[270][1]  ( .D(n8099), .E(n592), .CK(clk), .Q(
        \registers[270][1] ) );
  EDFFX1 \registers_reg[270][0]  ( .D(n8045), .E(n592), .CK(clk), .Q(
        \registers[270][0] ) );
  EDFFX1 \registers_reg[266][7]  ( .D(n8428), .E(n588), .CK(clk), .Q(
        \registers[266][7] ) );
  EDFFX1 \registers_reg[266][6]  ( .D(n8370), .E(n588), .CK(clk), .Q(
        \registers[266][6] ) );
  EDFFX1 \registers_reg[266][5]  ( .D(n8312), .E(n588), .CK(clk), .Q(
        \registers[266][5] ) );
  EDFFX1 \registers_reg[266][4]  ( .D(n8254), .E(n588), .CK(clk), .Q(
        \registers[266][4] ) );
  EDFFX1 \registers_reg[266][3]  ( .D(n8202), .E(n588), .CK(clk), .Q(
        \registers[266][3] ) );
  EDFFX1 \registers_reg[266][2]  ( .D(n8156), .E(n588), .CK(clk), .Q(
        \registers[266][2] ) );
  EDFFX1 \registers_reg[266][1]  ( .D(n8100), .E(n588), .CK(clk), .Q(
        \registers[266][1] ) );
  EDFFX1 \registers_reg[266][0]  ( .D(n8040), .E(n588), .CK(clk), .Q(
        \registers[266][0] ) );
  EDFFX1 \registers_reg[262][7]  ( .D(n8429), .E(n972), .CK(clk), .Q(
        \registers[262][7] ) );
  EDFFX1 \registers_reg[262][6]  ( .D(n8371), .E(n972), .CK(clk), .Q(
        \registers[262][6] ) );
  EDFFX1 \registers_reg[262][5]  ( .D(n8313), .E(n972), .CK(clk), .Q(
        \registers[262][5] ) );
  EDFFX1 \registers_reg[262][4]  ( .D(n8255), .E(n972), .CK(clk), .Q(
        \registers[262][4] ) );
  EDFFX1 \registers_reg[262][3]  ( .D(n8200), .E(n972), .CK(clk), .Q(
        \registers[262][3] ) );
  EDFFX1 \registers_reg[262][2]  ( .D(n8157), .E(n972), .CK(clk), .Q(
        \registers[262][2] ) );
  EDFFX1 \registers_reg[262][1]  ( .D(n8101), .E(n972), .CK(clk), .Q(
        \registers[262][1] ) );
  EDFFX1 \registers_reg[262][0]  ( .D(n8041), .E(n972), .CK(clk), .Q(
        \registers[262][0] ) );
  EDFFX1 \registers_reg[258][7]  ( .D(n8429), .E(n968), .CK(clk), .Q(
        \registers[258][7] ) );
  EDFFX1 \registers_reg[258][6]  ( .D(n8371), .E(n968), .CK(clk), .Q(
        \registers[258][6] ) );
  EDFFX1 \registers_reg[258][5]  ( .D(n8313), .E(n968), .CK(clk), .Q(
        \registers[258][5] ) );
  EDFFX1 \registers_reg[258][4]  ( .D(n8255), .E(n968), .CK(clk), .Q(
        \registers[258][4] ) );
  EDFFX1 \registers_reg[258][3]  ( .D(n8201), .E(n968), .CK(clk), .Q(
        \registers[258][3] ) );
  EDFFX1 \registers_reg[258][2]  ( .D(n8155), .E(n968), .CK(clk), .Q(
        \registers[258][2] ) );
  EDFFX1 \registers_reg[258][1]  ( .D(n8099), .E(n968), .CK(clk), .Q(
        \registers[258][1] ) );
  EDFFX1 \registers_reg[258][0]  ( .D(n8042), .E(n968), .CK(clk), .Q(
        \registers[258][0] ) );
  EDFFX1 \registers_reg[254][7]  ( .D(n8410), .E(n584), .CK(clk), .Q(
        \registers[254][7] ) );
  EDFFX1 \registers_reg[254][6]  ( .D(n8352), .E(n584), .CK(clk), .Q(
        \registers[254][6] ) );
  EDFFX1 \registers_reg[254][5]  ( .D(n8294), .E(n584), .CK(clk), .Q(
        \registers[254][5] ) );
  EDFFX1 \registers_reg[254][4]  ( .D(n8236), .E(n584), .CK(clk), .Q(
        \registers[254][4] ) );
  EDFFX1 \registers_reg[254][3]  ( .D(n8190), .E(n584), .CK(clk), .Q(
        \registers[254][3] ) );
  EDFFX1 \registers_reg[254][2]  ( .D(n8142), .E(n584), .CK(clk), .Q(
        \registers[254][2] ) );
  EDFFX1 \registers_reg[254][1]  ( .D(n8086), .E(n584), .CK(clk), .Q(
        \registers[254][1] ) );
  EDFFX1 \registers_reg[254][0]  ( .D(n8025), .E(n584), .CK(clk), .Q(
        \registers[254][0] ) );
  EDFFX1 \registers_reg[250][7]  ( .D(n8411), .E(n580), .CK(clk), .Q(
        \registers[250][7] ) );
  EDFFX1 \registers_reg[250][6]  ( .D(n8353), .E(n580), .CK(clk), .Q(
        \registers[250][6] ) );
  EDFFX1 \registers_reg[250][5]  ( .D(n8295), .E(n580), .CK(clk), .Q(
        \registers[250][5] ) );
  EDFFX1 \registers_reg[250][4]  ( .D(n8237), .E(n580), .CK(clk), .Q(
        \registers[250][4] ) );
  EDFFX1 \registers_reg[250][3]  ( .D(n8188), .E(n580), .CK(clk), .Q(
        \registers[250][3] ) );
  EDFFX1 \registers_reg[250][2]  ( .D(n8143), .E(n580), .CK(clk), .Q(
        \registers[250][2] ) );
  EDFFX1 \registers_reg[250][1]  ( .D(n8087), .E(n580), .CK(clk), .Q(
        \registers[250][1] ) );
  EDFFX1 \registers_reg[250][0]  ( .D(n8026), .E(n580), .CK(clk), .Q(
        \registers[250][0] ) );
  EDFFX1 \registers_reg[246][7]  ( .D(n8412), .E(n576), .CK(clk), .Q(
        \registers[246][7] ) );
  EDFFX1 \registers_reg[246][6]  ( .D(n8354), .E(n576), .CK(clk), .Q(
        \registers[246][6] ) );
  EDFFX1 \registers_reg[246][5]  ( .D(n8296), .E(n576), .CK(clk), .Q(
        \registers[246][5] ) );
  EDFFX1 \registers_reg[246][4]  ( .D(n8238), .E(n576), .CK(clk), .Q(
        \registers[246][4] ) );
  EDFFX1 \registers_reg[246][3]  ( .D(n8189), .E(n576), .CK(clk), .Q(
        \registers[246][3] ) );
  EDFFX1 \registers_reg[246][2]  ( .D(n8141), .E(n576), .CK(clk), .Q(
        \registers[246][2] ) );
  EDFFX1 \registers_reg[246][1]  ( .D(n8085), .E(n576), .CK(clk), .Q(
        \registers[246][1] ) );
  EDFFX1 \registers_reg[246][0]  ( .D(n8027), .E(n576), .CK(clk), .Q(
        \registers[246][0] ) );
  EDFFX1 \registers_reg[242][7]  ( .D(n8410), .E(n572), .CK(clk), .Q(
        \registers[242][7] ) );
  EDFFX1 \registers_reg[242][6]  ( .D(n8352), .E(n572), .CK(clk), .Q(
        \registers[242][6] ) );
  EDFFX1 \registers_reg[242][5]  ( .D(n8294), .E(n572), .CK(clk), .Q(
        \registers[242][5] ) );
  EDFFX1 \registers_reg[242][4]  ( .D(n8236), .E(n572), .CK(clk), .Q(
        \registers[242][4] ) );
  EDFFX1 \registers_reg[242][3]  ( .D(n8190), .E(n572), .CK(clk), .Q(
        \registers[242][3] ) );
  EDFFX1 \registers_reg[242][2]  ( .D(n8142), .E(n572), .CK(clk), .Q(
        \registers[242][2] ) );
  EDFFX1 \registers_reg[242][1]  ( .D(n8086), .E(n572), .CK(clk), .Q(
        \registers[242][1] ) );
  EDFFX1 \registers_reg[242][0]  ( .D(n8025), .E(n572), .CK(clk), .Q(
        \registers[242][0] ) );
  EDFFX1 \registers_reg[238][7]  ( .D(n8411), .E(n568), .CK(clk), .Q(
        \registers[238][7] ) );
  EDFFX1 \registers_reg[238][6]  ( .D(n8353), .E(n568), .CK(clk), .Q(
        \registers[238][6] ) );
  EDFFX1 \registers_reg[238][5]  ( .D(n8295), .E(n568), .CK(clk), .Q(
        \registers[238][5] ) );
  EDFFX1 \registers_reg[238][4]  ( .D(n8237), .E(n568), .CK(clk), .Q(
        \registers[238][4] ) );
  EDFFX1 \registers_reg[238][3]  ( .D(n8188), .E(n568), .CK(clk), .Q(
        \registers[238][3] ) );
  EDFFX1 \registers_reg[238][2]  ( .D(n8143), .E(n568), .CK(clk), .Q(
        \registers[238][2] ) );
  EDFFX1 \registers_reg[238][1]  ( .D(n8087), .E(n568), .CK(clk), .Q(
        \registers[238][1] ) );
  EDFFX1 \registers_reg[238][0]  ( .D(n8026), .E(n568), .CK(clk), .Q(
        \registers[238][0] ) );
  EDFFX1 \registers_reg[234][7]  ( .D(n8412), .E(n564), .CK(clk), .Q(
        \registers[234][7] ) );
  EDFFX1 \registers_reg[234][6]  ( .D(n8354), .E(n564), .CK(clk), .Q(
        \registers[234][6] ) );
  EDFFX1 \registers_reg[234][5]  ( .D(n8296), .E(n564), .CK(clk), .Q(
        \registers[234][5] ) );
  EDFFX1 \registers_reg[234][4]  ( .D(n8238), .E(n564), .CK(clk), .Q(
        \registers[234][4] ) );
  EDFFX1 \registers_reg[234][3]  ( .D(n8186), .E(n564), .CK(clk), .Q(
        \registers[234][3] ) );
  EDFFX1 \registers_reg[234][2]  ( .D(n8141), .E(n564), .CK(clk), .Q(
        \registers[234][2] ) );
  EDFFX1 \registers_reg[234][1]  ( .D(n8085), .E(n564), .CK(clk), .Q(
        \registers[234][1] ) );
  EDFFX1 \registers_reg[234][0]  ( .D(n8027), .E(n564), .CK(clk), .Q(
        \registers[234][0] ) );
  EDFFX1 \registers_reg[230][7]  ( .D(n8410), .E(n1032), .CK(clk), .Q(
        \registers[230][7] ) );
  EDFFX1 \registers_reg[230][6]  ( .D(n8352), .E(n1032), .CK(clk), .Q(
        \registers[230][6] ) );
  EDFFX1 \registers_reg[230][5]  ( .D(n8294), .E(n1032), .CK(clk), .Q(
        \registers[230][5] ) );
  EDFFX1 \registers_reg[230][4]  ( .D(n8236), .E(n1032), .CK(clk), .Q(
        \registers[230][4] ) );
  EDFFX1 \registers_reg[230][3]  ( .D(n8187), .E(n1032), .CK(clk), .Q(
        \registers[230][3] ) );
  EDFFX1 \registers_reg[230][2]  ( .D(n8142), .E(n1032), .CK(clk), .Q(
        \registers[230][2] ) );
  EDFFX1 \registers_reg[230][1]  ( .D(n8086), .E(n1032), .CK(clk), .Q(
        \registers[230][1] ) );
  EDFFX1 \registers_reg[230][0]  ( .D(n8025), .E(n1032), .CK(clk), .Q(
        \registers[230][0] ) );
  EDFFX1 \registers_reg[226][7]  ( .D(n8411), .E(n965), .CK(clk), .Q(
        \registers[226][7] ) );
  EDFFX1 \registers_reg[226][6]  ( .D(n8353), .E(n965), .CK(clk), .Q(
        \registers[226][6] ) );
  EDFFX1 \registers_reg[226][5]  ( .D(n8295), .E(n965), .CK(clk), .Q(
        \registers[226][5] ) );
  EDFFX1 \registers_reg[226][4]  ( .D(n8237), .E(n965), .CK(clk), .Q(
        \registers[226][4] ) );
  EDFFX1 \registers_reg[226][3]  ( .D(n8185), .E(n965), .CK(clk), .Q(
        \registers[226][3] ) );
  EDFFX1 \registers_reg[226][2]  ( .D(n8143), .E(n965), .CK(clk), .Q(
        \registers[226][2] ) );
  EDFFX1 \registers_reg[226][1]  ( .D(n8087), .E(n965), .CK(clk), .Q(
        \registers[226][1] ) );
  EDFFX1 \registers_reg[226][0]  ( .D(n8026), .E(n965), .CK(clk), .Q(
        \registers[226][0] ) );
  EDFFX1 \registers_reg[222][7]  ( .D(n8412), .E(n560), .CK(clk), .Q(
        \registers[222][7] ) );
  EDFFX1 \registers_reg[222][6]  ( .D(n8354), .E(n560), .CK(clk), .Q(
        \registers[222][6] ) );
  EDFFX1 \registers_reg[222][5]  ( .D(n8296), .E(n560), .CK(clk), .Q(
        \registers[222][5] ) );
  EDFFX1 \registers_reg[222][4]  ( .D(n8238), .E(n560), .CK(clk), .Q(
        \registers[222][4] ) );
  EDFFX1 \registers_reg[222][3]  ( .D(n8186), .E(n560), .CK(clk), .Q(
        \registers[222][3] ) );
  EDFFX1 \registers_reg[222][2]  ( .D(n8141), .E(n560), .CK(clk), .Q(
        \registers[222][2] ) );
  EDFFX1 \registers_reg[222][1]  ( .D(n8085), .E(n560), .CK(clk), .Q(
        \registers[222][1] ) );
  EDFFX1 \registers_reg[222][0]  ( .D(n8027), .E(n560), .CK(clk), .Q(
        \registers[222][0] ) );
  EDFFX1 \registers_reg[218][7]  ( .D(n8410), .E(n556), .CK(clk), .Q(
        \registers[218][7] ) );
  EDFFX1 \registers_reg[218][6]  ( .D(n8352), .E(n556), .CK(clk), .Q(
        \registers[218][6] ) );
  EDFFX1 \registers_reg[218][5]  ( .D(n8294), .E(n556), .CK(clk), .Q(
        \registers[218][5] ) );
  EDFFX1 \registers_reg[218][4]  ( .D(n8236), .E(n556), .CK(clk), .Q(
        \registers[218][4] ) );
  EDFFX1 \registers_reg[218][3]  ( .D(n8187), .E(n556), .CK(clk), .Q(
        \registers[218][3] ) );
  EDFFX1 \registers_reg[218][2]  ( .D(n8139), .E(n556), .CK(clk), .Q(
        \registers[218][2] ) );
  EDFFX1 \registers_reg[218][1]  ( .D(n8083), .E(n556), .CK(clk), .Q(
        \registers[218][1] ) );
  EDFFX1 \registers_reg[218][0]  ( .D(n8022), .E(n556), .CK(clk), .Q(
        \registers[218][0] ) );
  EDFFX1 \registers_reg[214][7]  ( .D(n8411), .E(n552), .CK(clk), .Q(
        \registers[214][7] ) );
  EDFFX1 \registers_reg[214][6]  ( .D(n8353), .E(n552), .CK(clk), .Q(
        \registers[214][6] ) );
  EDFFX1 \registers_reg[214][5]  ( .D(n8295), .E(n552), .CK(clk), .Q(
        \registers[214][5] ) );
  EDFFX1 \registers_reg[214][4]  ( .D(n8237), .E(n552), .CK(clk), .Q(
        \registers[214][4] ) );
  EDFFX1 \registers_reg[214][3]  ( .D(n8185), .E(n552), .CK(clk), .Q(
        \registers[214][3] ) );
  EDFFX1 \registers_reg[214][2]  ( .D(n8140), .E(n552), .CK(clk), .Q(
        \registers[214][2] ) );
  EDFFX1 \registers_reg[214][1]  ( .D(n8084), .E(n552), .CK(clk), .Q(
        \registers[214][1] ) );
  EDFFX1 \registers_reg[214][0]  ( .D(n8023), .E(n552), .CK(clk), .Q(
        \registers[214][0] ) );
  EDFFX1 \registers_reg[210][7]  ( .D(n8412), .E(n548), .CK(clk), .Q(
        \registers[210][7] ) );
  EDFFX1 \registers_reg[210][6]  ( .D(n8354), .E(n548), .CK(clk), .Q(
        \registers[210][6] ) );
  EDFFX1 \registers_reg[210][5]  ( .D(n8296), .E(n548), .CK(clk), .Q(
        \registers[210][5] ) );
  EDFFX1 \registers_reg[210][4]  ( .D(n8238), .E(n548), .CK(clk), .Q(
        \registers[210][4] ) );
  EDFFX1 \registers_reg[210][3]  ( .D(n8186), .E(n548), .CK(clk), .Q(
        \registers[210][3] ) );
  EDFFX1 \registers_reg[210][2]  ( .D(n8138), .E(n548), .CK(clk), .Q(
        \registers[210][2] ) );
  EDFFX1 \registers_reg[210][1]  ( .D(n8082), .E(n548), .CK(clk), .Q(
        \registers[210][1] ) );
  EDFFX1 \registers_reg[210][0]  ( .D(n8024), .E(n548), .CK(clk), .Q(
        \registers[210][0] ) );
  EDFFX1 \registers_reg[206][7]  ( .D(n8408), .E(n544), .CK(clk), .Q(
        \registers[206][7] ) );
  EDFFX1 \registers_reg[206][6]  ( .D(n8350), .E(n544), .CK(clk), .Q(
        \registers[206][6] ) );
  EDFFX1 \registers_reg[206][5]  ( .D(n8292), .E(n544), .CK(clk), .Q(
        \registers[206][5] ) );
  EDFFX1 \registers_reg[206][4]  ( .D(n8234), .E(n544), .CK(clk), .Q(
        \registers[206][4] ) );
  EDFFX1 \registers_reg[206][3]  ( .D(n8187), .E(n544), .CK(clk), .Q(
        \registers[206][3] ) );
  EDFFX1 \registers_reg[206][2]  ( .D(n8139), .E(n544), .CK(clk), .Q(
        \registers[206][2] ) );
  EDFFX1 \registers_reg[206][1]  ( .D(n8083), .E(n544), .CK(clk), .Q(
        \registers[206][1] ) );
  EDFFX1 \registers_reg[206][0]  ( .D(n8022), .E(n544), .CK(clk), .Q(
        \registers[206][0] ) );
  EDFFX1 \registers_reg[202][7]  ( .D(n8409), .E(n540), .CK(clk), .Q(
        \registers[202][7] ) );
  EDFFX1 \registers_reg[202][6]  ( .D(n8351), .E(n540), .CK(clk), .Q(
        \registers[202][6] ) );
  EDFFX1 \registers_reg[202][5]  ( .D(n8293), .E(n540), .CK(clk), .Q(
        \registers[202][5] ) );
  EDFFX1 \registers_reg[202][4]  ( .D(n8235), .E(n540), .CK(clk), .Q(
        \registers[202][4] ) );
  EDFFX1 \registers_reg[202][3]  ( .D(n8185), .E(n540), .CK(clk), .Q(
        \registers[202][3] ) );
  EDFFX1 \registers_reg[202][2]  ( .D(n8140), .E(n540), .CK(clk), .Q(
        \registers[202][2] ) );
  EDFFX1 \registers_reg[202][1]  ( .D(n8084), .E(n540), .CK(clk), .Q(
        \registers[202][1] ) );
  EDFFX1 \registers_reg[202][0]  ( .D(n8023), .E(n540), .CK(clk), .Q(
        \registers[202][0] ) );
  EDFFX1 \registers_reg[198][7]  ( .D(n8407), .E(n1028), .CK(clk), .Q(
        \registers[198][7] ) );
  EDFFX1 \registers_reg[198][6]  ( .D(n8349), .E(n1028), .CK(clk), .Q(
        \registers[198][6] ) );
  EDFFX1 \registers_reg[198][5]  ( .D(n8291), .E(n1028), .CK(clk), .Q(
        \registers[198][5] ) );
  EDFFX1 \registers_reg[198][4]  ( .D(n8233), .E(n1028), .CK(clk), .Q(
        \registers[198][4] ) );
  EDFFX1 \registers_reg[198][3]  ( .D(n8186), .E(n1028), .CK(clk), .Q(
        \registers[198][3] ) );
  EDFFX1 \registers_reg[198][2]  ( .D(n8138), .E(n1028), .CK(clk), .Q(
        \registers[198][2] ) );
  EDFFX1 \registers_reg[198][1]  ( .D(n8082), .E(n1028), .CK(clk), .Q(
        \registers[198][1] ) );
  EDFFX1 \registers_reg[198][0]  ( .D(n8024), .E(n1028), .CK(clk), .Q(
        \registers[198][0] ) );
  EDFFX1 \registers_reg[194][7]  ( .D(n8408), .E(n962), .CK(clk), .Q(
        \registers[194][7] ) );
  EDFFX1 \registers_reg[194][6]  ( .D(n8350), .E(n962), .CK(clk), .Q(
        \registers[194][6] ) );
  EDFFX1 \registers_reg[194][5]  ( .D(n8292), .E(n962), .CK(clk), .Q(
        \registers[194][5] ) );
  EDFFX1 \registers_reg[194][4]  ( .D(n8234), .E(n962), .CK(clk), .Q(
        \registers[194][4] ) );
  EDFFX1 \registers_reg[194][3]  ( .D(n8187), .E(n962), .CK(clk), .Q(
        \registers[194][3] ) );
  EDFFX1 \registers_reg[194][2]  ( .D(n8139), .E(n962), .CK(clk), .Q(
        \registers[194][2] ) );
  EDFFX1 \registers_reg[194][1]  ( .D(n8083), .E(n962), .CK(clk), .Q(
        \registers[194][1] ) );
  EDFFX1 \registers_reg[194][0]  ( .D(n8022), .E(n962), .CK(clk), .Q(
        \registers[194][0] ) );
  EDFFX1 \registers_reg[190][7]  ( .D(n8407), .E(n536), .CK(clk), .Q(
        \registers[190][7] ) );
  EDFFX1 \registers_reg[190][6]  ( .D(n8349), .E(n536), .CK(clk), .Q(
        \registers[190][6] ) );
  EDFFX1 \registers_reg[190][5]  ( .D(n8291), .E(n536), .CK(clk), .Q(
        \registers[190][5] ) );
  EDFFX1 \registers_reg[190][4]  ( .D(n8233), .E(n536), .CK(clk), .Q(
        \registers[190][4] ) );
  EDFFX1 \registers_reg[190][3]  ( .D(n8186), .E(n536), .CK(clk), .Q(
        \registers[190][3] ) );
  EDFFX1 \registers_reg[190][2]  ( .D(n8138), .E(n536), .CK(clk), .Q(
        \registers[190][2] ) );
  EDFFX1 \registers_reg[190][1]  ( .D(n8082), .E(n536), .CK(clk), .Q(
        \registers[190][1] ) );
  EDFFX1 \registers_reg[190][0]  ( .D(n8024), .E(n536), .CK(clk), .Q(
        \registers[190][0] ) );
  EDFFX1 \registers_reg[186][7]  ( .D(n8408), .E(n532), .CK(clk), .Q(
        \registers[186][7] ) );
  EDFFX1 \registers_reg[186][6]  ( .D(n8350), .E(n532), .CK(clk), .Q(
        \registers[186][6] ) );
  EDFFX1 \registers_reg[186][5]  ( .D(n8292), .E(n532), .CK(clk), .Q(
        \registers[186][5] ) );
  EDFFX1 \registers_reg[186][4]  ( .D(n8234), .E(n532), .CK(clk), .Q(
        \registers[186][4] ) );
  EDFFX1 \registers_reg[186][3]  ( .D(n8187), .E(n532), .CK(clk), .Q(
        \registers[186][3] ) );
  EDFFX1 \registers_reg[186][2]  ( .D(n8139), .E(n532), .CK(clk), .Q(
        \registers[186][2] ) );
  EDFFX1 \registers_reg[186][1]  ( .D(n8083), .E(n532), .CK(clk), .Q(
        \registers[186][1] ) );
  EDFFX1 \registers_reg[186][0]  ( .D(n8022), .E(n532), .CK(clk), .Q(
        \registers[186][0] ) );
  EDFFX1 \registers_reg[182][7]  ( .D(n8409), .E(n528), .CK(clk), .Q(
        \registers[182][7] ) );
  EDFFX1 \registers_reg[182][6]  ( .D(n8351), .E(n528), .CK(clk), .Q(
        \registers[182][6] ) );
  EDFFX1 \registers_reg[182][5]  ( .D(n8293), .E(n528), .CK(clk), .Q(
        \registers[182][5] ) );
  EDFFX1 \registers_reg[182][4]  ( .D(n8235), .E(n528), .CK(clk), .Q(
        \registers[182][4] ) );
  EDFFX1 \registers_reg[182][3]  ( .D(n8185), .E(n528), .CK(clk), .Q(
        \registers[182][3] ) );
  EDFFX1 \registers_reg[182][2]  ( .D(n8140), .E(n528), .CK(clk), .Q(
        \registers[182][2] ) );
  EDFFX1 \registers_reg[182][1]  ( .D(n8084), .E(n528), .CK(clk), .Q(
        \registers[182][1] ) );
  EDFFX1 \registers_reg[182][0]  ( .D(n8023), .E(n528), .CK(clk), .Q(
        \registers[182][0] ) );
  EDFFX1 \registers_reg[178][7]  ( .D(n8407), .E(n524), .CK(clk), .Q(
        \registers[178][7] ) );
  EDFFX1 \registers_reg[178][6]  ( .D(n8349), .E(n524), .CK(clk), .Q(
        \registers[178][6] ) );
  EDFFX1 \registers_reg[178][5]  ( .D(n8291), .E(n524), .CK(clk), .Q(
        \registers[178][5] ) );
  EDFFX1 \registers_reg[178][4]  ( .D(n8233), .E(n524), .CK(clk), .Q(
        \registers[178][4] ) );
  EDFFX1 \registers_reg[178][3]  ( .D(n8186), .E(n524), .CK(clk), .Q(
        \registers[178][3] ) );
  EDFFX1 \registers_reg[178][2]  ( .D(n8138), .E(n524), .CK(clk), .Q(
        \registers[178][2] ) );
  EDFFX1 \registers_reg[178][1]  ( .D(n8082), .E(n524), .CK(clk), .Q(
        \registers[178][1] ) );
  EDFFX1 \registers_reg[178][0]  ( .D(n8024), .E(n524), .CK(clk), .Q(
        \registers[178][0] ) );
  EDFFX1 \registers_reg[174][7]  ( .D(n8408), .E(n520), .CK(clk), .Q(
        \registers[174][7] ) );
  EDFFX1 \registers_reg[174][6]  ( .D(n8350), .E(n520), .CK(clk), .Q(
        \registers[174][6] ) );
  EDFFX1 \registers_reg[174][5]  ( .D(n8292), .E(n520), .CK(clk), .Q(
        \registers[174][5] ) );
  EDFFX1 \registers_reg[174][4]  ( .D(n8234), .E(n520), .CK(clk), .Q(
        \registers[174][4] ) );
  EDFFX1 \registers_reg[174][3]  ( .D(n8187), .E(n520), .CK(clk), .Q(
        \registers[174][3] ) );
  EDFFX1 \registers_reg[174][2]  ( .D(n8139), .E(n520), .CK(clk), .Q(
        \registers[174][2] ) );
  EDFFX1 \registers_reg[174][1]  ( .D(n8083), .E(n520), .CK(clk), .Q(
        \registers[174][1] ) );
  EDFFX1 \registers_reg[174][0]  ( .D(n8022), .E(n520), .CK(clk), .Q(
        \registers[174][0] ) );
  EDFFX1 \registers_reg[170][7]  ( .D(n8409), .E(n516), .CK(clk), .Q(
        \registers[170][7] ) );
  EDFFX1 \registers_reg[170][6]  ( .D(n8351), .E(n516), .CK(clk), .Q(
        \registers[170][6] ) );
  EDFFX1 \registers_reg[170][5]  ( .D(n8293), .E(n516), .CK(clk), .Q(
        \registers[170][5] ) );
  EDFFX1 \registers_reg[170][4]  ( .D(n8235), .E(n516), .CK(clk), .Q(
        \registers[170][4] ) );
  EDFFX1 \registers_reg[170][3]  ( .D(n8182), .E(n516), .CK(clk), .Q(
        \registers[170][3] ) );
  EDFFX1 \registers_reg[170][2]  ( .D(n8140), .E(n516), .CK(clk), .Q(
        \registers[170][2] ) );
  EDFFX1 \registers_reg[170][1]  ( .D(n8084), .E(n516), .CK(clk), .Q(
        \registers[170][1] ) );
  EDFFX1 \registers_reg[170][0]  ( .D(n8023), .E(n516), .CK(clk), .Q(
        \registers[170][0] ) );
  EDFFX1 \registers_reg[166][7]  ( .D(n8407), .E(n1024), .CK(clk), .Q(
        \registers[166][7] ) );
  EDFFX1 \registers_reg[166][6]  ( .D(n8349), .E(n1024), .CK(clk), .Q(
        \registers[166][6] ) );
  EDFFX1 \registers_reg[166][5]  ( .D(n8291), .E(n1024), .CK(clk), .Q(
        \registers[166][5] ) );
  EDFFX1 \registers_reg[166][4]  ( .D(n8233), .E(n1024), .CK(clk), .Q(
        \registers[166][4] ) );
  EDFFX1 \registers_reg[166][3]  ( .D(n8183), .E(n1024), .CK(clk), .Q(
        \registers[166][3] ) );
  EDFFX1 \registers_reg[166][2]  ( .D(n8135), .E(n1024), .CK(clk), .Q(
        \registers[166][2] ) );
  EDFFX1 \registers_reg[166][1]  ( .D(n8079), .E(n1024), .CK(clk), .Q(
        \registers[166][1] ) );
  EDFFX1 \registers_reg[166][0]  ( .D(n8021), .E(n1024), .CK(clk), .Q(
        \registers[166][0] ) );
  EDFFX1 \registers_reg[162][7]  ( .D(n8408), .E(n959), .CK(clk), .Q(
        \registers[162][7] ) );
  EDFFX1 \registers_reg[162][6]  ( .D(n8350), .E(n959), .CK(clk), .Q(
        \registers[162][6] ) );
  EDFFX1 \registers_reg[162][5]  ( .D(n8292), .E(n959), .CK(clk), .Q(
        \registers[162][5] ) );
  EDFFX1 \registers_reg[162][4]  ( .D(n8234), .E(n959), .CK(clk), .Q(
        \registers[162][4] ) );
  EDFFX1 \registers_reg[162][3]  ( .D(n8184), .E(n959), .CK(clk), .Q(
        \registers[162][3] ) );
  EDFFX1 \registers_reg[162][2]  ( .D(n8136), .E(n959), .CK(clk), .Q(
        \registers[162][2] ) );
  EDFFX1 \registers_reg[162][1]  ( .D(n8080), .E(n959), .CK(clk), .Q(
        \registers[162][1] ) );
  EDFFX1 \registers_reg[162][0]  ( .D(n8019), .E(n959), .CK(clk), .Q(
        \registers[162][0] ) );
  EDFFX1 \registers_reg[158][7]  ( .D(n8404), .E(n512), .CK(clk), .Q(
        \registers[158][7] ) );
  EDFFX1 \registers_reg[158][6]  ( .D(n8346), .E(n512), .CK(clk), .Q(
        \registers[158][6] ) );
  EDFFX1 \registers_reg[158][5]  ( .D(n8288), .E(n512), .CK(clk), .Q(
        \registers[158][5] ) );
  EDFFX1 \registers_reg[158][4]  ( .D(n8230), .E(n512), .CK(clk), .Q(
        \registers[158][4] ) );
  EDFFX1 \registers_reg[158][3]  ( .D(n8182), .E(n512), .CK(clk), .Q(
        \registers[158][3] ) );
  EDFFX1 \registers_reg[158][2]  ( .D(n8137), .E(n512), .CK(clk), .Q(
        \registers[158][2] ) );
  EDFFX1 \registers_reg[158][1]  ( .D(n8081), .E(n512), .CK(clk), .Q(
        \registers[158][1] ) );
  EDFFX1 \registers_reg[158][0]  ( .D(n8020), .E(n512), .CK(clk), .Q(
        \registers[158][0] ) );
  EDFFX1 \registers_reg[154][7]  ( .D(n8405), .E(n508), .CK(clk), .Q(
        \registers[154][7] ) );
  EDFFX1 \registers_reg[154][6]  ( .D(n8347), .E(n508), .CK(clk), .Q(
        \registers[154][6] ) );
  EDFFX1 \registers_reg[154][5]  ( .D(n8289), .E(n508), .CK(clk), .Q(
        \registers[154][5] ) );
  EDFFX1 \registers_reg[154][4]  ( .D(n8231), .E(n508), .CK(clk), .Q(
        \registers[154][4] ) );
  EDFFX1 \registers_reg[154][3]  ( .D(n8183), .E(n508), .CK(clk), .Q(
        \registers[154][3] ) );
  EDFFX1 \registers_reg[154][2]  ( .D(n8135), .E(n508), .CK(clk), .Q(
        \registers[154][2] ) );
  EDFFX1 \registers_reg[154][1]  ( .D(n8079), .E(n508), .CK(clk), .Q(
        \registers[154][1] ) );
  EDFFX1 \registers_reg[154][0]  ( .D(n8021), .E(n508), .CK(clk), .Q(
        \registers[154][0] ) );
  EDFFX1 \registers_reg[150][7]  ( .D(n8406), .E(n504), .CK(clk), .Q(
        \registers[150][7] ) );
  EDFFX1 \registers_reg[150][6]  ( .D(n8348), .E(n504), .CK(clk), .Q(
        \registers[150][6] ) );
  EDFFX1 \registers_reg[150][5]  ( .D(n8290), .E(n504), .CK(clk), .Q(
        \registers[150][5] ) );
  EDFFX1 \registers_reg[150][4]  ( .D(n8232), .E(n504), .CK(clk), .Q(
        \registers[150][4] ) );
  EDFFX1 \registers_reg[150][3]  ( .D(n8184), .E(n504), .CK(clk), .Q(
        \registers[150][3] ) );
  EDFFX1 \registers_reg[150][2]  ( .D(n8136), .E(n504), .CK(clk), .Q(
        \registers[150][2] ) );
  EDFFX1 \registers_reg[150][1]  ( .D(n8080), .E(n504), .CK(clk), .Q(
        \registers[150][1] ) );
  EDFFX1 \registers_reg[150][0]  ( .D(n8019), .E(n504), .CK(clk), .Q(
        \registers[150][0] ) );
  EDFFX1 \registers_reg[146][7]  ( .D(n8404), .E(n500), .CK(clk), .Q(
        \registers[146][7] ) );
  EDFFX1 \registers_reg[146][6]  ( .D(n8346), .E(n500), .CK(clk), .Q(
        \registers[146][6] ) );
  EDFFX1 \registers_reg[146][5]  ( .D(n8288), .E(n500), .CK(clk), .Q(
        \registers[146][5] ) );
  EDFFX1 \registers_reg[146][4]  ( .D(n8230), .E(n500), .CK(clk), .Q(
        \registers[146][4] ) );
  EDFFX1 \registers_reg[146][3]  ( .D(n8182), .E(n500), .CK(clk), .Q(
        \registers[146][3] ) );
  EDFFX1 \registers_reg[146][2]  ( .D(n8137), .E(n500), .CK(clk), .Q(
        \registers[146][2] ) );
  EDFFX1 \registers_reg[146][1]  ( .D(n8081), .E(n500), .CK(clk), .Q(
        \registers[146][1] ) );
  EDFFX1 \registers_reg[146][0]  ( .D(n8020), .E(n500), .CK(clk), .Q(
        \registers[146][0] ) );
  EDFFX1 \registers_reg[142][7]  ( .D(n8405), .E(n496), .CK(clk), .Q(
        \registers[142][7] ) );
  EDFFX1 \registers_reg[142][6]  ( .D(n8347), .E(n496), .CK(clk), .Q(
        \registers[142][6] ) );
  EDFFX1 \registers_reg[142][5]  ( .D(n8289), .E(n496), .CK(clk), .Q(
        \registers[142][5] ) );
  EDFFX1 \registers_reg[142][4]  ( .D(n8231), .E(n496), .CK(clk), .Q(
        \registers[142][4] ) );
  EDFFX1 \registers_reg[142][3]  ( .D(n8183), .E(n496), .CK(clk), .Q(
        \registers[142][3] ) );
  EDFFX1 \registers_reg[142][2]  ( .D(n8135), .E(n496), .CK(clk), .Q(
        \registers[142][2] ) );
  EDFFX1 \registers_reg[142][1]  ( .D(n8079), .E(n496), .CK(clk), .Q(
        \registers[142][1] ) );
  EDFFX1 \registers_reg[142][0]  ( .D(n8021), .E(n496), .CK(clk), .Q(
        \registers[142][0] ) );
  EDFFX1 \registers_reg[138][7]  ( .D(n8406), .E(n492), .CK(clk), .Q(
        \registers[138][7] ) );
  EDFFX1 \registers_reg[138][6]  ( .D(n8348), .E(n492), .CK(clk), .Q(
        \registers[138][6] ) );
  EDFFX1 \registers_reg[138][5]  ( .D(n8290), .E(n492), .CK(clk), .Q(
        \registers[138][5] ) );
  EDFFX1 \registers_reg[138][4]  ( .D(n8232), .E(n492), .CK(clk), .Q(
        \registers[138][4] ) );
  EDFFX1 \registers_reg[138][3]  ( .D(n8184), .E(n492), .CK(clk), .Q(
        \registers[138][3] ) );
  EDFFX1 \registers_reg[138][2]  ( .D(n8136), .E(n492), .CK(clk), .Q(
        \registers[138][2] ) );
  EDFFX1 \registers_reg[138][1]  ( .D(n8080), .E(n492), .CK(clk), .Q(
        \registers[138][1] ) );
  EDFFX1 \registers_reg[138][0]  ( .D(n8019), .E(n492), .CK(clk), .Q(
        \registers[138][0] ) );
  EDFFX1 \registers_reg[134][7]  ( .D(n8404), .E(n1020), .CK(clk), .Q(
        \registers[134][7] ) );
  EDFFX1 \registers_reg[134][6]  ( .D(n8346), .E(n1020), .CK(clk), .Q(
        \registers[134][6] ) );
  EDFFX1 \registers_reg[134][5]  ( .D(n8288), .E(n1020), .CK(clk), .Q(
        \registers[134][5] ) );
  EDFFX1 \registers_reg[134][4]  ( .D(n8230), .E(n1020), .CK(clk), .Q(
        \registers[134][4] ) );
  EDFFX1 \registers_reg[134][3]  ( .D(n8182), .E(n1020), .CK(clk), .Q(
        \registers[134][3] ) );
  EDFFX1 \registers_reg[134][2]  ( .D(n8137), .E(n1020), .CK(clk), .Q(
        \registers[134][2] ) );
  EDFFX1 \registers_reg[134][1]  ( .D(n8081), .E(n1020), .CK(clk), .Q(
        \registers[134][1] ) );
  EDFFX1 \registers_reg[134][0]  ( .D(n8020), .E(n1020), .CK(clk), .Q(
        \registers[134][0] ) );
  EDFFX1 \registers_reg[130][7]  ( .D(n8405), .E(n956), .CK(clk), .Q(
        \registers[130][7] ) );
  EDFFX1 \registers_reg[130][6]  ( .D(n8347), .E(n956), .CK(clk), .Q(
        \registers[130][6] ) );
  EDFFX1 \registers_reg[130][5]  ( .D(n8289), .E(n956), .CK(clk), .Q(
        \registers[130][5] ) );
  EDFFX1 \registers_reg[130][4]  ( .D(n8231), .E(n956), .CK(clk), .Q(
        \registers[130][4] ) );
  EDFFX1 \registers_reg[130][3]  ( .D(n8183), .E(n956), .CK(clk), .Q(
        \registers[130][3] ) );
  EDFFX1 \registers_reg[130][2]  ( .D(n8135), .E(n956), .CK(clk), .Q(
        \registers[130][2] ) );
  EDFFX1 \registers_reg[130][1]  ( .D(n8079), .E(n956), .CK(clk), .Q(
        \registers[130][1] ) );
  EDFFX1 \registers_reg[130][0]  ( .D(n8021), .E(n956), .CK(clk), .Q(
        \registers[130][0] ) );
  EDFFX1 \registers_reg[126][7]  ( .D(n8420), .E(n488), .CK(clk), .Q(
        \registers[126][7] ) );
  EDFFX1 \registers_reg[126][6]  ( .D(n8362), .E(n488), .CK(clk), .Q(
        \registers[126][6] ) );
  EDFFX1 \registers_reg[126][5]  ( .D(n8304), .E(n488), .CK(clk), .Q(
        \registers[126][5] ) );
  EDFFX1 \registers_reg[126][4]  ( .D(n8246), .E(n488), .CK(clk), .Q(
        \registers[126][4] ) );
  EDFFX1 \registers_reg[126][3]  ( .D(n8194), .E(n488), .CK(clk), .Q(
        \registers[126][3] ) );
  EDFFX1 \registers_reg[126][2]  ( .D(n8728), .E(n488), .CK(clk), .Q(
        \registers[126][2] ) );
  EDFFX1 \registers_reg[126][1]  ( .D(n8700), .E(n488), .CK(clk), .Q(
        \registers[126][1] ) );
  EDFFX1 \registers_reg[126][0]  ( .D(n8036), .E(n488), .CK(clk), .Q(
        \registers[126][0] ) );
  EDFFX1 \registers_reg[122][7]  ( .D(n8421), .E(n484), .CK(clk), .Q(
        \registers[122][7] ) );
  EDFFX1 \registers_reg[122][6]  ( .D(n8363), .E(n484), .CK(clk), .Q(
        \registers[122][6] ) );
  EDFFX1 \registers_reg[122][5]  ( .D(n8305), .E(n484), .CK(clk), .Q(
        \registers[122][5] ) );
  EDFFX1 \registers_reg[122][4]  ( .D(n8247), .E(n484), .CK(clk), .Q(
        \registers[122][4] ) );
  EDFFX1 \registers_reg[122][3]  ( .D(n8195), .E(n484), .CK(clk), .Q(
        \registers[122][3] ) );
  EDFFX1 \registers_reg[122][2]  ( .D(n8150), .E(n484), .CK(clk), .Q(
        \registers[122][2] ) );
  EDFFX1 \registers_reg[122][1]  ( .D(n8094), .E(n484), .CK(clk), .Q(
        \registers[122][1] ) );
  EDFFX1 \registers_reg[122][0]  ( .D(n8034), .E(n484), .CK(clk), .Q(
        \registers[122][0] ) );
  EDFFX1 \registers_reg[118][7]  ( .D(n8419), .E(n480), .CK(clk), .Q(
        \registers[118][7] ) );
  EDFFX1 \registers_reg[118][6]  ( .D(n8361), .E(n480), .CK(clk), .Q(
        \registers[118][6] ) );
  EDFFX1 \registers_reg[118][5]  ( .D(n8303), .E(n480), .CK(clk), .Q(
        \registers[118][5] ) );
  EDFFX1 \registers_reg[118][4]  ( .D(n8245), .E(n480), .CK(clk), .Q(
        \registers[118][4] ) );
  EDFFX1 \registers_reg[118][3]  ( .D(n8196), .E(n480), .CK(clk), .Q(
        \registers[118][3] ) );
  EDFFX1 \registers_reg[118][2]  ( .D(n8151), .E(n480), .CK(clk), .Q(
        \registers[118][2] ) );
  EDFFX1 \registers_reg[118][1]  ( .D(n8095), .E(n480), .CK(clk), .Q(
        \registers[118][1] ) );
  EDFFX1 \registers_reg[118][0]  ( .D(n8035), .E(n480), .CK(clk), .Q(
        \registers[118][0] ) );
  EDFFX1 \registers_reg[114][7]  ( .D(n8420), .E(n476), .CK(clk), .Q(
        \registers[114][7] ) );
  EDFFX1 \registers_reg[114][6]  ( .D(n8362), .E(n476), .CK(clk), .Q(
        \registers[114][6] ) );
  EDFFX1 \registers_reg[114][5]  ( .D(n8304), .E(n476), .CK(clk), .Q(
        \registers[114][5] ) );
  EDFFX1 \registers_reg[114][4]  ( .D(n8246), .E(n476), .CK(clk), .Q(
        \registers[114][4] ) );
  EDFFX1 \registers_reg[114][3]  ( .D(n8194), .E(n476), .CK(clk), .Q(
        \registers[114][3] ) );
  EDFFX1 \registers_reg[114][2]  ( .D(n8149), .E(n476), .CK(clk), .Q(
        \registers[114][2] ) );
  EDFFX1 \registers_reg[114][1]  ( .D(n8093), .E(n476), .CK(clk), .Q(
        \registers[114][1] ) );
  EDFFX1 \registers_reg[114][0]  ( .D(n8033), .E(n476), .CK(clk), .Q(
        \registers[114][0] ) );
  EDFFX1 \registers_reg[110][7]  ( .D(n8421), .E(n472), .CK(clk), .Q(
        \registers[110][7] ) );
  EDFFX1 \registers_reg[110][6]  ( .D(n8363), .E(n472), .CK(clk), .Q(
        \registers[110][6] ) );
  EDFFX1 \registers_reg[110][5]  ( .D(n8305), .E(n472), .CK(clk), .Q(
        \registers[110][5] ) );
  EDFFX1 \registers_reg[110][4]  ( .D(n8247), .E(n472), .CK(clk), .Q(
        \registers[110][4] ) );
  EDFFX1 \registers_reg[110][3]  ( .D(n8195), .E(n472), .CK(clk), .Q(
        \registers[110][3] ) );
  EDFFX1 \registers_reg[110][2]  ( .D(n8147), .E(n472), .CK(clk), .Q(
        \registers[110][2] ) );
  EDFFX1 \registers_reg[110][1]  ( .D(n8091), .E(n472), .CK(clk), .Q(
        \registers[110][1] ) );
  EDFFX1 \registers_reg[110][0]  ( .D(n8031), .E(n472), .CK(clk), .Q(
        \registers[110][0] ) );
  EDFFX1 \registers_reg[106][7]  ( .D(n8419), .E(n468), .CK(clk), .Q(
        \registers[106][7] ) );
  EDFFX1 \registers_reg[106][6]  ( .D(n8361), .E(n468), .CK(clk), .Q(
        \registers[106][6] ) );
  EDFFX1 \registers_reg[106][5]  ( .D(n8303), .E(n468), .CK(clk), .Q(
        \registers[106][5] ) );
  EDFFX1 \registers_reg[106][4]  ( .D(n8245), .E(n468), .CK(clk), .Q(
        \registers[106][4] ) );
  EDFFX1 \registers_reg[106][3]  ( .D(n8196), .E(n468), .CK(clk), .Q(
        \registers[106][3] ) );
  EDFFX1 \registers_reg[106][2]  ( .D(n8148), .E(n468), .CK(clk), .Q(
        \registers[106][2] ) );
  EDFFX1 \registers_reg[106][1]  ( .D(n8092), .E(n468), .CK(clk), .Q(
        \registers[106][1] ) );
  EDFFX1 \registers_reg[106][0]  ( .D(n8032), .E(n468), .CK(clk), .Q(
        \registers[106][0] ) );
  EDFFX1 \registers_reg[102][7]  ( .D(n8420), .E(n953), .CK(clk), .Q(
        \registers[102][7] ) );
  EDFFX1 \registers_reg[102][6]  ( .D(n8362), .E(n953), .CK(clk), .Q(
        \registers[102][6] ) );
  EDFFX1 \registers_reg[102][5]  ( .D(n8304), .E(n953), .CK(clk), .Q(
        \registers[102][5] ) );
  EDFFX1 \registers_reg[102][4]  ( .D(n8246), .E(n953), .CK(clk), .Q(
        \registers[102][4] ) );
  EDFFX1 \registers_reg[102][3]  ( .D(n8191), .E(n953), .CK(clk), .Q(
        \registers[102][3] ) );
  EDFFX1 \registers_reg[102][2]  ( .D(n8149), .E(n953), .CK(clk), .Q(
        \registers[102][2] ) );
  EDFFX1 \registers_reg[102][1]  ( .D(n8093), .E(n953), .CK(clk), .Q(
        \registers[102][1] ) );
  EDFFX1 \registers_reg[102][0]  ( .D(n8033), .E(n953), .CK(clk), .Q(
        \registers[102][0] ) );
  EDFFX1 \registers_reg[98][7]  ( .D(n8416), .E(n949), .CK(clk), .Q(
        \registers[98][7] ) );
  EDFFX1 \registers_reg[98][6]  ( .D(n8358), .E(n949), .CK(clk), .Q(
        \registers[98][6] ) );
  EDFFX1 \registers_reg[98][5]  ( .D(n8300), .E(n949), .CK(clk), .Q(
        \registers[98][5] ) );
  EDFFX1 \registers_reg[98][4]  ( .D(n8242), .E(n949), .CK(clk), .Q(
        \registers[98][4] ) );
  EDFFX1 \registers_reg[98][3]  ( .D(n8192), .E(n949), .CK(clk), .Q(
        \registers[98][3] ) );
  EDFFX1 \registers_reg[98][2]  ( .D(n8147), .E(n949), .CK(clk), .Q(
        \registers[98][2] ) );
  EDFFX1 \registers_reg[98][1]  ( .D(n8091), .E(n949), .CK(clk), .Q(
        \registers[98][1] ) );
  EDFFX1 \registers_reg[98][0]  ( .D(n8031), .E(n949), .CK(clk), .Q(
        \registers[98][0] ) );
  EDFFX1 \registers_reg[94][7]  ( .D(n8417), .E(n464), .CK(clk), .Q(
        \registers[94][7] ) );
  EDFFX1 \registers_reg[94][6]  ( .D(n8359), .E(n464), .CK(clk), .Q(
        \registers[94][6] ) );
  EDFFX1 \registers_reg[94][5]  ( .D(n8301), .E(n464), .CK(clk), .Q(
        \registers[94][5] ) );
  EDFFX1 \registers_reg[94][4]  ( .D(n8243), .E(n464), .CK(clk), .Q(
        \registers[94][4] ) );
  EDFFX1 \registers_reg[94][3]  ( .D(n8193), .E(n464), .CK(clk), .Q(
        \registers[94][3] ) );
  EDFFX1 \registers_reg[94][2]  ( .D(n8148), .E(n464), .CK(clk), .Q(
        \registers[94][2] ) );
  EDFFX1 \registers_reg[94][1]  ( .D(n8092), .E(n464), .CK(clk), .Q(
        \registers[94][1] ) );
  EDFFX1 \registers_reg[94][0]  ( .D(n8032), .E(n464), .CK(clk), .Q(
        \registers[94][0] ) );
  EDFFX1 \registers_reg[90][7]  ( .D(n8418), .E(n460), .CK(clk), .Q(
        \registers[90][7] ) );
  EDFFX1 \registers_reg[90][6]  ( .D(n8360), .E(n460), .CK(clk), .Q(
        \registers[90][6] ) );
  EDFFX1 \registers_reg[90][5]  ( .D(n8302), .E(n460), .CK(clk), .Q(
        \registers[90][5] ) );
  EDFFX1 \registers_reg[90][4]  ( .D(n8244), .E(n460), .CK(clk), .Q(
        \registers[90][4] ) );
  EDFFX1 \registers_reg[90][3]  ( .D(n8191), .E(n460), .CK(clk), .Q(
        \registers[90][3] ) );
  EDFFX1 \registers_reg[90][2]  ( .D(n8149), .E(n460), .CK(clk), .Q(
        \registers[90][2] ) );
  EDFFX1 \registers_reg[90][1]  ( .D(n8093), .E(n460), .CK(clk), .Q(
        \registers[90][1] ) );
  EDFFX1 \registers_reg[90][0]  ( .D(n8033), .E(n460), .CK(clk), .Q(
        \registers[90][0] ) );
  EDFFX1 \registers_reg[86][7]  ( .D(n8416), .E(n456), .CK(clk), .Q(
        \registers[86][7] ) );
  EDFFX1 \registers_reg[86][6]  ( .D(n8358), .E(n456), .CK(clk), .Q(
        \registers[86][6] ) );
  EDFFX1 \registers_reg[86][5]  ( .D(n8300), .E(n456), .CK(clk), .Q(
        \registers[86][5] ) );
  EDFFX1 \registers_reg[86][4]  ( .D(n8242), .E(n456), .CK(clk), .Q(
        \registers[86][4] ) );
  EDFFX1 \registers_reg[86][3]  ( .D(n8192), .E(n456), .CK(clk), .Q(
        \registers[86][3] ) );
  EDFFX1 \registers_reg[86][2]  ( .D(n8147), .E(n456), .CK(clk), .Q(
        \registers[86][2] ) );
  EDFFX1 \registers_reg[86][1]  ( .D(n8091), .E(n456), .CK(clk), .Q(
        \registers[86][1] ) );
  EDFFX1 \registers_reg[86][0]  ( .D(n8031), .E(n456), .CK(clk), .Q(
        \registers[86][0] ) );
  EDFFX1 \registers_reg[82][7]  ( .D(n8417), .E(n452), .CK(clk), .Q(
        \registers[82][7] ) );
  EDFFX1 \registers_reg[82][6]  ( .D(n8359), .E(n452), .CK(clk), .Q(
        \registers[82][6] ) );
  EDFFX1 \registers_reg[82][5]  ( .D(n8301), .E(n452), .CK(clk), .Q(
        \registers[82][5] ) );
  EDFFX1 \registers_reg[82][4]  ( .D(n8243), .E(n452), .CK(clk), .Q(
        \registers[82][4] ) );
  EDFFX1 \registers_reg[82][3]  ( .D(n8193), .E(n452), .CK(clk), .Q(
        \registers[82][3] ) );
  EDFFX1 \registers_reg[82][2]  ( .D(n8148), .E(n452), .CK(clk), .Q(
        \registers[82][2] ) );
  EDFFX1 \registers_reg[82][1]  ( .D(n8092), .E(n452), .CK(clk), .Q(
        \registers[82][1] ) );
  EDFFX1 \registers_reg[82][0]  ( .D(n8032), .E(n452), .CK(clk), .Q(
        \registers[82][0] ) );
  EDFFX1 \registers_reg[78][7]  ( .D(n8418), .E(n448), .CK(clk), .Q(
        \registers[78][7] ) );
  EDFFX1 \registers_reg[78][6]  ( .D(n8360), .E(n448), .CK(clk), .Q(
        \registers[78][6] ) );
  EDFFX1 \registers_reg[78][5]  ( .D(n8302), .E(n448), .CK(clk), .Q(
        \registers[78][5] ) );
  EDFFX1 \registers_reg[78][4]  ( .D(n8244), .E(n448), .CK(clk), .Q(
        \registers[78][4] ) );
  EDFFX1 \registers_reg[78][3]  ( .D(n8191), .E(n448), .CK(clk), .Q(
        \registers[78][3] ) );
  EDFFX1 \registers_reg[78][2]  ( .D(n8149), .E(n448), .CK(clk), .Q(
        \registers[78][2] ) );
  EDFFX1 \registers_reg[78][1]  ( .D(n8093), .E(n448), .CK(clk), .Q(
        \registers[78][1] ) );
  EDFFX1 \registers_reg[78][0]  ( .D(n8033), .E(n448), .CK(clk), .Q(
        \registers[78][0] ) );
  EDFFX1 \registers_reg[74][7]  ( .D(n8416), .E(n444), .CK(clk), .Q(
        \registers[74][7] ) );
  EDFFX1 \registers_reg[74][6]  ( .D(n8358), .E(n444), .CK(clk), .Q(
        \registers[74][6] ) );
  EDFFX1 \registers_reg[74][5]  ( .D(n8300), .E(n444), .CK(clk), .Q(
        \registers[74][5] ) );
  EDFFX1 \registers_reg[74][4]  ( .D(n8242), .E(n444), .CK(clk), .Q(
        \registers[74][4] ) );
  EDFFX1 \registers_reg[74][3]  ( .D(n8192), .E(n444), .CK(clk), .Q(
        \registers[74][3] ) );
  EDFFX1 \registers_reg[74][2]  ( .D(n8147), .E(n444), .CK(clk), .Q(
        \registers[74][2] ) );
  EDFFX1 \registers_reg[74][1]  ( .D(n8091), .E(n444), .CK(clk), .Q(
        \registers[74][1] ) );
  EDFFX1 \registers_reg[74][0]  ( .D(n8031), .E(n444), .CK(clk), .Q(
        \registers[74][0] ) );
  EDFFX1 \registers_reg[70][7]  ( .D(n8417), .E(n946), .CK(clk), .Q(
        \registers[70][7] ) );
  EDFFX1 \registers_reg[70][6]  ( .D(n8359), .E(n946), .CK(clk), .Q(
        \registers[70][6] ) );
  EDFFX1 \registers_reg[70][5]  ( .D(n8301), .E(n946), .CK(clk), .Q(
        \registers[70][5] ) );
  EDFFX1 \registers_reg[70][4]  ( .D(n8243), .E(n946), .CK(clk), .Q(
        \registers[70][4] ) );
  EDFFX1 \registers_reg[70][3]  ( .D(n8193), .E(n946), .CK(clk), .Q(
        \registers[70][3] ) );
  EDFFX1 \registers_reg[70][2]  ( .D(n8148), .E(n946), .CK(clk), .Q(
        \registers[70][2] ) );
  EDFFX1 \registers_reg[70][1]  ( .D(n8092), .E(n946), .CK(clk), .Q(
        \registers[70][1] ) );
  EDFFX1 \registers_reg[70][0]  ( .D(n8032), .E(n946), .CK(clk), .Q(
        \registers[70][0] ) );
  EDFFX1 \registers_reg[66][7]  ( .D(n8418), .E(n942), .CK(clk), .Q(
        \registers[66][7] ) );
  EDFFX1 \registers_reg[66][6]  ( .D(n8360), .E(n942), .CK(clk), .Q(
        \registers[66][6] ) );
  EDFFX1 \registers_reg[66][5]  ( .D(n8302), .E(n942), .CK(clk), .Q(
        \registers[66][5] ) );
  EDFFX1 \registers_reg[66][4]  ( .D(n8244), .E(n942), .CK(clk), .Q(
        \registers[66][4] ) );
  EDFFX1 \registers_reg[66][3]  ( .D(n8191), .E(n942), .CK(clk), .Q(
        \registers[66][3] ) );
  EDFFX1 \registers_reg[66][2]  ( .D(n8149), .E(n942), .CK(clk), .Q(
        \registers[66][2] ) );
  EDFFX1 \registers_reg[66][1]  ( .D(n8093), .E(n942), .CK(clk), .Q(
        \registers[66][1] ) );
  EDFFX1 \registers_reg[66][0]  ( .D(n8033), .E(n942), .CK(clk), .Q(
        \registers[66][0] ) );
  EDFFX1 \registers_reg[62][7]  ( .D(n8417), .E(n440), .CK(clk), .Q(
        \registers[62][7] ) );
  EDFFX1 \registers_reg[62][6]  ( .D(n8359), .E(n440), .CK(clk), .Q(
        \registers[62][6] ) );
  EDFFX1 \registers_reg[62][5]  ( .D(n8301), .E(n440), .CK(clk), .Q(
        \registers[62][5] ) );
  EDFFX1 \registers_reg[62][4]  ( .D(n8243), .E(n440), .CK(clk), .Q(
        \registers[62][4] ) );
  EDFFX1 \registers_reg[62][3]  ( .D(n8193), .E(n440), .CK(clk), .Q(
        \registers[62][3] ) );
  EDFFX1 \registers_reg[62][2]  ( .D(n8145), .E(n440), .CK(clk), .Q(
        \registers[62][2] ) );
  EDFFX1 \registers_reg[62][1]  ( .D(n8089), .E(n440), .CK(clk), .Q(
        \registers[62][1] ) );
  EDFFX1 \registers_reg[62][0]  ( .D(n8029), .E(n440), .CK(clk), .Q(
        \registers[62][0] ) );
  EDFFX1 \registers_reg[58][7]  ( .D(n8418), .E(n436), .CK(clk), .Q(
        \registers[58][7] ) );
  EDFFX1 \registers_reg[58][6]  ( .D(n8360), .E(n436), .CK(clk), .Q(
        \registers[58][6] ) );
  EDFFX1 \registers_reg[58][5]  ( .D(n8302), .E(n436), .CK(clk), .Q(
        \registers[58][5] ) );
  EDFFX1 \registers_reg[58][4]  ( .D(n8244), .E(n436), .CK(clk), .Q(
        \registers[58][4] ) );
  EDFFX1 \registers_reg[58][3]  ( .D(n8191), .E(n436), .CK(clk), .Q(
        \registers[58][3] ) );
  EDFFX1 \registers_reg[58][2]  ( .D(n8146), .E(n436), .CK(clk), .Q(
        \registers[58][2] ) );
  EDFFX1 \registers_reg[58][1]  ( .D(n8090), .E(n436), .CK(clk), .Q(
        \registers[58][1] ) );
  EDFFX1 \registers_reg[58][0]  ( .D(n8030), .E(n436), .CK(clk), .Q(
        \registers[58][0] ) );
  EDFFX1 \registers_reg[54][7]  ( .D(n8416), .E(n432), .CK(clk), .Q(
        \registers[54][7] ) );
  EDFFX1 \registers_reg[54][6]  ( .D(n8358), .E(n432), .CK(clk), .Q(
        \registers[54][6] ) );
  EDFFX1 \registers_reg[54][5]  ( .D(n8300), .E(n432), .CK(clk), .Q(
        \registers[54][5] ) );
  EDFFX1 \registers_reg[54][4]  ( .D(n8242), .E(n432), .CK(clk), .Q(
        \registers[54][4] ) );
  EDFFX1 \registers_reg[54][3]  ( .D(n8192), .E(n432), .CK(clk), .Q(
        \registers[54][3] ) );
  EDFFX1 \registers_reg[54][2]  ( .D(n8144), .E(n432), .CK(clk), .Q(
        \registers[54][2] ) );
  EDFFX1 \registers_reg[54][1]  ( .D(n8088), .E(n432), .CK(clk), .Q(
        \registers[54][1] ) );
  EDFFX1 \registers_reg[54][0]  ( .D(n8028), .E(n432), .CK(clk), .Q(
        \registers[54][0] ) );
  EDFFX1 \registers_reg[50][7]  ( .D(n8415), .E(n428), .CK(clk), .Q(
        \registers[50][7] ) );
  EDFFX1 \registers_reg[50][6]  ( .D(n8357), .E(n428), .CK(clk), .Q(
        \registers[50][6] ) );
  EDFFX1 \registers_reg[50][5]  ( .D(n8299), .E(n428), .CK(clk), .Q(
        \registers[50][5] ) );
  EDFFX1 \registers_reg[50][4]  ( .D(n8241), .E(n428), .CK(clk), .Q(
        \registers[50][4] ) );
  EDFFX1 \registers_reg[50][3]  ( .D(n8193), .E(n428), .CK(clk), .Q(
        \registers[50][3] ) );
  EDFFX1 \registers_reg[50][2]  ( .D(n8145), .E(n428), .CK(clk), .Q(
        \registers[50][2] ) );
  EDFFX1 \registers_reg[50][1]  ( .D(n8089), .E(n428), .CK(clk), .Q(
        \registers[50][1] ) );
  EDFFX1 \registers_reg[50][0]  ( .D(n8029), .E(n428), .CK(clk), .Q(
        \registers[50][0] ) );
  EDFFX1 \registers_reg[46][7]  ( .D(n8413), .E(n424), .CK(clk), .Q(
        \registers[46][7] ) );
  EDFFX1 \registers_reg[46][6]  ( .D(n8355), .E(n424), .CK(clk), .Q(
        \registers[46][6] ) );
  EDFFX1 \registers_reg[46][5]  ( .D(n8297), .E(n424), .CK(clk), .Q(
        \registers[46][5] ) );
  EDFFX1 \registers_reg[46][4]  ( .D(n8239), .E(n424), .CK(clk), .Q(
        \registers[46][4] ) );
  EDFFX1 \registers_reg[46][3]  ( .D(n8191), .E(n424), .CK(clk), .Q(
        \registers[46][3] ) );
  EDFFX1 \registers_reg[46][2]  ( .D(n8146), .E(n424), .CK(clk), .Q(
        \registers[46][2] ) );
  EDFFX1 \registers_reg[46][1]  ( .D(n8090), .E(n424), .CK(clk), .Q(
        \registers[46][1] ) );
  EDFFX1 \registers_reg[46][0]  ( .D(n8030), .E(n424), .CK(clk), .Q(
        \registers[46][0] ) );
  EDFFX1 \registers_reg[42][7]  ( .D(n8414), .E(n420), .CK(clk), .Q(
        \registers[42][7] ) );
  EDFFX1 \registers_reg[42][6]  ( .D(n8356), .E(n420), .CK(clk), .Q(
        \registers[42][6] ) );
  EDFFX1 \registers_reg[42][5]  ( .D(n8298), .E(n420), .CK(clk), .Q(
        \registers[42][5] ) );
  EDFFX1 \registers_reg[42][4]  ( .D(n8240), .E(n420), .CK(clk), .Q(
        \registers[42][4] ) );
  EDFFX1 \registers_reg[42][3]  ( .D(n8189), .E(n420), .CK(clk), .Q(
        \registers[42][3] ) );
  EDFFX1 \registers_reg[42][2]  ( .D(n8144), .E(n420), .CK(clk), .Q(
        \registers[42][2] ) );
  EDFFX1 \registers_reg[42][1]  ( .D(n8088), .E(n420), .CK(clk), .Q(
        \registers[42][1] ) );
  EDFFX1 \registers_reg[42][0]  ( .D(n8028), .E(n420), .CK(clk), .Q(
        \registers[42][0] ) );
  EDFFX1 \registers_reg[38][7]  ( .D(n8415), .E(n939), .CK(clk), .Q(
        \registers[38][7] ) );
  EDFFX1 \registers_reg[38][6]  ( .D(n8357), .E(n939), .CK(clk), .Q(
        \registers[38][6] ) );
  EDFFX1 \registers_reg[38][5]  ( .D(n8299), .E(n939), .CK(clk), .Q(
        \registers[38][5] ) );
  EDFFX1 \registers_reg[38][4]  ( .D(n8241), .E(n939), .CK(clk), .Q(
        \registers[38][4] ) );
  EDFFX1 \registers_reg[38][3]  ( .D(n8190), .E(n939), .CK(clk), .Q(
        \registers[38][3] ) );
  EDFFX1 \registers_reg[38][2]  ( .D(n8145), .E(n939), .CK(clk), .Q(
        \registers[38][2] ) );
  EDFFX1 \registers_reg[38][1]  ( .D(n8089), .E(n939), .CK(clk), .Q(
        \registers[38][1] ) );
  EDFFX1 \registers_reg[38][0]  ( .D(n8029), .E(n939), .CK(clk), .Q(
        \registers[38][0] ) );
  EDFFX1 \registers_reg[34][7]  ( .D(n8413), .E(n935), .CK(clk), .Q(
        \registers[34][7] ) );
  EDFFX1 \registers_reg[34][6]  ( .D(n8355), .E(n935), .CK(clk), .Q(
        \registers[34][6] ) );
  EDFFX1 \registers_reg[34][5]  ( .D(n8297), .E(n935), .CK(clk), .Q(
        \registers[34][5] ) );
  EDFFX1 \registers_reg[34][4]  ( .D(n8239), .E(n935), .CK(clk), .Q(
        \registers[34][4] ) );
  EDFFX1 \registers_reg[34][3]  ( .D(n8188), .E(n935), .CK(clk), .Q(
        \registers[34][3] ) );
  EDFFX1 \registers_reg[34][2]  ( .D(n8146), .E(n935), .CK(clk), .Q(
        \registers[34][2] ) );
  EDFFX1 \registers_reg[34][1]  ( .D(n8090), .E(n935), .CK(clk), .Q(
        \registers[34][1] ) );
  EDFFX1 \registers_reg[34][0]  ( .D(n8030), .E(n935), .CK(clk), .Q(
        \registers[34][0] ) );
  EDFFX1 \registers_reg[30][7]  ( .D(n8414), .E(n416), .CK(clk), .Q(
        \registers[30][7] ) );
  EDFFX1 \registers_reg[30][6]  ( .D(n8356), .E(n416), .CK(clk), .Q(
        \registers[30][6] ) );
  EDFFX1 \registers_reg[30][5]  ( .D(n8298), .E(n416), .CK(clk), .Q(
        \registers[30][5] ) );
  EDFFX1 \registers_reg[30][4]  ( .D(n8240), .E(n416), .CK(clk), .Q(
        \registers[30][4] ) );
  EDFFX1 \registers_reg[30][3]  ( .D(n8189), .E(n416), .CK(clk), .Q(
        \registers[30][3] ) );
  EDFFX1 \registers_reg[30][2]  ( .D(n8144), .E(n416), .CK(clk), .Q(
        \registers[30][2] ) );
  EDFFX1 \registers_reg[30][1]  ( .D(n8088), .E(n416), .CK(clk), .Q(
        \registers[30][1] ) );
  EDFFX1 \registers_reg[30][0]  ( .D(n8028), .E(n416), .CK(clk), .Q(
        \registers[30][0] ) );
  EDFFX1 \registers_reg[26][7]  ( .D(n8415), .E(n412), .CK(clk), .Q(
        \registers[26][7] ) );
  EDFFX1 \registers_reg[26][6]  ( .D(n8357), .E(n412), .CK(clk), .Q(
        \registers[26][6] ) );
  EDFFX1 \registers_reg[26][5]  ( .D(n8299), .E(n412), .CK(clk), .Q(
        \registers[26][5] ) );
  EDFFX1 \registers_reg[26][4]  ( .D(n8241), .E(n412), .CK(clk), .Q(
        \registers[26][4] ) );
  EDFFX1 \registers_reg[26][3]  ( .D(n8190), .E(n412), .CK(clk), .Q(
        \registers[26][3] ) );
  EDFFX1 \registers_reg[26][2]  ( .D(n8145), .E(n412), .CK(clk), .Q(
        \registers[26][2] ) );
  EDFFX1 \registers_reg[26][1]  ( .D(n8089), .E(n412), .CK(clk), .Q(
        \registers[26][1] ) );
  EDFFX1 \registers_reg[26][0]  ( .D(n8029), .E(n412), .CK(clk), .Q(
        \registers[26][0] ) );
  EDFFX1 \registers_reg[22][7]  ( .D(n8413), .E(n408), .CK(clk), .Q(
        \registers[22][7] ) );
  EDFFX1 \registers_reg[22][6]  ( .D(n8355), .E(n408), .CK(clk), .Q(
        \registers[22][6] ) );
  EDFFX1 \registers_reg[22][5]  ( .D(n8297), .E(n408), .CK(clk), .Q(
        \registers[22][5] ) );
  EDFFX1 \registers_reg[22][4]  ( .D(n8239), .E(n408), .CK(clk), .Q(
        \registers[22][4] ) );
  EDFFX1 \registers_reg[22][3]  ( .D(n8188), .E(n408), .CK(clk), .Q(
        \registers[22][3] ) );
  EDFFX1 \registers_reg[22][2]  ( .D(n8146), .E(n408), .CK(clk), .Q(
        \registers[22][2] ) );
  EDFFX1 \registers_reg[22][1]  ( .D(n8090), .E(n408), .CK(clk), .Q(
        \registers[22][1] ) );
  EDFFX1 \registers_reg[22][0]  ( .D(n8030), .E(n408), .CK(clk), .Q(
        \registers[22][0] ) );
  EDFFX1 \registers_reg[18][7]  ( .D(n8414), .E(n404), .CK(clk), .Q(
        \registers[18][7] ) );
  EDFFX1 \registers_reg[18][6]  ( .D(n8356), .E(n404), .CK(clk), .Q(
        \registers[18][6] ) );
  EDFFX1 \registers_reg[18][5]  ( .D(n8298), .E(n404), .CK(clk), .Q(
        \registers[18][5] ) );
  EDFFX1 \registers_reg[18][4]  ( .D(n8240), .E(n404), .CK(clk), .Q(
        \registers[18][4] ) );
  EDFFX1 \registers_reg[18][3]  ( .D(n8189), .E(n404), .CK(clk), .Q(
        \registers[18][3] ) );
  EDFFX1 \registers_reg[18][2]  ( .D(n8144), .E(n404), .CK(clk), .Q(
        \registers[18][2] ) );
  EDFFX1 \registers_reg[18][1]  ( .D(n8088), .E(n404), .CK(clk), .Q(
        \registers[18][1] ) );
  EDFFX1 \registers_reg[18][0]  ( .D(n8028), .E(n404), .CK(clk), .Q(
        \registers[18][0] ) );
  EDFFX1 \registers_reg[14][7]  ( .D(n8415), .E(n400), .CK(clk), .Q(
        \registers[14][7] ) );
  EDFFX1 \registers_reg[14][6]  ( .D(n8357), .E(n400), .CK(clk), .Q(
        \registers[14][6] ) );
  EDFFX1 \registers_reg[14][5]  ( .D(n8299), .E(n400), .CK(clk), .Q(
        \registers[14][5] ) );
  EDFFX1 \registers_reg[14][4]  ( .D(n8241), .E(n400), .CK(clk), .Q(
        \registers[14][4] ) );
  EDFFX1 \registers_reg[14][3]  ( .D(n8190), .E(n400), .CK(clk), .Q(
        \registers[14][3] ) );
  EDFFX1 \registers_reg[14][2]  ( .D(n8142), .E(n400), .CK(clk), .Q(
        \registers[14][2] ) );
  EDFFX1 \registers_reg[14][1]  ( .D(n8086), .E(n400), .CK(clk), .Q(
        \registers[14][1] ) );
  EDFFX1 \registers_reg[14][0]  ( .D(n8026), .E(n400), .CK(clk), .Q(
        \registers[14][0] ) );
  EDFFX1 \registers_reg[10][7]  ( .D(n8413), .E(n396), .CK(clk), .Q(
        \registers[10][7] ) );
  EDFFX1 \registers_reg[10][6]  ( .D(n8355), .E(n396), .CK(clk), .Q(
        \registers[10][6] ) );
  EDFFX1 \registers_reg[10][5]  ( .D(n8297), .E(n396), .CK(clk), .Q(
        \registers[10][5] ) );
  EDFFX1 \registers_reg[10][4]  ( .D(n8239), .E(n396), .CK(clk), .Q(
        \registers[10][4] ) );
  EDFFX1 \registers_reg[10][3]  ( .D(n8188), .E(n396), .CK(clk), .Q(
        \registers[10][3] ) );
  EDFFX1 \registers_reg[10][2]  ( .D(n8143), .E(n396), .CK(clk), .Q(
        \registers[10][2] ) );
  EDFFX1 \registers_reg[10][1]  ( .D(n8087), .E(n396), .CK(clk), .Q(
        \registers[10][1] ) );
  EDFFX1 \registers_reg[10][0]  ( .D(n8027), .E(n396), .CK(clk), .Q(
        \registers[10][0] ) );
  EDFFX1 \registers_reg[6][7]  ( .D(n8414), .E(n1016), .CK(clk), .Q(
        \registers[6][7] ) );
  EDFFX1 \registers_reg[6][6]  ( .D(n8356), .E(n1016), .CK(clk), .Q(
        \registers[6][6] ), .QN(n1127) );
  EDFFX1 \registers_reg[6][5]  ( .D(n8298), .E(n1016), .CK(clk), .Q(
        \registers[6][5] ), .QN(n1128) );
  EDFFX1 \registers_reg[6][4]  ( .D(n8240), .E(n1016), .CK(clk), .Q(
        \registers[6][4] ), .QN(n1129) );
  EDFFX1 \registers_reg[6][3]  ( .D(n8189), .E(n1016), .CK(clk), .Q(
        \registers[6][3] ), .QN(n1130) );
  EDFFX1 \registers_reg[6][2]  ( .D(n8141), .E(n1016), .CK(clk), .Q(
        \registers[6][2] ), .QN(n1131) );
  EDFFX1 \registers_reg[6][1]  ( .D(n8085), .E(n1016), .CK(clk), .Q(
        \registers[6][1] ), .QN(n1132) );
  EDFFX1 \registers_reg[6][0]  ( .D(n8025), .E(n1016), .CK(clk), .Q(
        \registers[6][0] ), .QN(n1133) );
  EDFFX1 \registers_reg[2][7]  ( .D(n8410), .E(n392), .CK(clk), .Q(
        \registers[2][7] ) );
  EDFFX1 \registers_reg[2][6]  ( .D(n8352), .E(n392), .CK(clk), .Q(
        \registers[2][6] ) );
  EDFFX1 \registers_reg[2][5]  ( .D(n8294), .E(n392), .CK(clk), .Q(
        \registers[2][5] ) );
  EDFFX1 \registers_reg[2][4]  ( .D(n8236), .E(n392), .CK(clk), .Q(
        \registers[2][4] ) );
  EDFFX1 \registers_reg[2][3]  ( .D(n8190), .E(n392), .CK(clk), .Q(
        \registers[2][3] ) );
  EDFFX1 \registers_reg[2][2]  ( .D(n8142), .E(n392), .CK(clk), .Q(
        \registers[2][2] ) );
  EDFFX1 \registers_reg[2][1]  ( .D(n8086), .E(n392), .CK(clk), .Q(
        \registers[2][1] ) );
  EDFFX1 \registers_reg[2][0]  ( .D(n8026), .E(n392), .CK(clk), .Q(
        \registers[2][0] ) );
  EDFFX1 \registers_reg[4][1]  ( .D(n8087), .E(n1014), .CK(clk), .Q(
        \registers[4][1] ) );
  EDFFX1 \registers_reg[4][0]  ( .D(n8027), .E(n1014), .CK(clk), .Q(
        \registers[4][0] ) );
  DFFHQX1 \registers_reg[0][7]  ( .D(n2436), .CK(clk), .Q(\registers[0][7] )
         );
  DFFHQX1 \registers_reg[0][6]  ( .D(n2435), .CK(clk), .Q(\registers[0][6] )
         );
  DFFHQX1 \registers_reg[0][5]  ( .D(n2434), .CK(clk), .Q(\registers[0][5] )
         );
  DFFHQX1 \registers_reg[0][4]  ( .D(n2433), .CK(clk), .Q(\registers[0][4] )
         );
  DFFHQX1 \registers_reg[0][3]  ( .D(n2432), .CK(clk), .Q(\registers[0][3] )
         );
  DFFHQX1 \registers_reg[0][2]  ( .D(n2431), .CK(clk), .Q(\registers[0][2] )
         );
  DFFHQX1 \registers_reg[0][1]  ( .D(n2430), .CK(clk), .Q(\registers[0][1] )
         );
  DFFHQX1 \registers_reg[0][0]  ( .D(n2429), .CK(clk), .Q(\registers[0][0] )
         );
  DFFHQX1 \param_i_reg[2]  ( .D(n2426), .CK(clk), .Q(param_i[2]) );
  DFFHQX1 \param_i_reg[1]  ( .D(n2427), .CK(clk), .Q(param_i[1]) );
  DFFHQX1 StartBit_reg ( .D(n8957), .CK(clk), .Q(StartBit) );
  DFFHQX1 \state_reg[0]  ( .D(n8921), .CK(clk), .Q(state[0]) );
  DFFHQX1 \state_reg[1]  ( .D(n8922), .CK(clk), .Q(state[1]) );
  DFFTRX1 ena_out_reg ( .D(n1261), .RN(n1212), .CK(clk), .Q(ena_out) );
  DFFHQX1 \params_reg[20]  ( .D(n2409), .CK(clk), .Q(params[20]) );
  DFFHQX1 \params_reg[19]  ( .D(n2410), .CK(clk), .Q(params[19]) );
  DFFHQX1 \block_i_reg[18]  ( .D(n8938), .CK(clk), .Q(block_i[18]) );
  DFFHQX1 \block_i_reg[17]  ( .D(n8956), .CK(clk), .Q(block_i[17]) );
  DFFHQX1 \params_reg[16]  ( .D(n2413), .CK(clk), .Q(params[16]) );
  DFFHQX1 \pixel_i_reg[12]  ( .D(n8924), .CK(clk), .Q(pixel_i[12]) );
  DFFHQX1 \params_reg[13]  ( .D(n2416), .CK(clk), .Q(params[13]) );
  DFFHQX1 \params_reg[14]  ( .D(n2415), .CK(clk), .Q(params[14]) );
  DFFHQX1 \block_i_reg[15]  ( .D(n8954), .CK(clk), .Q(block_i[15]) );
  DFFHQX1 \block_i_reg[16]  ( .D(n8955), .CK(clk), .Q(block_i[16]) );
  DFFHQX1 \params_reg[15]  ( .D(n2414), .CK(clk), .Q(params[15]) );
  DFFHQX1 \params_reg[18]  ( .D(n2411), .CK(clk), .Q(params[18]) );
  DFFHQX1 \pixel_i_reg[11]  ( .D(n8936), .CK(clk), .Q(pixel_i[11]) );
  DFFHQX1 \pixel_i_reg[10]  ( .D(n8935), .CK(clk), .Q(pixel_i[10]) );
  DFFHQX1 \block_i_reg[13]  ( .D(n8952), .CK(clk), .Q(block_i[13]) );
  DFFHQX1 \block_i_reg[14]  ( .D(n8953), .CK(clk), .Q(block_i[14]) );
  DFFHQX1 \params_reg[17]  ( .D(n2412), .CK(clk), .Q(params[17]) );
  DFFHQX1 \block_i_reg[12]  ( .D(n8951), .CK(clk), .Q(block_i[12]) );
  DFFHQX1 \block_i_reg[10]  ( .D(n8949), .CK(clk), .Q(block_i[10]) );
  DFFHQX1 \block_i_reg[11]  ( .D(n8950), .CK(clk), .Q(block_i[11]) );
  DFFHQX1 \block_i_reg[9]  ( .D(n8948), .CK(clk), .Q(block_i[9]) );
  DFFHQX1 \block_i_reg[8]  ( .D(n8947), .CK(clk), .Q(block_i[8]) );
  DFFHQX1 \block_i_reg[5]  ( .D(n8944), .CK(clk), .Q(block_i[5]) );
  DFFHQX1 \block_i_reg[6]  ( .D(n8945), .CK(clk), .Q(block_i[6]) );
  DFFHQX1 \block_i_reg[7]  ( .D(n8946), .CK(clk), .Q(block_i[7]) );
  DFFHQX1 \block_i_reg[4]  ( .D(n8943), .CK(clk), .Q(block_i[4]) );
  DFFHQX1 \block_i_reg[1]  ( .D(n8940), .CK(clk), .Q(block_i[1]) );
  DFFHQX1 \block_i_reg[2]  ( .D(n8941), .CK(clk), .Q(block_i[2]) );
  DFFHQX1 \block_i_reg[3]  ( .D(n8942), .CK(clk), .Q(block_i[3]) );
  EDFFX1 \params_reg[11]  ( .D(\registers[4][0] ), .E(n1044), .CK(clk), .Q(
        params[11]) );
  EDFFX1 \N2_reg[0]  ( .D(N128), .E(n8438), .CK(clk), .Q(N2[0]) );
  EDFFX1 \N2_reg[1]  ( .D(1'b0), .E(n1034), .CK(clk), .Q(N2[1]) );
  EDFFX1 \N2_reg[2]  ( .D(N130), .E(n1034), .CK(clk), .Q(N2[2]) );
  EDFFX1 \N2_reg[3]  ( .D(N131), .E(n1034), .CK(clk), .Q(N2[3]) );
  EDFFX1 \N2_reg[4]  ( .D(N132), .E(n1034), .CK(clk), .Q(N2[4]) );
  EDFFX1 \W_block_reg[31]  ( .D(N1308), .E(n1043), .CK(clk), .Q(W_block[31])
         );
  EDFFX1 \W_block_reg[30]  ( .D(N1309), .E(n1043), .CK(clk), .Q(W_block[30])
         );
  EDFFX1 \W_block_reg[15]  ( .D(N1308), .E(n1041), .CK(clk), .Q(W_block[15])
         );
  EDFFX1 \W_block_reg[14]  ( .D(N1309), .E(n1041), .CK(clk), .Q(W_block[14])
         );
  EDFFX1 \W_block_reg[23]  ( .D(N1308), .E(n1037), .CK(clk), .Q(W_block[23])
         );
  EDFFX1 \W_block_reg[22]  ( .D(N1309), .E(n1037), .CK(clk), .Q(W_block[22])
         );
  EDFFX1 \W_block_reg[7]  ( .D(N1308), .E(n1036), .CK(clk), .Q(W_block[7]) );
  EDFFX1 \W_block_reg[6]  ( .D(N1309), .E(n1036), .CK(clk), .Q(W_block[6]) );
  EDFFX1 \N2_reg[5]  ( .D(N133), .E(n1034), .CK(clk), .Q(N2[5]) );
  EDFFX1 \W_block_reg[29]  ( .D(N1310), .E(n1043), .CK(clk), .Q(W_block[29])
         );
  EDFFX1 \W_block_reg[28]  ( .D(N1311), .E(n1043), .CK(clk), .Q(W_block[28])
         );
  EDFFX1 \W_block_reg[27]  ( .D(N1312), .E(n1043), .CK(clk), .Q(W_block[27])
         );
  EDFFX1 \W_block_reg[26]  ( .D(N1313), .E(n1043), .CK(clk), .Q(W_block[26])
         );
  EDFFX1 \W_block_reg[25]  ( .D(N1314), .E(n1043), .CK(clk), .Q(W_block[25])
         );
  EDFFX1 \W_block_reg[24]  ( .D(N1315), .E(n1043), .CK(clk), .Q(W_block[24])
         );
  EDFFX1 \W_block_reg[13]  ( .D(N1310), .E(n1041), .CK(clk), .Q(W_block[13])
         );
  EDFFX1 \W_block_reg[12]  ( .D(N1311), .E(n1041), .CK(clk), .Q(W_block[12])
         );
  EDFFX1 \W_block_reg[11]  ( .D(N1312), .E(n1041), .CK(clk), .Q(W_block[11])
         );
  EDFFX1 \W_block_reg[10]  ( .D(N1313), .E(n1041), .CK(clk), .Q(W_block[10])
         );
  EDFFX1 \W_block_reg[9]  ( .D(N1314), .E(n1041), .CK(clk), .Q(W_block[9]) );
  EDFFX1 \W_block_reg[8]  ( .D(N1315), .E(n1041), .CK(clk), .Q(W_block[8]) );
  EDFFX1 \W_block_reg[21]  ( .D(N1310), .E(n1037), .CK(clk), .Q(W_block[21])
         );
  EDFFX1 \W_block_reg[20]  ( .D(N1311), .E(n1037), .CK(clk), .Q(W_block[20])
         );
  EDFFX1 \W_block_reg[19]  ( .D(N1312), .E(n1037), .CK(clk), .Q(W_block[19])
         );
  EDFFX1 \W_block_reg[18]  ( .D(N1313), .E(n1037), .CK(clk), .Q(W_block[18])
         );
  EDFFX1 \W_block_reg[17]  ( .D(N1314), .E(n1037), .CK(clk), .Q(W_block[17])
         );
  EDFFX1 \W_block_reg[16]  ( .D(N1315), .E(n1037), .CK(clk), .Q(W_block[16])
         );
  EDFFX1 \W_block_reg[5]  ( .D(N1310), .E(n1036), .CK(clk), .Q(W_block[5]) );
  EDFFX1 \W_block_reg[4]  ( .D(N1311), .E(n1036), .CK(clk), .Q(W_block[4]) );
  EDFFX1 \W_block_reg[3]  ( .D(N1312), .E(n1036), .CK(clk), .Q(W_block[3]) );
  EDFFX1 \W_block_reg[2]  ( .D(N1313), .E(n1036), .CK(clk), .Q(W_block[2]) );
  EDFFX1 \W_block_reg[1]  ( .D(N1314), .E(n1036), .CK(clk), .Q(W_block[1]) );
  EDFFX1 \W_block_reg[0]  ( .D(N1315), .E(n1036), .CK(clk), .Q(W_block[0]) );
  EDFFX1 \Im_block_reg[31]  ( .D(N1227), .E(n1040), .CK(clk), .Q(Im_block[31])
         );
  EDFFX1 \Im_block_reg[30]  ( .D(N1228), .E(n1040), .CK(clk), .Q(Im_block[30])
         );
  EDFFX1 \Im_block_reg[29]  ( .D(N1229), .E(n1040), .CK(clk), .Q(Im_block[29])
         );
  EDFFX1 \Im_block_reg[15]  ( .D(N1227), .E(n1042), .CK(clk), .Q(Im_block[15])
         );
  EDFFX1 \Im_block_reg[14]  ( .D(N1228), .E(n1042), .CK(clk), .Q(Im_block[14])
         );
  EDFFX1 \Im_block_reg[23]  ( .D(N1227), .E(n1039), .CK(clk), .Q(Im_block[23])
         );
  EDFFX1 \Im_block_reg[22]  ( .D(N1228), .E(n1039), .CK(clk), .Q(Im_block[22])
         );
  EDFFX1 \Im_block_reg[21]  ( .D(N1229), .E(n1039), .CK(clk), .Q(Im_block[21])
         );
  EDFFX1 \Im_block_reg[7]  ( .D(N1227), .E(n1038), .CK(clk), .Q(Im_block[7])
         );
  EDFFX1 \Im_block_reg[6]  ( .D(N1228), .E(n1038), .CK(clk), .Q(Im_block[6])
         );
  EDFFX1 \Im_block_reg[28]  ( .D(N1230), .E(n1040), .CK(clk), .Q(Im_block[28])
         );
  EDFFX1 \Im_block_reg[27]  ( .D(N1231), .E(n1040), .CK(clk), .Q(Im_block[27])
         );
  EDFFX1 \Im_block_reg[26]  ( .D(N1232), .E(n1040), .CK(clk), .Q(Im_block[26])
         );
  EDFFX1 \Im_block_reg[25]  ( .D(N1233), .E(n1040), .CK(clk), .Q(Im_block[25])
         );
  EDFFX1 \Im_block_reg[24]  ( .D(N1234), .E(n1040), .CK(clk), .Q(Im_block[24])
         );
  EDFFX1 \Im_block_reg[13]  ( .D(N1229), .E(n1042), .CK(clk), .Q(Im_block[13])
         );
  EDFFX1 \Im_block_reg[12]  ( .D(N1230), .E(n1042), .CK(clk), .Q(Im_block[12])
         );
  EDFFX1 \Im_block_reg[11]  ( .D(N1231), .E(n1042), .CK(clk), .Q(Im_block[11])
         );
  EDFFX1 \Im_block_reg[10]  ( .D(N1232), .E(n1042), .CK(clk), .Q(Im_block[10])
         );
  EDFFX1 \Im_block_reg[9]  ( .D(N1233), .E(n1042), .CK(clk), .Q(Im_block[9])
         );
  EDFFX1 \Im_block_reg[8]  ( .D(N1234), .E(n1042), .CK(clk), .Q(Im_block[8])
         );
  EDFFX1 \Im_block_reg[20]  ( .D(N1230), .E(n1039), .CK(clk), .Q(Im_block[20])
         );
  EDFFX1 \Im_block_reg[19]  ( .D(N1231), .E(n1039), .CK(clk), .Q(Im_block[19])
         );
  EDFFX1 \Im_block_reg[18]  ( .D(N1232), .E(n1039), .CK(clk), .Q(Im_block[18])
         );
  EDFFX1 \Im_block_reg[17]  ( .D(N1233), .E(n1039), .CK(clk), .Q(Im_block[17])
         );
  EDFFX1 \Im_block_reg[16]  ( .D(N1234), .E(n1039), .CK(clk), .Q(Im_block[16])
         );
  EDFFX1 \Im_block_reg[5]  ( .D(N1229), .E(n1038), .CK(clk), .Q(Im_block[5])
         );
  EDFFX1 \Im_block_reg[4]  ( .D(N1230), .E(n1038), .CK(clk), .Q(Im_block[4])
         );
  EDFFX1 \Im_block_reg[3]  ( .D(N1231), .E(n1038), .CK(clk), .Q(Im_block[3])
         );
  EDFFX1 \Im_block_reg[2]  ( .D(N1232), .E(n1038), .CK(clk), .Q(Im_block[2])
         );
  EDFFX1 \Im_block_reg[1]  ( .D(N1233), .E(n1038), .CK(clk), .Q(Im_block[1])
         );
  EDFFX1 \Im_block_reg[0]  ( .D(N1234), .E(n1038), .CK(clk), .Q(Im_block[0])
         );
  EDFFX1 \N2_reg[6]  ( .D(N134), .E(n1034), .CK(clk), .Q(N2[6]) );
  EDFFX1 \N2_reg[7]  ( .D(N135), .E(n1034), .CK(clk), .Q(N2[7]) );
  EDFFX1 \N2_reg[8]  ( .D(N136), .E(n1034), .CK(clk), .Q(N2[8]) );
  EDFFX1 \N2_reg[9]  ( .D(N137), .E(n1034), .CK(clk), .Q(N2[9]) );
  EDFFX1 \N2_reg[10]  ( .D(N138), .E(n8438), .CK(clk), .Q(N2[10]) );
  EDFFX1 \N2_reg[11]  ( .D(N139), .E(n8438), .CK(clk), .Q(N2[11]) );
  EDFFX1 \N2_reg[12]  ( .D(N140), .E(n8438), .CK(clk), .Q(N2[12]) );
  EDFFX1 \N2_reg[13]  ( .D(N141), .E(n8438), .CK(clk), .Q(N2[13]) );
  EDFFX1 \N2_reg[14]  ( .D(N142), .E(n8438), .CK(clk), .Q(N2[14]) );
  EDFFX1 \N2_reg[15]  ( .D(N143), .E(n8438), .CK(clk), .Q(N2[15]) );
  EDFFX1 \N2_reg[16]  ( .D(N144), .E(n8438), .CK(clk), .Q(N2[16]) );
  EDFFX1 \N2_reg[17]  ( .D(N145), .E(n8438), .CK(clk), .Q(N2[17]) );
  EDFFX1 \N2_reg[18]  ( .D(N146), .E(n8438), .CK(clk), .Q(N2[18]) );
  DFFHQX1 \params_reg[7]  ( .D(n2417), .CK(clk), .Q(params[7]) );
  DFFHQX1 \params_reg[6]  ( .D(n2418), .CK(clk), .Q(params[6]) );
  DFFHQX1 \params_reg[5]  ( .D(n2419), .CK(clk), .Q(params[5]) );
  EDFFX1 \N2_reg[19]  ( .D(N147), .E(n8438), .CK(clk), .Q(N2[19]) );
  DFFHQX1 \params_reg[4]  ( .D(n2420), .CK(clk), .Q(params[4]) );
  EDFFX2 \M2_reg[1]  ( .D(1'b0), .E(n8437), .CK(clk), .Q(M2[1]) );
  EDFFX2 \M2_reg[2]  ( .D(N110), .E(n8437), .CK(clk), .Q(M2[2]) );
  DFFHQX1 \params_reg[3]  ( .D(n2421), .CK(clk), .Q(params[3]) );
  DFFHQX1 \params_reg[2]  ( .D(n2422), .CK(clk), .Q(params[2]) );
  DFFHQX1 \params_reg[1]  ( .D(n2423), .CK(clk), .Q(params[1]) );
  EDFFX2 \M2_reg[4]  ( .D(N112), .E(n8437), .CK(clk), .Q(M2[4]) );
  EDFFX2 \M2_reg[5]  ( .D(N113), .E(n8437), .CK(clk), .Q(M2[5]) );
  EDFFX2 \params_reg[10]  ( .D(M2[2]), .E(n1044), .CK(clk), .Q(params[10]) );
  EDFFX1 \M2_reg[0]  ( .D(N108), .E(n8437), .CK(clk), .Q(M2[0]) );
  EDFFX1 \params_reg[8]  ( .D(M2[0]), .E(n1044), .CK(clk), .Q(params[8]) );
  EDFFX1 \M2_reg[6]  ( .D(N114), .E(n8437), .CK(clk), .Q(M2[6]), .QN(n7) );
  DFFHQX1 \params_reg[0]  ( .D(n2424), .CK(clk), .Q(params[0]) );
  EDFFX2 \M2_reg[7]  ( .D(N115), .E(n8437), .CK(clk), .Q(M2[7]) );
  EDFFX2 \M2_reg[8]  ( .D(N116), .E(n8437), .CK(clk), .Q(M2[8]) );
  EDFFX2 \params_reg[9]  ( .D(M2[1]), .E(n1044), .CK(clk), .Q(params[9]) );
  EDFFX1 \M2_reg[9]  ( .D(N117), .E(n8437), .CK(clk), .Q(M2[9]), .QN(n6) );
  EDFFX1 \M2_reg[11]  ( .D(N119), .E(n1035), .CK(clk), .Q(M2[11]) );
  EDFFX1 \M2_reg[10]  ( .D(N118), .E(n1035), .CK(clk), .Q(M2[10]) );
  EDFFX1 \M2_reg[15]  ( .D(N123), .E(n1035), .CK(clk), .Q(M2[15]) );
  EDFFX1 \M2_reg[13]  ( .D(N121), .E(n1035), .CK(clk), .Q(M2[13]) );
  EDFFX1 \M2_reg[14]  ( .D(N122), .E(n1035), .CK(clk), .Q(M2[14]) );
  EDFFX1 \M2_reg[12]  ( .D(N120), .E(n1035), .CK(clk), .Q(M2[12]) );
  EDFFX1 \M2_reg[18]  ( .D(N126), .E(n1035), .CK(clk), .Q(M2[18]) );
  EDFFX1 \M2_reg[16]  ( .D(N124), .E(n1035), .CK(clk), .Q(M2[16]) );
  EDFFX1 \M2_reg[19]  ( .D(N127), .E(n1035), .CK(clk), .Q(M2[19]) );
  EDFFX1 \M2_reg[17]  ( .D(N125), .E(n1035), .CK(clk), .Q(M2[17]) );
  DFFHQX1 \params_reg[46]  ( .D(n2383), .CK(clk), .Q(params[46]) );
  DFFHQX1 \params_reg[45]  ( .D(n2384), .CK(clk), .Q(params[45]) );
  DFFHQX1 \params_reg[40]  ( .D(n2389), .CK(clk), .Q(params[40]) );
  DFFHQX1 \params_reg[44]  ( .D(n2385), .CK(clk), .Q(params[44]) );
  DFFHQX1 \params_reg[43]  ( .D(n2386), .CK(clk), .Q(params[43]) );
  DFFHQX1 \params_reg[42]  ( .D(n2387), .CK(clk), .Q(params[42]) );
  DFFHQX1 \params_reg[41]  ( .D(n2388), .CK(clk), .Q(params[41]) );
  DFFHQX1 \params_reg[39]  ( .D(n2390), .CK(clk), .Q(params[39]) );
  DFFHQX1 \params_reg[37]  ( .D(n2392), .CK(clk), .Q(params[37]) );
  DFFHQX1 \params_reg[38]  ( .D(n2391), .CK(clk), .Q(params[38]) );
  DFFHQX1 \params_reg[36]  ( .D(n2393), .CK(clk), .Q(params[36]) );
  DFFHQX1 \params_reg[34]  ( .D(n2395), .CK(clk), .Q(params[34]) );
  DFFHQX1 \params_reg[33]  ( .D(n2396), .CK(clk), .Q(params[33]) );
  DFFHQX1 \params_reg[26]  ( .D(n2403), .CK(clk), .Q(params[26]) );
  DFFHQX1 \params_reg[27]  ( .D(n2402), .CK(clk), .Q(params[27]) );
  DFFHQX1 \params_reg[32]  ( .D(n2397), .CK(clk), .Q(params[32]) );
  DFFHQX1 \params_reg[31]  ( .D(n2398), .CK(clk), .Q(params[31]) );
  DFFHQX1 \params_reg[25]  ( .D(n2404), .CK(clk), .Q(params[25]) );
  DFFHQX1 \params_reg[24]  ( .D(n2405), .CK(clk), .Q(params[24]) );
  DFFHQX1 \params_reg[30]  ( .D(n2399), .CK(clk), .Q(params[30]) );
  DFFHQX1 \params_reg[23]  ( .D(n2406), .CK(clk), .Q(params[23]) );
  DFFHQX1 \params_reg[29]  ( .D(n2400), .CK(clk), .Q(params[29]) );
  DFFHQX1 \params_reg[22]  ( .D(n2407), .CK(clk), .Q(params[22]) );
  DFFHQX1 \params_reg[28]  ( .D(n2401), .CK(clk), .Q(params[28]) );
  DFFHQX1 \params_reg[21]  ( .D(n2408), .CK(clk), .Q(params[21]) );
  DFFHQX1 \pixel_i_reg[8]  ( .D(n8933), .CK(clk), .Q(pixel_i[8]) );
  DFFHQX1 \pixel_i_reg[5]  ( .D(n8930), .CK(clk), .Q(pixel_i[5]) );
  EDFFX1 \params_reg[12]  ( .D(\registers[4][1] ), .E(n1044), .CK(clk), .Q(
        params[12]) );
  DFFHQX1 \params_reg[35]  ( .D(n2394), .CK(clk), .Q(params[35]) );
  EDFFX1 \M2_reg[3]  ( .D(N111), .E(n8437), .CK(clk), .Q(M2[3]), .QN(n5) );
  DFFHQX4 \pixel_i_reg[0]  ( .D(n8925), .CK(clk), .Q(N1197) );
  DFFHQX2 \pixel_i_reg[3]  ( .D(n8928), .CK(clk), .Q(pixel_i[3]) );
  DFFHQX2 \pixel_i_reg[6]  ( .D(n8931), .CK(clk), .Q(pixel_i[6]) );
  DFFHQX2 \pixel_i_reg[1]  ( .D(n8926), .CK(clk), .Q(pixel_i[1]) );
  DFFHQX2 \param_i_reg[0]  ( .D(n2428), .CK(clk), .Q(param_i[0]) );
  DFFHQX2 \pixel_i_reg[9]  ( .D(n8934), .CK(clk), .Q(pixel_i[9]) );
  DFFHQX2 \pixel_i_reg[4]  ( .D(n8929), .CK(clk), .Q(pixel_i[4]) );
  DFFHQX2 \pixel_i_reg[7]  ( .D(n8932), .CK(clk), .Q(pixel_i[7]) );
  DFFHQX2 \pixel_i_reg[2]  ( .D(n8927), .CK(clk), .Q(pixel_i[2]) );
  DFFHQX2 \block_i_reg[0]  ( .D(n8939), .CK(clk), .Q(block_i[0]) );
  OAI31X1 U3 ( .A0(n8963), .A1(n1241), .A2(n8960), .B0(n8973), .Y(n1261) );
  INVX1 U4 ( .A(n8), .Y(n9) );
  INVX1 U5 ( .A(pixel_i[5]), .Y(n8) );
  OR4X1 U6 ( .A(pixel_i[6]), .B(pixel_i[7]), .C(pixel_i[8]), .D(pixel_i[9]), 
        .Y(n1215) );
  NOR4BX2 U7 ( .AN(n8914), .B(M2[14]), .C(n8913), .D(M2[13]), .Y(N1195) );
  AOI22XL U8 ( .A0(N1349), .A1(n8442), .B0(block_i[0]), .B1(n8435), .Y(n1235)
         );
  NOR4XL U9 ( .A(pixel_i[3]), .B(n1215), .C(n9), .D(pixel_i[4]), .Y(n1214) );
  AOI22XL U10 ( .A0(n8440), .A1(n9), .B0(N1240), .B1(n8441), .Y(n1250) );
  AOI22XL U16 ( .A0(n8440), .A1(pixel_i[8]), .B0(N1243), .B1(n8441), .Y(n1247)
         );
  INVX1 U17 ( .A(param_i[2]), .Y(n8966) );
  INVX1 U18 ( .A(param_i[0]), .Y(n8964) );
  CLKINVX3 U19 ( .A(n7443), .Y(n7461) );
  CLKINVX3 U20 ( .A(n7442), .Y(n7462) );
  CLKINVX3 U21 ( .A(n7444), .Y(n7458) );
  CLKINVX3 U22 ( .A(n7443), .Y(n7460) );
  CLKINVX3 U23 ( .A(n7443), .Y(n7459) );
  CLKINVX3 U24 ( .A(n7441), .Y(n7466) );
  CLKINVX3 U25 ( .A(n7441), .Y(n7467) );
  CLKINVX3 U26 ( .A(n7442), .Y(n7463) );
  CLKINVX3 U27 ( .A(n7442), .Y(n7464) );
  CLKINVX3 U28 ( .A(n7441), .Y(n7465) );
  CLKINVX3 U29 ( .A(n7446), .Y(n7450) );
  CLKINVX3 U30 ( .A(n7446), .Y(n7451) );
  CLKINVX3 U31 ( .A(n7447), .Y(n7448) );
  CLKINVX3 U32 ( .A(n7447), .Y(n7449) );
  CLKINVX3 U33 ( .A(n7444), .Y(n7456) );
  CLKINVX3 U34 ( .A(n7444), .Y(n7457) );
  CLKINVX3 U35 ( .A(n7446), .Y(n7452) );
  CLKINVX3 U36 ( .A(n7445), .Y(n7453) );
  CLKINVX3 U37 ( .A(n7445), .Y(n7455) );
  CLKINVX3 U38 ( .A(n7445), .Y(n7454) );
  CLKINVX3 U39 ( .A(n7436), .Y(n7482) );
  CLKINVX3 U40 ( .A(n7435), .Y(n7483) );
  CLKINVX3 U41 ( .A(n7436), .Y(n7480) );
  CLKINVX3 U42 ( .A(n7436), .Y(n7481) );
  CLKINVX3 U43 ( .A(n7434), .Y(n7488) );
  CLKINVX3 U44 ( .A(n7433), .Y(n7489) );
  CLKINVX3 U45 ( .A(n7435), .Y(n7484) );
  CLKINVX3 U46 ( .A(n7435), .Y(n7485) );
  CLKINVX3 U47 ( .A(n7434), .Y(n7487) );
  CLKINVX3 U48 ( .A(n7434), .Y(n7486) );
  CLKINVX3 U49 ( .A(n7439), .Y(n7472) );
  CLKINVX3 U50 ( .A(n7439), .Y(n7473) );
  CLKINVX3 U51 ( .A(n7440), .Y(n7468) );
  CLKINVX3 U52 ( .A(n7440), .Y(n7469) );
  CLKINVX3 U53 ( .A(n7439), .Y(n7471) );
  CLKINVX3 U54 ( .A(n7440), .Y(n7470) );
  CLKINVX3 U55 ( .A(n7437), .Y(n7477) );
  CLKINVX3 U56 ( .A(n7437), .Y(n7479) );
  CLKINVX3 U57 ( .A(n7437), .Y(n7478) );
  CLKINVX3 U58 ( .A(n7438), .Y(n7474) );
  CLKINVX3 U59 ( .A(n7438), .Y(n7476) );
  CLKINVX3 U60 ( .A(n7438), .Y(n7475) );
  CLKINVX3 U61 ( .A(n7428), .Y(n7504) );
  CLKINVX3 U62 ( .A(n7428), .Y(n7505) );
  CLKINVX3 U63 ( .A(n7429), .Y(n7501) );
  CLKINVX3 U64 ( .A(n7429), .Y(n7503) );
  CLKINVX3 U65 ( .A(n7429), .Y(n7502) );
  CLKINVX3 U66 ( .A(n7427), .Y(n7509) );
  CLKINVX3 U67 ( .A(n7426), .Y(n7510) );
  CLKINVX3 U68 ( .A(n7428), .Y(n7506) );
  CLKINVX3 U69 ( .A(n7427), .Y(n7508) );
  CLKINVX3 U70 ( .A(n7427), .Y(n7507) );
  CLKINVX3 U71 ( .A(n7432), .Y(n7493) );
  CLKINVX3 U72 ( .A(n7432), .Y(n7494) );
  CLKINVX3 U73 ( .A(n7433), .Y(n7490) );
  CLKINVX3 U74 ( .A(n7432), .Y(n7492) );
  CLKINVX3 U75 ( .A(n7433), .Y(n7491) );
  CLKINVX3 U76 ( .A(n7430), .Y(n7498) );
  CLKINVX3 U77 ( .A(n7430), .Y(n7500) );
  CLKINVX3 U78 ( .A(n7430), .Y(n7499) );
  CLKINVX3 U79 ( .A(n7431), .Y(n7495) );
  CLKINVX3 U80 ( .A(n7431), .Y(n7496) );
  CLKINVX3 U81 ( .A(n7431), .Y(n7497) );
  CLKINVX3 U82 ( .A(n7421), .Y(n7525) );
  CLKINVX3 U83 ( .A(n7421), .Y(n7526) );
  CLKINVX3 U84 ( .A(n7422), .Y(n7522) );
  CLKINVX3 U85 ( .A(n7422), .Y(n7524) );
  CLKINVX3 U86 ( .A(n7422), .Y(n7523) );
  CLKINVX3 U87 ( .A(n7420), .Y(n7530) );
  CLKINVX3 U88 ( .A(n7419), .Y(n7531) );
  CLKINVX3 U89 ( .A(n7421), .Y(n7527) );
  CLKINVX3 U90 ( .A(n7420), .Y(n7528) );
  CLKINVX3 U91 ( .A(n7420), .Y(n7529) );
  CLKINVX3 U92 ( .A(n7425), .Y(n7514) );
  CLKINVX3 U93 ( .A(n7425), .Y(n7515) );
  CLKINVX3 U94 ( .A(n7426), .Y(n7511) );
  CLKINVX3 U95 ( .A(n7426), .Y(n7512) );
  CLKINVX3 U96 ( .A(n7425), .Y(n7513) );
  CLKINVX3 U97 ( .A(n7423), .Y(n7520) );
  CLKINVX3 U98 ( .A(n7423), .Y(n7521) );
  CLKINVX3 U99 ( .A(n7424), .Y(n7516) );
  CLKINVX3 U100 ( .A(n7424), .Y(n7517) );
  CLKINVX3 U101 ( .A(n7423), .Y(n7519) );
  CLKINVX3 U102 ( .A(n7424), .Y(n7518) );
  CLKINVX3 U103 ( .A(n7414), .Y(n7546) );
  CLKINVX3 U104 ( .A(n7414), .Y(n7547) );
  CLKINVX3 U105 ( .A(n7415), .Y(n7544) );
  CLKINVX3 U106 ( .A(n7415), .Y(n7545) );
  CLKINVX3 U107 ( .A(n7412), .Y(n7552) );
  CLKINVX3 U108 ( .A(n7412), .Y(n7553) );
  CLKINVX3 U109 ( .A(n7414), .Y(n7548) );
  CLKINVX3 U110 ( .A(n7413), .Y(n7549) );
  CLKINVX3 U111 ( .A(n7413), .Y(n7551) );
  CLKINVX3 U112 ( .A(n7413), .Y(n7550) );
  CLKINVX3 U113 ( .A(n7418), .Y(n7536) );
  CLKINVX3 U114 ( .A(n7417), .Y(n7537) );
  CLKINVX3 U115 ( .A(n7419), .Y(n7532) );
  CLKINVX3 U116 ( .A(n7419), .Y(n7533) );
  CLKINVX3 U117 ( .A(n7418), .Y(n7535) );
  CLKINVX3 U118 ( .A(n7418), .Y(n7534) );
  CLKINVX3 U119 ( .A(n7416), .Y(n7541) );
  CLKINVX3 U120 ( .A(n7415), .Y(n7543) );
  CLKINVX3 U121 ( .A(n7416), .Y(n7542) );
  CLKINVX3 U122 ( .A(n7417), .Y(n7538) );
  CLKINVX3 U123 ( .A(n7416), .Y(n7540) );
  CLKINVX3 U124 ( .A(n7417), .Y(n7539) );
  CLKINVX3 U125 ( .A(n7407), .Y(n7568) );
  CLKINVX3 U126 ( .A(n7407), .Y(n7569) );
  CLKINVX3 U127 ( .A(n7408), .Y(n7565) );
  CLKINVX3 U128 ( .A(n7407), .Y(n7567) );
  CLKINVX3 U129 ( .A(n7408), .Y(n7566) );
  CLKINVX3 U130 ( .A(n7405), .Y(n7573) );
  CLKINVX3 U131 ( .A(n7405), .Y(n7574) );
  CLKINVX3 U132 ( .A(n7406), .Y(n7570) );
  CLKINVX3 U133 ( .A(n7406), .Y(n7572) );
  CLKINVX3 U134 ( .A(n7406), .Y(n7571) );
  CLKINVX3 U135 ( .A(n7411), .Y(n7557) );
  CLKINVX3 U136 ( .A(n7410), .Y(n7558) );
  CLKINVX3 U137 ( .A(n7412), .Y(n7554) );
  CLKINVX3 U138 ( .A(n7411), .Y(n7556) );
  CLKINVX3 U139 ( .A(n7411), .Y(n7555) );
  CLKINVX3 U140 ( .A(n7409), .Y(n7562) );
  CLKINVX3 U141 ( .A(n7408), .Y(n7564) );
  CLKINVX3 U142 ( .A(n7409), .Y(n7563) );
  CLKINVX3 U143 ( .A(n7410), .Y(n7559) );
  CLKINVX3 U144 ( .A(n7410), .Y(n7560) );
  CLKINVX3 U145 ( .A(n7409), .Y(n7561) );
  CLKINVX3 U146 ( .A(n7402), .Y(n7589) );
  CLKINVX3 U147 ( .A(n7402), .Y(n7590) );
  CLKINVX3 U148 ( .A(n7398), .Y(n7586) );
  CLKINVX3 U149 ( .A(n7402), .Y(n7588) );
  CLKINVX3 U150 ( .A(n7402), .Y(n7587) );
  CLKINVX3 U151 ( .A(n7400), .Y(n7594) );
  CLKINVX3 U152 ( .A(n7400), .Y(n7595) );
  CLKINVX3 U153 ( .A(n7401), .Y(n7591) );
  CLKINVX3 U154 ( .A(n7401), .Y(n7592) );
  CLKINVX3 U155 ( .A(n7401), .Y(n7593) );
  CLKINVX3 U156 ( .A(n7404), .Y(n7578) );
  CLKINVX3 U157 ( .A(n7404), .Y(n7579) );
  CLKINVX3 U158 ( .A(n7405), .Y(n7575) );
  CLKINVX3 U159 ( .A(n7404), .Y(n7576) );
  CLKINVX3 U160 ( .A(n7404), .Y(n7577) );
  CLKINVX3 U161 ( .A(n7403), .Y(n7584) );
  CLKINVX3 U162 ( .A(n7403), .Y(n7585) );
  CLKINVX3 U163 ( .A(n7405), .Y(n7580) );
  CLKINVX3 U164 ( .A(n7411), .Y(n7581) );
  CLKINVX3 U165 ( .A(n7403), .Y(n7583) );
  CLKINVX3 U166 ( .A(n7403), .Y(n7582) );
  CLKINVX3 U167 ( .A(n7404), .Y(n7608) );
  CLKINVX3 U168 ( .A(n7398), .Y(n7600) );
  CLKINVX3 U169 ( .A(n7398), .Y(n7601) );
  CLKINVX3 U170 ( .A(n7400), .Y(n7596) );
  CLKINVX3 U171 ( .A(n7399), .Y(n7597) );
  CLKINVX3 U172 ( .A(n7399), .Y(n7599) );
  CLKINVX3 U173 ( .A(n7399), .Y(n7598) );
  CLKINVX3 U174 ( .A(n7410), .Y(n7605) );
  CLKINVX3 U175 ( .A(n7405), .Y(n7607) );
  CLKINVX3 U176 ( .A(n7408), .Y(n7606) );
  CLKINVX3 U177 ( .A(n7398), .Y(n7602) );
  CLKINVX3 U178 ( .A(n7407), .Y(n7604) );
  CLKINVX3 U179 ( .A(n7406), .Y(n7603) );
  CLKINVX3 U180 ( .A(n7687), .Y(n7703) );
  CLKINVX3 U181 ( .A(n7687), .Y(n7704) );
  CLKINVX3 U182 ( .A(n7687), .Y(n7702) );
  CLKINVX3 U183 ( .A(n7688), .Y(n7701) );
  CLKINVX3 U184 ( .A(n7685), .Y(n7708) );
  CLKINVX3 U185 ( .A(n7685), .Y(n7709) );
  CLKINVX3 U186 ( .A(n7686), .Y(n7705) );
  CLKINVX3 U187 ( .A(n7686), .Y(n7707) );
  CLKINVX3 U188 ( .A(n7686), .Y(n7706) );
  CLKINVX3 U189 ( .A(n7690), .Y(n7693) );
  CLKINVX3 U190 ( .A(n7690), .Y(n7694) );
  CLKINVX3 U191 ( .A(n7653), .Y(n7691) );
  CLKINVX3 U192 ( .A(n7652), .Y(n7692) );
  CLKINVX3 U193 ( .A(n7689), .Y(n7698) );
  CLKINVX3 U194 ( .A(n7688), .Y(n7700) );
  CLKINVX3 U195 ( .A(n7688), .Y(n7699) );
  CLKINVX3 U196 ( .A(n7690), .Y(n7695) );
  CLKINVX3 U197 ( .A(n7689), .Y(n7696) );
  CLKINVX3 U198 ( .A(n7689), .Y(n7697) );
  CLKINVX3 U199 ( .A(n7680), .Y(n7723) );
  CLKINVX3 U200 ( .A(n7681), .Y(n7720) );
  CLKINVX3 U201 ( .A(n7681), .Y(n7722) );
  CLKINVX3 U202 ( .A(n7681), .Y(n7721) );
  CLKINVX3 U203 ( .A(n7679), .Y(n7728) );
  CLKINVX3 U204 ( .A(n7680), .Y(n7724) );
  CLKINVX3 U205 ( .A(n7680), .Y(n7725) );
  CLKINVX3 U206 ( .A(n7679), .Y(n7727) );
  CLKINVX3 U207 ( .A(n7679), .Y(n7726) );
  CLKINVX3 U208 ( .A(n7684), .Y(n7713) );
  CLKINVX3 U209 ( .A(n7683), .Y(n7714) );
  CLKINVX3 U210 ( .A(n7685), .Y(n7710) );
  CLKINVX3 U211 ( .A(n7684), .Y(n7712) );
  CLKINVX3 U212 ( .A(n7684), .Y(n7711) );
  CLKINVX3 U213 ( .A(n7682), .Y(n7718) );
  CLKINVX3 U214 ( .A(n7682), .Y(n7719) );
  CLKINVX3 U215 ( .A(n7683), .Y(n7715) );
  CLKINVX3 U216 ( .A(n7682), .Y(n7717) );
  CLKINVX3 U217 ( .A(n7683), .Y(n7716) );
  CLKINVX3 U218 ( .A(n7674), .Y(n7743) );
  CLKINVX3 U219 ( .A(n7674), .Y(n7742) );
  CLKINVX3 U220 ( .A(n7675), .Y(n7740) );
  CLKINVX3 U221 ( .A(n7674), .Y(n7741) );
  CLKINVX3 U222 ( .A(n7672), .Y(n7748) );
  CLKINVX3 U223 ( .A(n7673), .Y(n7744) );
  CLKINVX3 U224 ( .A(n7672), .Y(n7747) );
  CLKINVX3 U225 ( .A(n7673), .Y(n7745) );
  CLKINVX3 U226 ( .A(n7673), .Y(n7746) );
  CLKINVX3 U227 ( .A(n7677), .Y(n7733) );
  CLKINVX3 U228 ( .A(n7678), .Y(n7729) );
  CLKINVX3 U229 ( .A(n7678), .Y(n7730) );
  CLKINVX3 U230 ( .A(n7677), .Y(n7732) );
  CLKINVX3 U231 ( .A(n7678), .Y(n7731) );
  CLKINVX3 U232 ( .A(n7675), .Y(n7739) );
  CLKINVX3 U233 ( .A(n7675), .Y(n7738) );
  CLKINVX3 U234 ( .A(n7677), .Y(n7734) );
  CLKINVX3 U235 ( .A(n7676), .Y(n7735) );
  CLKINVX3 U236 ( .A(n7676), .Y(n7737) );
  CLKINVX3 U237 ( .A(n7676), .Y(n7736) );
  CLKINVX3 U238 ( .A(n7667), .Y(n7762) );
  CLKINVX3 U239 ( .A(n7667), .Y(n7763) );
  CLKINVX3 U240 ( .A(n7668), .Y(n7760) );
  CLKINVX3 U241 ( .A(n7668), .Y(n7761) );
  CLKINVX3 U242 ( .A(n7666), .Y(n7767) );
  CLKINVX3 U243 ( .A(n7665), .Y(n7768) );
  CLKINVX3 U244 ( .A(n7667), .Y(n7764) );
  CLKINVX3 U245 ( .A(n7666), .Y(n7766) );
  CLKINVX3 U246 ( .A(n7666), .Y(n7765) );
  CLKINVX3 U247 ( .A(n7671), .Y(n7752) );
  CLKINVX3 U248 ( .A(n7670), .Y(n7753) );
  CLKINVX3 U249 ( .A(n7672), .Y(n7749) );
  CLKINVX3 U250 ( .A(n7671), .Y(n7750) );
  CLKINVX3 U251 ( .A(n7671), .Y(n7751) );
  CLKINVX3 U252 ( .A(n7669), .Y(n7757) );
  CLKINVX3 U253 ( .A(n7668), .Y(n7759) );
  CLKINVX3 U254 ( .A(n7669), .Y(n7758) );
  CLKINVX3 U255 ( .A(n7670), .Y(n7754) );
  CLKINVX3 U256 ( .A(n7670), .Y(n7755) );
  CLKINVX3 U257 ( .A(n7669), .Y(n7756) );
  CLKINVX3 U258 ( .A(n7661), .Y(n7782) );
  CLKINVX3 U259 ( .A(n7660), .Y(n7783) );
  CLKINVX3 U260 ( .A(n7661), .Y(n7781) );
  CLKINVX3 U261 ( .A(n7661), .Y(n7780) );
  CLKINVX3 U262 ( .A(n7659), .Y(n7787) );
  CLKINVX3 U263 ( .A(n7660), .Y(n7784) );
  CLKINVX3 U264 ( .A(n7659), .Y(n7786) );
  CLKINVX3 U265 ( .A(n7660), .Y(n7785) );
  CLKINVX3 U266 ( .A(n7664), .Y(n7772) );
  CLKINVX3 U267 ( .A(n7664), .Y(n7773) );
  CLKINVX3 U268 ( .A(n7665), .Y(n7769) );
  CLKINVX3 U269 ( .A(n7664), .Y(n7771) );
  CLKINVX3 U270 ( .A(n7665), .Y(n7770) );
  CLKINVX3 U271 ( .A(n7662), .Y(n7779) );
  CLKINVX3 U272 ( .A(n7662), .Y(n7777) );
  CLKINVX3 U273 ( .A(n7662), .Y(n7778) );
  CLKINVX3 U274 ( .A(n7663), .Y(n7774) );
  CLKINVX3 U275 ( .A(n7663), .Y(n7776) );
  CLKINVX3 U276 ( .A(n7663), .Y(n7775) );
  CLKINVX3 U277 ( .A(n7657), .Y(n7792) );
  CLKINVX3 U278 ( .A(n7659), .Y(n7788) );
  CLKINVX3 U279 ( .A(n7658), .Y(n7789) );
  CLKINVX3 U280 ( .A(n7658), .Y(n7791) );
  CLKINVX3 U281 ( .A(n7658), .Y(n7790) );
  CLKINVX3 U282 ( .A(n7657), .Y(n7793) );
  CLKINVX3 U283 ( .A(n7657), .Y(n7794) );
  CLKINVX3 U284 ( .A(n4100), .Y(n4118) );
  CLKINVX3 U285 ( .A(n4099), .Y(n4119) );
  CLKINVX3 U286 ( .A(n4101), .Y(n4115) );
  CLKINVX3 U287 ( .A(n4100), .Y(n4117) );
  CLKINVX3 U288 ( .A(n4100), .Y(n4116) );
  CLKINVX3 U289 ( .A(n4098), .Y(n4123) );
  CLKINVX3 U290 ( .A(n4098), .Y(n4124) );
  CLKINVX3 U291 ( .A(n4099), .Y(n4120) );
  CLKINVX3 U292 ( .A(n4099), .Y(n4121) );
  CLKINVX3 U293 ( .A(n4098), .Y(n4122) );
  CLKINVX3 U294 ( .A(n4103), .Y(n4107) );
  CLKINVX3 U295 ( .A(n4103), .Y(n4108) );
  CLKINVX3 U296 ( .A(n4104), .Y(n4105) );
  CLKINVX3 U297 ( .A(n4104), .Y(n4106) );
  CLKINVX3 U298 ( .A(n4101), .Y(n4113) );
  CLKINVX3 U299 ( .A(n4101), .Y(n4114) );
  CLKINVX3 U300 ( .A(n4103), .Y(n4109) );
  CLKINVX3 U301 ( .A(n4102), .Y(n4110) );
  CLKINVX3 U302 ( .A(n4102), .Y(n4112) );
  CLKINVX3 U303 ( .A(n4102), .Y(n4111) );
  CLKINVX3 U304 ( .A(n4093), .Y(n4139) );
  CLKINVX3 U305 ( .A(n4092), .Y(n4140) );
  CLKINVX3 U306 ( .A(n4093), .Y(n4137) );
  CLKINVX3 U307 ( .A(n4093), .Y(n4138) );
  CLKINVX3 U308 ( .A(n4091), .Y(n4145) );
  CLKINVX3 U309 ( .A(n4090), .Y(n4146) );
  CLKINVX3 U310 ( .A(n4092), .Y(n4141) );
  CLKINVX3 U311 ( .A(n4092), .Y(n4142) );
  CLKINVX3 U312 ( .A(n4091), .Y(n4144) );
  CLKINVX3 U313 ( .A(n4091), .Y(n4143) );
  CLKINVX3 U314 ( .A(n4096), .Y(n4129) );
  CLKINVX3 U315 ( .A(n4096), .Y(n4130) );
  CLKINVX3 U316 ( .A(n4097), .Y(n4125) );
  CLKINVX3 U317 ( .A(n4097), .Y(n4126) );
  CLKINVX3 U318 ( .A(n4096), .Y(n4128) );
  CLKINVX3 U319 ( .A(n4097), .Y(n4127) );
  CLKINVX3 U320 ( .A(n4094), .Y(n4134) );
  CLKINVX3 U321 ( .A(n4094), .Y(n4136) );
  CLKINVX3 U322 ( .A(n4094), .Y(n4135) );
  CLKINVX3 U323 ( .A(n4095), .Y(n4131) );
  CLKINVX3 U324 ( .A(n4095), .Y(n4133) );
  CLKINVX3 U325 ( .A(n4095), .Y(n4132) );
  CLKINVX3 U326 ( .A(n4085), .Y(n4161) );
  CLKINVX3 U327 ( .A(n4085), .Y(n4162) );
  CLKINVX3 U328 ( .A(n4086), .Y(n4158) );
  CLKINVX3 U329 ( .A(n4086), .Y(n4160) );
  CLKINVX3 U330 ( .A(n4086), .Y(n4159) );
  CLKINVX3 U331 ( .A(n4084), .Y(n4166) );
  CLKINVX3 U332 ( .A(n4083), .Y(n4167) );
  CLKINVX3 U333 ( .A(n4085), .Y(n4163) );
  CLKINVX3 U334 ( .A(n4084), .Y(n4165) );
  CLKINVX3 U335 ( .A(n4084), .Y(n4164) );
  CLKINVX3 U336 ( .A(n4089), .Y(n4150) );
  CLKINVX3 U337 ( .A(n4089), .Y(n4151) );
  CLKINVX3 U338 ( .A(n4090), .Y(n4147) );
  CLKINVX3 U339 ( .A(n4089), .Y(n4149) );
  CLKINVX3 U340 ( .A(n4090), .Y(n4148) );
  CLKINVX3 U341 ( .A(n4087), .Y(n4155) );
  CLKINVX3 U342 ( .A(n4087), .Y(n4157) );
  CLKINVX3 U343 ( .A(n4087), .Y(n4156) );
  CLKINVX3 U344 ( .A(n4088), .Y(n4152) );
  CLKINVX3 U345 ( .A(n4088), .Y(n4153) );
  CLKINVX3 U346 ( .A(n4088), .Y(n4154) );
  CLKINVX3 U347 ( .A(n4078), .Y(n4182) );
  CLKINVX3 U348 ( .A(n4078), .Y(n4183) );
  CLKINVX3 U349 ( .A(n4079), .Y(n4179) );
  CLKINVX3 U350 ( .A(n4079), .Y(n4181) );
  CLKINVX3 U351 ( .A(n4079), .Y(n4180) );
  CLKINVX3 U352 ( .A(n4077), .Y(n4187) );
  CLKINVX3 U353 ( .A(n4076), .Y(n4188) );
  CLKINVX3 U354 ( .A(n4078), .Y(n4184) );
  CLKINVX3 U355 ( .A(n4077), .Y(n4185) );
  CLKINVX3 U356 ( .A(n4077), .Y(n4186) );
  CLKINVX3 U357 ( .A(n4082), .Y(n4171) );
  CLKINVX3 U358 ( .A(n4082), .Y(n4172) );
  CLKINVX3 U359 ( .A(n4083), .Y(n4168) );
  CLKINVX3 U360 ( .A(n4083), .Y(n4169) );
  CLKINVX3 U361 ( .A(n4082), .Y(n4170) );
  CLKINVX3 U362 ( .A(n4080), .Y(n4177) );
  CLKINVX3 U363 ( .A(n4080), .Y(n4178) );
  CLKINVX3 U364 ( .A(n4081), .Y(n4173) );
  CLKINVX3 U365 ( .A(n4081), .Y(n4174) );
  CLKINVX3 U366 ( .A(n4080), .Y(n4176) );
  CLKINVX3 U367 ( .A(n4081), .Y(n4175) );
  CLKINVX3 U368 ( .A(n4071), .Y(n4203) );
  CLKINVX3 U369 ( .A(n4071), .Y(n4204) );
  CLKINVX3 U370 ( .A(n4072), .Y(n4201) );
  CLKINVX3 U371 ( .A(n4072), .Y(n4202) );
  CLKINVX3 U372 ( .A(n4069), .Y(n4209) );
  CLKINVX3 U373 ( .A(n4069), .Y(n4210) );
  CLKINVX3 U374 ( .A(n4071), .Y(n4205) );
  CLKINVX3 U375 ( .A(n4070), .Y(n4206) );
  CLKINVX3 U376 ( .A(n4070), .Y(n4208) );
  CLKINVX3 U377 ( .A(n4070), .Y(n4207) );
  CLKINVX3 U378 ( .A(n4075), .Y(n4193) );
  CLKINVX3 U379 ( .A(n4074), .Y(n4194) );
  CLKINVX3 U380 ( .A(n4076), .Y(n4189) );
  CLKINVX3 U381 ( .A(n4076), .Y(n4190) );
  CLKINVX3 U382 ( .A(n4075), .Y(n4192) );
  CLKINVX3 U383 ( .A(n4075), .Y(n4191) );
  CLKINVX3 U384 ( .A(n4073), .Y(n4198) );
  CLKINVX3 U385 ( .A(n4072), .Y(n4200) );
  CLKINVX3 U386 ( .A(n4073), .Y(n4199) );
  CLKINVX3 U387 ( .A(n4074), .Y(n4195) );
  CLKINVX3 U388 ( .A(n4073), .Y(n4197) );
  CLKINVX3 U389 ( .A(n4074), .Y(n4196) );
  CLKINVX3 U390 ( .A(n4065), .Y(n4225) );
  CLKINVX3 U391 ( .A(n4065), .Y(n4226) );
  CLKINVX3 U392 ( .A(n4064), .Y(n4222) );
  CLKINVX3 U393 ( .A(n4065), .Y(n4224) );
  CLKINVX3 U394 ( .A(n4049), .Y(n4223) );
  CLKINVX3 U395 ( .A(n4063), .Y(n4230) );
  CLKINVX3 U396 ( .A(n4063), .Y(n4231) );
  CLKINVX3 U397 ( .A(n4064), .Y(n4227) );
  CLKINVX3 U398 ( .A(n4064), .Y(n4229) );
  CLKINVX3 U399 ( .A(n4064), .Y(n4228) );
  CLKINVX3 U400 ( .A(n4068), .Y(n4214) );
  CLKINVX3 U401 ( .A(n4067), .Y(n4215) );
  CLKINVX3 U402 ( .A(n4069), .Y(n4211) );
  CLKINVX3 U403 ( .A(n4068), .Y(n4213) );
  CLKINVX3 U404 ( .A(n4068), .Y(n4212) );
  CLKINVX3 U405 ( .A(n4066), .Y(n4219) );
  CLKINVX3 U406 ( .A(n4065), .Y(n4221) );
  CLKINVX3 U407 ( .A(n4066), .Y(n4220) );
  CLKINVX3 U408 ( .A(n4067), .Y(n4216) );
  CLKINVX3 U409 ( .A(n4067), .Y(n4217) );
  CLKINVX3 U410 ( .A(n4066), .Y(n4218) );
  CLKINVX3 U411 ( .A(n4058), .Y(n4246) );
  CLKINVX3 U412 ( .A(n4058), .Y(n4247) );
  CLKINVX3 U413 ( .A(n4059), .Y(n4243) );
  CLKINVX3 U414 ( .A(n4058), .Y(n4245) );
  CLKINVX3 U415 ( .A(n4059), .Y(n4244) );
  CLKINVX3 U416 ( .A(n4056), .Y(n4251) );
  CLKINVX3 U417 ( .A(n4056), .Y(n4252) );
  CLKINVX3 U418 ( .A(n4057), .Y(n4248) );
  CLKINVX3 U419 ( .A(n4057), .Y(n4249) );
  CLKINVX3 U420 ( .A(n4057), .Y(n4250) );
  CLKINVX3 U421 ( .A(n4062), .Y(n4235) );
  CLKINVX3 U422 ( .A(n4061), .Y(n4236) );
  CLKINVX3 U423 ( .A(n4063), .Y(n4232) );
  CLKINVX3 U424 ( .A(n4062), .Y(n4233) );
  CLKINVX3 U425 ( .A(n4062), .Y(n4234) );
  CLKINVX3 U426 ( .A(n4060), .Y(n4241) );
  CLKINVX3 U427 ( .A(n4059), .Y(n4242) );
  CLKINVX3 U428 ( .A(n4061), .Y(n4237) );
  CLKINVX3 U429 ( .A(n4061), .Y(n4238) );
  CLKINVX3 U430 ( .A(n4060), .Y(n4240) );
  CLKINVX3 U431 ( .A(n4060), .Y(n4239) );
  CLKINVX3 U432 ( .A(n4052), .Y(n4265) );
  CLKINVX3 U433 ( .A(n4054), .Y(n4257) );
  CLKINVX3 U434 ( .A(n4054), .Y(n4258) );
  CLKINVX3 U435 ( .A(n4056), .Y(n4253) );
  CLKINVX3 U436 ( .A(n4055), .Y(n4254) );
  CLKINVX3 U437 ( .A(n4055), .Y(n4256) );
  CLKINVX3 U438 ( .A(n4055), .Y(n4255) );
  CLKINVX3 U439 ( .A(n4053), .Y(n4262) );
  CLKINVX3 U440 ( .A(n4052), .Y(n4264) );
  CLKINVX3 U441 ( .A(n4052), .Y(n4263) );
  CLKINVX3 U442 ( .A(n4054), .Y(n4259) );
  CLKINVX3 U443 ( .A(n4053), .Y(n4261) );
  CLKINVX3 U444 ( .A(n4053), .Y(n4260) );
  CLKINVX3 U445 ( .A(n7400), .Y(n7610) );
  CLKINVX3 U446 ( .A(n7401), .Y(n7609) );
  CLKINVX3 U447 ( .A(n7399), .Y(n7611) );
  CLKINVX3 U448 ( .A(n7397), .Y(n7612) );
  CLKINVX3 U449 ( .A(n7397), .Y(n7613) );
  CLKINVX3 U450 ( .A(n7396), .Y(n7616) );
  CLKINVX3 U451 ( .A(n7396), .Y(n7617) );
  CLKINVX3 U452 ( .A(n7396), .Y(n7615) );
  CLKINVX3 U453 ( .A(n7397), .Y(n7614) );
  CLKINVX3 U454 ( .A(n4345), .Y(n4359) );
  CLKINVX3 U455 ( .A(n4345), .Y(n4360) );
  CLKINVX3 U456 ( .A(n4345), .Y(n4358) );
  CLKINVX3 U457 ( .A(n4346), .Y(n4357) );
  CLKINVX3 U458 ( .A(n4343), .Y(n4364) );
  CLKINVX3 U459 ( .A(n4343), .Y(n4365) );
  CLKINVX3 U460 ( .A(n4344), .Y(n4361) );
  CLKINVX3 U461 ( .A(n4344), .Y(n4363) );
  CLKINVX3 U462 ( .A(n4344), .Y(n4362) );
  CLKINVX3 U463 ( .A(n4348), .Y(n4349) );
  CLKINVX3 U464 ( .A(n4348), .Y(n4350) );
  CLKINVX3 U465 ( .A(n4347), .Y(n4354) );
  CLKINVX3 U466 ( .A(n4346), .Y(n4356) );
  CLKINVX3 U467 ( .A(n4346), .Y(n4355) );
  CLKINVX3 U468 ( .A(n4337), .Y(n4351) );
  CLKINVX3 U469 ( .A(n4347), .Y(n4352) );
  CLKINVX3 U470 ( .A(n4347), .Y(n4353) );
  CLKINVX3 U471 ( .A(n4338), .Y(n4379) );
  CLKINVX3 U472 ( .A(n4339), .Y(n4376) );
  CLKINVX3 U473 ( .A(n4339), .Y(n4378) );
  CLKINVX3 U474 ( .A(n4339), .Y(n4377) );
  CLKINVX3 U475 ( .A(n4337), .Y(n4384) );
  CLKINVX3 U476 ( .A(n4338), .Y(n4380) );
  CLKINVX3 U477 ( .A(n4338), .Y(n4381) );
  CLKINVX3 U478 ( .A(n4337), .Y(n4383) );
  CLKINVX3 U479 ( .A(n4337), .Y(n4382) );
  CLKINVX3 U480 ( .A(n4342), .Y(n4369) );
  CLKINVX3 U481 ( .A(n4341), .Y(n4370) );
  CLKINVX3 U482 ( .A(n4343), .Y(n4366) );
  CLKINVX3 U483 ( .A(n4342), .Y(n4368) );
  CLKINVX3 U484 ( .A(n4342), .Y(n4367) );
  CLKINVX3 U485 ( .A(n4340), .Y(n4374) );
  CLKINVX3 U486 ( .A(n4340), .Y(n4375) );
  CLKINVX3 U487 ( .A(n4341), .Y(n4371) );
  CLKINVX3 U488 ( .A(n4340), .Y(n4373) );
  CLKINVX3 U489 ( .A(n4341), .Y(n4372) );
  CLKINVX3 U490 ( .A(n4332), .Y(n4399) );
  CLKINVX3 U491 ( .A(n4332), .Y(n4398) );
  CLKINVX3 U492 ( .A(n4333), .Y(n4396) );
  CLKINVX3 U493 ( .A(n4332), .Y(n4397) );
  CLKINVX3 U494 ( .A(n4330), .Y(n4404) );
  CLKINVX3 U495 ( .A(n4331), .Y(n4400) );
  CLKINVX3 U496 ( .A(n4330), .Y(n4403) );
  CLKINVX3 U497 ( .A(n4331), .Y(n4401) );
  CLKINVX3 U498 ( .A(n4331), .Y(n4402) );
  CLKINVX3 U499 ( .A(n4335), .Y(n4389) );
  CLKINVX3 U500 ( .A(n4336), .Y(n4385) );
  CLKINVX3 U501 ( .A(n4336), .Y(n4386) );
  CLKINVX3 U502 ( .A(n4335), .Y(n4388) );
  CLKINVX3 U503 ( .A(n4336), .Y(n4387) );
  CLKINVX3 U504 ( .A(n4333), .Y(n4395) );
  CLKINVX3 U505 ( .A(n4333), .Y(n4394) );
  CLKINVX3 U506 ( .A(n4335), .Y(n4390) );
  CLKINVX3 U507 ( .A(n4334), .Y(n4391) );
  CLKINVX3 U508 ( .A(n4334), .Y(n4393) );
  CLKINVX3 U509 ( .A(n4334), .Y(n4392) );
  CLKINVX3 U510 ( .A(n4325), .Y(n4418) );
  CLKINVX3 U511 ( .A(n4325), .Y(n4419) );
  CLKINVX3 U512 ( .A(n4326), .Y(n4416) );
  CLKINVX3 U513 ( .A(n4326), .Y(n4417) );
  CLKINVX3 U514 ( .A(n4324), .Y(n4423) );
  CLKINVX3 U515 ( .A(n4323), .Y(n4424) );
  CLKINVX3 U516 ( .A(n4325), .Y(n4420) );
  CLKINVX3 U517 ( .A(n4324), .Y(n4422) );
  CLKINVX3 U518 ( .A(n4324), .Y(n4421) );
  CLKINVX3 U519 ( .A(n4329), .Y(n4408) );
  CLKINVX3 U520 ( .A(n4328), .Y(n4409) );
  CLKINVX3 U521 ( .A(n4330), .Y(n4405) );
  CLKINVX3 U522 ( .A(n4329), .Y(n4406) );
  CLKINVX3 U523 ( .A(n4329), .Y(n4407) );
  CLKINVX3 U524 ( .A(n4327), .Y(n4413) );
  CLKINVX3 U525 ( .A(n4326), .Y(n4415) );
  CLKINVX3 U526 ( .A(n4327), .Y(n4414) );
  CLKINVX3 U527 ( .A(n4328), .Y(n4410) );
  CLKINVX3 U528 ( .A(n4328), .Y(n4411) );
  CLKINVX3 U529 ( .A(n4327), .Y(n4412) );
  CLKINVX3 U530 ( .A(n4319), .Y(n4438) );
  CLKINVX3 U531 ( .A(n4318), .Y(n4439) );
  CLKINVX3 U532 ( .A(n4319), .Y(n4437) );
  CLKINVX3 U533 ( .A(n4319), .Y(n4436) );
  CLKINVX3 U534 ( .A(n4317), .Y(n4443) );
  CLKINVX3 U535 ( .A(n4318), .Y(n4440) );
  CLKINVX3 U536 ( .A(n4317), .Y(n4442) );
  CLKINVX3 U537 ( .A(n4318), .Y(n4441) );
  CLKINVX3 U538 ( .A(n4322), .Y(n4428) );
  CLKINVX3 U539 ( .A(n4322), .Y(n4429) );
  CLKINVX3 U540 ( .A(n4323), .Y(n4425) );
  CLKINVX3 U541 ( .A(n4322), .Y(n4427) );
  CLKINVX3 U542 ( .A(n4323), .Y(n4426) );
  CLKINVX3 U543 ( .A(n4320), .Y(n4435) );
  CLKINVX3 U544 ( .A(n4320), .Y(n4433) );
  CLKINVX3 U545 ( .A(n4320), .Y(n4434) );
  CLKINVX3 U546 ( .A(n4321), .Y(n4430) );
  CLKINVX3 U547 ( .A(n4321), .Y(n4432) );
  CLKINVX3 U548 ( .A(n4321), .Y(n4431) );
  CLKINVX3 U549 ( .A(n4315), .Y(n4448) );
  CLKINVX3 U550 ( .A(n4317), .Y(n4444) );
  CLKINVX3 U551 ( .A(n4316), .Y(n4445) );
  CLKINVX3 U552 ( .A(n4316), .Y(n4447) );
  CLKINVX3 U553 ( .A(n4316), .Y(n4446) );
  CLKINVX3 U554 ( .A(n4315), .Y(n4449) );
  CLKINVX3 U555 ( .A(n4315), .Y(n4450) );
  CLKINVX3 U556 ( .A(n7654), .Y(n7802) );
  CLKINVX3 U557 ( .A(n7655), .Y(n7799) );
  CLKINVX3 U558 ( .A(n7654), .Y(n7801) );
  CLKINVX3 U559 ( .A(n7655), .Y(n7800) );
  CLKINVX3 U560 ( .A(n7653), .Y(n7806) );
  CLKINVX3 U561 ( .A(n7654), .Y(n7803) );
  CLKINVX3 U562 ( .A(n7653), .Y(n7805) );
  CLKINVX3 U563 ( .A(n7652), .Y(n7804) );
  CLKINVX3 U564 ( .A(n7655), .Y(n7798) );
  CLKINVX3 U565 ( .A(n7656), .Y(n7797) );
  CLKINVX3 U566 ( .A(n7656), .Y(n7796) );
  CLKINVX3 U567 ( .A(n7656), .Y(n7795) );
  CLKINVX3 U568 ( .A(n7649), .Y(n7820) );
  CLKINVX3 U569 ( .A(n7648), .Y(n7821) );
  CLKINVX3 U570 ( .A(n7649), .Y(n7818) );
  CLKINVX3 U571 ( .A(n7649), .Y(n7819) );
  CLKINVX3 U572 ( .A(n7647), .Y(n7825) );
  CLKINVX3 U573 ( .A(n7647), .Y(n7826) );
  CLKINVX3 U574 ( .A(n7648), .Y(n7822) );
  CLKINVX3 U575 ( .A(n7648), .Y(n7823) );
  CLKINVX3 U576 ( .A(n7647), .Y(n7824) );
  CLKINVX3 U577 ( .A(n7652), .Y(n7811) );
  CLKINVX3 U578 ( .A(n7653), .Y(n7807) );
  CLKINVX3 U579 ( .A(n7652), .Y(n7810) );
  CLKINVX3 U580 ( .A(n7653), .Y(n7808) );
  CLKINVX3 U581 ( .A(n7652), .Y(n7809) );
  CLKINVX3 U582 ( .A(n7650), .Y(n7815) );
  CLKINVX3 U583 ( .A(n7650), .Y(n7817) );
  CLKINVX3 U584 ( .A(n7650), .Y(n7816) );
  CLKINVX3 U585 ( .A(n7651), .Y(n7812) );
  CLKINVX3 U586 ( .A(n7651), .Y(n7813) );
  CLKINVX3 U587 ( .A(n7651), .Y(n7814) );
  CLKINVX3 U588 ( .A(n7643), .Y(n7839) );
  CLKINVX3 U589 ( .A(n7651), .Y(n7838) );
  CLKINVX3 U590 ( .A(n7643), .Y(n7840) );
  CLKINVX3 U591 ( .A(n7643), .Y(n7841) );
  CLKINVX3 U592 ( .A(n7642), .Y(n7842) );
  CLKINVX3 U593 ( .A(n7643), .Y(n7845) );
  CLKINVX3 U594 ( .A(n7642), .Y(n7846) );
  CLKINVX3 U595 ( .A(n7642), .Y(n7844) );
  CLKINVX3 U596 ( .A(n7642), .Y(n7843) );
  CLKINVX3 U597 ( .A(n7645), .Y(n7830) );
  CLKINVX3 U598 ( .A(n7645), .Y(n7831) );
  CLKINVX3 U599 ( .A(n7646), .Y(n7827) );
  CLKINVX3 U600 ( .A(n7646), .Y(n7829) );
  CLKINVX3 U601 ( .A(n7646), .Y(n7828) );
  CLKINVX3 U602 ( .A(n7650), .Y(n7837) );
  CLKINVX3 U603 ( .A(n7644), .Y(n7835) );
  CLKINVX3 U604 ( .A(n7646), .Y(n7836) );
  CLKINVX3 U605 ( .A(n7645), .Y(n7832) );
  CLKINVX3 U606 ( .A(n7644), .Y(n7834) );
  CLKINVX3 U607 ( .A(n7644), .Y(n7833) );
  INVX1 U608 ( .A(n7628), .Y(n7687) );
  INVX1 U609 ( .A(n7382), .Y(n7443) );
  INVX1 U610 ( .A(n7382), .Y(n7442) );
  INVX1 U611 ( .A(n7383), .Y(n7441) );
  INVX1 U612 ( .A(n7629), .Y(n7686) );
  INVX1 U613 ( .A(n7382), .Y(n7444) );
  INVX1 U614 ( .A(n7628), .Y(n7688) );
  INVX1 U615 ( .A(n7381), .Y(n7446) );
  INVX1 U616 ( .A(n7381), .Y(n7445) );
  INVX1 U617 ( .A(n7628), .Y(n7689) );
  INVX1 U618 ( .A(n7384), .Y(n7436) );
  INVX1 U619 ( .A(n7630), .Y(n7681) );
  INVX1 U620 ( .A(n7385), .Y(n7435) );
  INVX1 U621 ( .A(n7631), .Y(n7680) );
  INVX1 U622 ( .A(n7385), .Y(n7434) );
  INVX1 U623 ( .A(n7631), .Y(n7679) );
  INVX1 U624 ( .A(n7629), .Y(n7685) );
  INVX1 U625 ( .A(n7383), .Y(n7439) );
  INVX1 U626 ( .A(n7383), .Y(n7440) );
  INVX1 U627 ( .A(n7629), .Y(n7684) );
  INVX1 U628 ( .A(n7384), .Y(n7437) );
  INVX1 U629 ( .A(n7630), .Y(n7682) );
  INVX1 U630 ( .A(n7384), .Y(n7438) );
  INVX1 U631 ( .A(n7630), .Y(n7683) );
  INVX1 U632 ( .A(n7387), .Y(n7429) );
  INVX1 U633 ( .A(n7633), .Y(n7674) );
  INVX1 U634 ( .A(n7387), .Y(n7428) );
  INVX1 U635 ( .A(n7387), .Y(n7427) );
  INVX1 U636 ( .A(n7633), .Y(n7673) );
  INVX1 U637 ( .A(n7386), .Y(n7432) );
  INVX1 U638 ( .A(n7385), .Y(n7433) );
  INVX1 U639 ( .A(n7631), .Y(n7678) );
  INVX1 U640 ( .A(n7386), .Y(n7430) );
  INVX1 U641 ( .A(n7632), .Y(n7675) );
  INVX1 U642 ( .A(n7632), .Y(n7677) );
  INVX1 U643 ( .A(n7386), .Y(n7431) );
  INVX1 U644 ( .A(n7632), .Y(n7676) );
  INVX1 U645 ( .A(n7389), .Y(n7422) );
  INVX1 U646 ( .A(n7389), .Y(n7421) );
  INVX1 U647 ( .A(n7635), .Y(n7667) );
  INVX1 U648 ( .A(n7390), .Y(n7420) );
  INVX1 U649 ( .A(n7635), .Y(n7666) );
  INVX1 U650 ( .A(n7633), .Y(n7672) );
  INVX1 U651 ( .A(n7388), .Y(n7426) );
  INVX1 U652 ( .A(n7388), .Y(n7425) );
  INVX1 U653 ( .A(n7634), .Y(n7671) );
  INVX1 U654 ( .A(n7635), .Y(n7668) );
  INVX1 U655 ( .A(n7389), .Y(n7423) );
  INVX1 U656 ( .A(n7634), .Y(n7670) );
  INVX1 U657 ( .A(n7388), .Y(n7424) );
  INVX1 U658 ( .A(n7634), .Y(n7669) );
  INVX1 U659 ( .A(n7637), .Y(n7661) );
  INVX1 U660 ( .A(n7392), .Y(n7414) );
  INVX1 U661 ( .A(n7392), .Y(n7413) );
  INVX1 U662 ( .A(n7637), .Y(n7660) );
  INVX1 U663 ( .A(n7390), .Y(n7419) );
  INVX1 U664 ( .A(n7636), .Y(n7664) );
  INVX1 U665 ( .A(n7390), .Y(n7418) );
  INVX1 U666 ( .A(n7636), .Y(n7665) );
  INVX1 U667 ( .A(n7391), .Y(n7415) );
  INVX1 U668 ( .A(n7637), .Y(n7662) );
  INVX1 U669 ( .A(n7391), .Y(n7416) );
  INVX1 U670 ( .A(n7391), .Y(n7417) );
  INVX1 U671 ( .A(n7636), .Y(n7663) );
  INVX1 U672 ( .A(n7394), .Y(n7407) );
  INVX1 U673 ( .A(n7394), .Y(n7406) );
  INVX1 U674 ( .A(n7638), .Y(n7659) );
  INVX1 U675 ( .A(n7392), .Y(n7412) );
  INVX1 U676 ( .A(n7393), .Y(n7411) );
  INVX1 U677 ( .A(n7638), .Y(n7658) );
  INVX1 U678 ( .A(n7394), .Y(n7408) );
  INVX1 U679 ( .A(n7638), .Y(n7657) );
  INVX1 U680 ( .A(n7393), .Y(n7410) );
  INVX1 U681 ( .A(n7393), .Y(n7409) );
  INVX1 U682 ( .A(n7393), .Y(n7402) );
  INVX1 U683 ( .A(n7395), .Y(n7401) );
  INVX1 U684 ( .A(n7395), .Y(n7405) );
  INVX1 U685 ( .A(N78), .Y(n7404) );
  INVX1 U686 ( .A(n7394), .Y(n7403) );
  INVX1 U687 ( .A(n7395), .Y(n7400) );
  INVX1 U688 ( .A(n7395), .Y(n7399) );
  INVX1 U689 ( .A(n7395), .Y(n7398) );
  INVX1 U690 ( .A(n7639), .Y(n7690) );
  INVX1 U691 ( .A(n7381), .Y(n7447) );
  CLKINVX3 U692 ( .A(n4586), .Y(n4587) );
  CLKINVX3 U693 ( .A(n4586), .Y(n4592) );
  CLKINVX3 U694 ( .A(n4584), .Y(n4593) );
  CLKINVX3 U695 ( .A(n4586), .Y(n4588) );
  CLKINVX3 U696 ( .A(n4585), .Y(n4589) );
  CLKINVX3 U697 ( .A(n4584), .Y(n4591) );
  CLKINVX3 U698 ( .A(n4585), .Y(n4590) );
  CLKINVX3 U699 ( .A(n4582), .Y(n4597) );
  CLKINVX3 U700 ( .A(n4582), .Y(n4598) );
  CLKINVX3 U701 ( .A(n4584), .Y(n4594) );
  CLKINVX3 U702 ( .A(n4583), .Y(n4596) );
  CLKINVX3 U703 ( .A(n4583), .Y(n4595) );
  CLKINVX3 U704 ( .A(n4583), .Y(n4602) );
  CLKINVX3 U705 ( .A(n4580), .Y(n4603) );
  CLKINVX3 U706 ( .A(n4581), .Y(n4599) );
  CLKINVX3 U707 ( .A(n4581), .Y(n4600) );
  CLKINVX3 U708 ( .A(n4582), .Y(n4601) );
  CLKINVX3 U709 ( .A(n4578), .Y(n4608) );
  CLKINVX3 U710 ( .A(n4577), .Y(n4609) );
  CLKINVX3 U711 ( .A(n4580), .Y(n4604) );
  CLKINVX3 U712 ( .A(n4579), .Y(n4605) );
  CLKINVX3 U713 ( .A(n4578), .Y(n4607) );
  CLKINVX3 U714 ( .A(n4579), .Y(n4606) );
  CLKINVX3 U715 ( .A(n4575), .Y(n4613) );
  CLKINVX3 U716 ( .A(n4575), .Y(n4614) );
  CLKINVX3 U717 ( .A(n4577), .Y(n4610) );
  CLKINVX3 U718 ( .A(n4576), .Y(n4612) );
  CLKINVX3 U719 ( .A(n4576), .Y(n4611) );
  CLKINVX3 U720 ( .A(n4573), .Y(n4618) );
  CLKINVX3 U721 ( .A(n4572), .Y(n4619) );
  CLKINVX3 U722 ( .A(n4574), .Y(n4615) );
  CLKINVX3 U723 ( .A(n4574), .Y(n4616) );
  CLKINVX3 U724 ( .A(n4573), .Y(n4617) );
  CLKINVX3 U725 ( .A(n4570), .Y(n4624) );
  CLKINVX3 U726 ( .A(n4572), .Y(n4620) );
  CLKINVX3 U727 ( .A(n4571), .Y(n4621) );
  CLKINVX3 U728 ( .A(n4570), .Y(n4623) );
  CLKINVX3 U729 ( .A(n4571), .Y(n4622) );
  CLKINVX3 U730 ( .A(n7929), .Y(n7930) );
  CLKINVX3 U731 ( .A(n7927), .Y(n7935) );
  CLKINVX3 U732 ( .A(n7926), .Y(n7936) );
  CLKINVX3 U733 ( .A(n7929), .Y(n7931) );
  CLKINVX3 U734 ( .A(n7928), .Y(n7932) );
  CLKINVX3 U735 ( .A(n7927), .Y(n7934) );
  CLKINVX3 U736 ( .A(n7928), .Y(n7933) );
  CLKINVX3 U737 ( .A(n7924), .Y(n7940) );
  CLKINVX3 U738 ( .A(n7924), .Y(n7941) );
  CLKINVX3 U739 ( .A(n7926), .Y(n7937) );
  CLKINVX3 U740 ( .A(n7925), .Y(n7939) );
  CLKINVX3 U741 ( .A(n7925), .Y(n7938) );
  CLKINVX3 U742 ( .A(n7925), .Y(n7945) );
  CLKINVX3 U743 ( .A(n7922), .Y(n7946) );
  CLKINVX3 U744 ( .A(n7923), .Y(n7942) );
  CLKINVX3 U745 ( .A(n7923), .Y(n7943) );
  CLKINVX3 U746 ( .A(n7924), .Y(n7944) );
  CLKINVX3 U747 ( .A(n7920), .Y(n7951) );
  CLKINVX3 U748 ( .A(n7919), .Y(n7952) );
  CLKINVX3 U749 ( .A(n7922), .Y(n7947) );
  CLKINVX3 U750 ( .A(n7921), .Y(n7948) );
  CLKINVX3 U751 ( .A(n7920), .Y(n7950) );
  CLKINVX3 U752 ( .A(n7921), .Y(n7949) );
  CLKINVX3 U753 ( .A(n7917), .Y(n7956) );
  CLKINVX3 U754 ( .A(n7917), .Y(n7957) );
  CLKINVX3 U755 ( .A(n7919), .Y(n7953) );
  CLKINVX3 U756 ( .A(n7918), .Y(n7955) );
  CLKINVX3 U757 ( .A(n7918), .Y(n7954) );
  CLKINVX3 U758 ( .A(n7915), .Y(n7961) );
  CLKINVX3 U759 ( .A(n7914), .Y(n7962) );
  CLKINVX3 U760 ( .A(n7916), .Y(n7958) );
  CLKINVX3 U761 ( .A(n7916), .Y(n7959) );
  CLKINVX3 U762 ( .A(n7915), .Y(n7960) );
  CLKINVX3 U763 ( .A(n7912), .Y(n7967) );
  CLKINVX3 U764 ( .A(n7914), .Y(n7963) );
  CLKINVX3 U765 ( .A(n7913), .Y(n7964) );
  CLKINVX3 U766 ( .A(n7912), .Y(n7966) );
  CLKINVX3 U767 ( .A(n7913), .Y(n7965) );
  CLKINVX3 U768 ( .A(n4523), .Y(n4529) );
  CLKINVX3 U769 ( .A(n4524), .Y(n4528) );
  CLKINVX3 U770 ( .A(n4524), .Y(n4526) );
  CLKINVX3 U771 ( .A(n4524), .Y(n4527) );
  CLKINVX3 U772 ( .A(n4523), .Y(n4533) );
  CLKINVX3 U773 ( .A(n4522), .Y(n4534) );
  CLKINVX3 U774 ( .A(n4523), .Y(n4530) );
  CLKINVX3 U775 ( .A(n4522), .Y(n4531) );
  CLKINVX3 U776 ( .A(n4522), .Y(n4532) );
  CLKINVX3 U777 ( .A(n4520), .Y(n4538) );
  CLKINVX3 U778 ( .A(n4519), .Y(n4539) );
  CLKINVX3 U779 ( .A(n4521), .Y(n4535) );
  CLKINVX3 U780 ( .A(n4521), .Y(n4536) );
  CLKINVX3 U781 ( .A(n4520), .Y(n4537) );
  CLKINVX3 U782 ( .A(n4517), .Y(n4543) );
  CLKINVX3 U783 ( .A(n4519), .Y(n4540) );
  CLKINVX3 U784 ( .A(n4518), .Y(n4541) );
  CLKINVX3 U785 ( .A(n4518), .Y(n4542) );
  CLKINVX3 U786 ( .A(n4516), .Y(n4547) );
  CLKINVX3 U787 ( .A(n4515), .Y(n4548) );
  CLKINVX3 U788 ( .A(n4517), .Y(n4544) );
  CLKINVX3 U789 ( .A(n4516), .Y(n4546) );
  CLKINVX3 U790 ( .A(n4517), .Y(n4545) );
  CLKINVX3 U791 ( .A(n4513), .Y(n4552) );
  CLKINVX3 U792 ( .A(n4513), .Y(n4553) );
  CLKINVX3 U793 ( .A(n4515), .Y(n4549) );
  CLKINVX3 U794 ( .A(n4514), .Y(n4551) );
  CLKINVX3 U795 ( .A(n4514), .Y(n4550) );
  CLKINVX3 U796 ( .A(n4511), .Y(n4557) );
  CLKINVX3 U797 ( .A(n4512), .Y(n4554) );
  CLKINVX3 U798 ( .A(n4511), .Y(n4556) );
  CLKINVX3 U799 ( .A(n4512), .Y(n4555) );
  CLKINVX3 U800 ( .A(n7864), .Y(n7870) );
  CLKINVX3 U801 ( .A(n7865), .Y(n7869) );
  CLKINVX3 U802 ( .A(n7853), .Y(n7867) );
  CLKINVX3 U803 ( .A(n7865), .Y(n7868) );
  CLKINVX3 U804 ( .A(n7862), .Y(n7874) );
  CLKINVX3 U805 ( .A(n7862), .Y(n7875) );
  CLKINVX3 U806 ( .A(n7864), .Y(n7871) );
  CLKINVX3 U807 ( .A(n7863), .Y(n7872) );
  CLKINVX3 U808 ( .A(n7863), .Y(n7873) );
  CLKINVX3 U809 ( .A(n7860), .Y(n7879) );
  CLKINVX3 U810 ( .A(n7859), .Y(n7880) );
  CLKINVX3 U811 ( .A(n7861), .Y(n7876) );
  CLKINVX3 U812 ( .A(n7861), .Y(n7877) );
  CLKINVX3 U813 ( .A(n7860), .Y(n7878) );
  CLKINVX3 U814 ( .A(n7857), .Y(n7884) );
  CLKINVX3 U815 ( .A(n7857), .Y(n7885) );
  CLKINVX3 U816 ( .A(n7859), .Y(n7881) );
  CLKINVX3 U817 ( .A(n7858), .Y(n7882) );
  CLKINVX3 U818 ( .A(n7858), .Y(n7883) );
  CLKINVX3 U819 ( .A(n7855), .Y(n7889) );
  CLKINVX3 U820 ( .A(n7855), .Y(n7890) );
  CLKINVX3 U821 ( .A(n7856), .Y(n7886) );
  CLKINVX3 U822 ( .A(n7855), .Y(n7888) );
  CLKINVX3 U823 ( .A(n7856), .Y(n7887) );
  CLKINVX3 U824 ( .A(n7854), .Y(n7894) );
  CLKINVX3 U825 ( .A(n7853), .Y(n7895) );
  CLKINVX3 U826 ( .A(n7853), .Y(n7891) );
  CLKINVX3 U827 ( .A(n7855), .Y(n7893) );
  CLKINVX3 U828 ( .A(n7854), .Y(n7892) );
  CLKINVX3 U829 ( .A(n7854), .Y(n7897) );
  CLKINVX3 U830 ( .A(n7855), .Y(n7896) );
  INVX1 U831 ( .A(n4510), .Y(n4525) );
  INVX1 U832 ( .A(n7848), .Y(n7866) );
  CLKINVX3 U833 ( .A(n4051), .Y(n4267) );
  CLKINVX3 U834 ( .A(n4051), .Y(n4268) );
  CLKINVX3 U835 ( .A(n4051), .Y(n4266) );
  CLKINVX3 U836 ( .A(n4049), .Y(n4273) );
  CLKINVX3 U837 ( .A(n4049), .Y(n4274) );
  CLKINVX3 U838 ( .A(n4050), .Y(n4269) );
  CLKINVX3 U839 ( .A(n4050), .Y(n4270) );
  CLKINVX3 U840 ( .A(n4049), .Y(n4272) );
  CLKINVX3 U841 ( .A(n4050), .Y(n4271) );
  CLKINVX3 U842 ( .A(n4312), .Y(n4458) );
  CLKINVX3 U843 ( .A(n4313), .Y(n4455) );
  CLKINVX3 U844 ( .A(n4312), .Y(n4457) );
  CLKINVX3 U845 ( .A(n4313), .Y(n4456) );
  CLKINVX3 U846 ( .A(n4310), .Y(n4463) );
  CLKINVX3 U847 ( .A(n4312), .Y(n4459) );
  CLKINVX3 U848 ( .A(n4311), .Y(n4462) );
  CLKINVX3 U849 ( .A(n4311), .Y(n4460) );
  CLKINVX3 U850 ( .A(n4311), .Y(n4461) );
  CLKINVX3 U851 ( .A(n4313), .Y(n4454) );
  CLKINVX3 U852 ( .A(n4314), .Y(n4453) );
  CLKINVX3 U853 ( .A(n4314), .Y(n4452) );
  CLKINVX3 U854 ( .A(n4314), .Y(n4451) );
  CLKINVX3 U855 ( .A(n4312), .Y(n4477) );
  CLKINVX3 U856 ( .A(n4307), .Y(n4478) );
  CLKINVX3 U857 ( .A(n4314), .Y(n4475) );
  CLKINVX3 U858 ( .A(n4313), .Y(n4476) );
  CLKINVX3 U859 ( .A(n4306), .Y(n4482) );
  CLKINVX3 U860 ( .A(n4306), .Y(n4483) );
  CLKINVX3 U861 ( .A(n4307), .Y(n4479) );
  CLKINVX3 U862 ( .A(n4307), .Y(n4480) );
  CLKINVX3 U863 ( .A(n4306), .Y(n4481) );
  CLKINVX3 U864 ( .A(n4309), .Y(n4468) );
  CLKINVX3 U865 ( .A(n4310), .Y(n4464) );
  CLKINVX3 U866 ( .A(n4309), .Y(n4467) );
  CLKINVX3 U867 ( .A(n4310), .Y(n4465) );
  CLKINVX3 U868 ( .A(n4309), .Y(n4466) );
  CLKINVX3 U869 ( .A(n4311), .Y(n4472) );
  CLKINVX3 U870 ( .A(n4303), .Y(n4474) );
  CLKINVX3 U871 ( .A(n4308), .Y(n4473) );
  CLKINVX3 U872 ( .A(n4308), .Y(n4469) );
  CLKINVX3 U873 ( .A(n4308), .Y(n4470) );
  CLKINVX3 U874 ( .A(n4308), .Y(n4471) );
  CLKINVX3 U875 ( .A(n4302), .Y(n4497) );
  CLKINVX3 U876 ( .A(n4304), .Y(n4496) );
  CLKINVX3 U877 ( .A(n4302), .Y(n4495) );
  CLKINVX3 U878 ( .A(n4301), .Y(n4501) );
  CLKINVX3 U879 ( .A(n4301), .Y(n4498) );
  CLKINVX3 U880 ( .A(n4301), .Y(n4500) );
  CLKINVX3 U881 ( .A(n4301), .Y(n4499) );
  CLKINVX3 U882 ( .A(n4304), .Y(n4487) );
  CLKINVX3 U883 ( .A(n4304), .Y(n4488) );
  CLKINVX3 U884 ( .A(n4305), .Y(n4484) );
  CLKINVX3 U885 ( .A(n4305), .Y(n4486) );
  CLKINVX3 U886 ( .A(n4305), .Y(n4485) );
  CLKINVX3 U887 ( .A(n4302), .Y(n4494) );
  CLKINVX3 U888 ( .A(n4303), .Y(n4492) );
  CLKINVX3 U889 ( .A(n4302), .Y(n4493) );
  CLKINVX3 U890 ( .A(n4304), .Y(n4489) );
  CLKINVX3 U891 ( .A(n4303), .Y(n4491) );
  CLKINVX3 U892 ( .A(n4303), .Y(n4490) );
  INVX1 U893 ( .A(n4286), .Y(n4345) );
  INVX1 U894 ( .A(n4033), .Y(n4100) );
  INVX1 U895 ( .A(n4033), .Y(n4099) );
  INVX1 U896 ( .A(n4034), .Y(n4098) );
  INVX1 U897 ( .A(n4287), .Y(n4344) );
  INVX1 U898 ( .A(n4033), .Y(n4101) );
  INVX1 U899 ( .A(n4286), .Y(n4346) );
  INVX1 U900 ( .A(n4032), .Y(n4103) );
  INVX1 U901 ( .A(n4032), .Y(n4102) );
  INVX1 U902 ( .A(n4286), .Y(n4347) );
  INVX1 U903 ( .A(n4035), .Y(n4093) );
  INVX1 U904 ( .A(n4288), .Y(n4339) );
  INVX1 U905 ( .A(n4036), .Y(n4092) );
  INVX1 U906 ( .A(n4289), .Y(n4338) );
  INVX1 U907 ( .A(n4036), .Y(n4091) );
  INVX1 U908 ( .A(n4289), .Y(n4337) );
  INVX1 U909 ( .A(n4287), .Y(n4343) );
  INVX1 U910 ( .A(n4034), .Y(n4096) );
  INVX1 U911 ( .A(n4034), .Y(n4097) );
  INVX1 U912 ( .A(n4287), .Y(n4342) );
  INVX1 U913 ( .A(n4035), .Y(n4094) );
  INVX1 U914 ( .A(n4288), .Y(n4340) );
  INVX1 U915 ( .A(n4035), .Y(n4095) );
  INVX1 U916 ( .A(n4288), .Y(n4341) );
  INVX1 U917 ( .A(n4038), .Y(n4086) );
  INVX1 U918 ( .A(n4291), .Y(n4332) );
  INVX1 U919 ( .A(n4038), .Y(n4085) );
  INVX1 U920 ( .A(n4038), .Y(n4084) );
  INVX1 U921 ( .A(n4291), .Y(n4331) );
  INVX1 U922 ( .A(n4037), .Y(n4089) );
  INVX1 U923 ( .A(n4036), .Y(n4090) );
  INVX1 U924 ( .A(n4289), .Y(n4336) );
  INVX1 U925 ( .A(n4037), .Y(n4087) );
  INVX1 U926 ( .A(n4290), .Y(n4333) );
  INVX1 U927 ( .A(n4290), .Y(n4335) );
  INVX1 U928 ( .A(n4037), .Y(n4088) );
  INVX1 U929 ( .A(n4290), .Y(n4334) );
  INVX1 U930 ( .A(n4040), .Y(n4079) );
  INVX1 U931 ( .A(n4040), .Y(n4078) );
  INVX1 U932 ( .A(n4293), .Y(n4325) );
  INVX1 U933 ( .A(n4041), .Y(n4077) );
  INVX1 U934 ( .A(n4293), .Y(n4324) );
  INVX1 U935 ( .A(n4291), .Y(n4330) );
  INVX1 U936 ( .A(n4039), .Y(n4083) );
  INVX1 U937 ( .A(n4039), .Y(n4082) );
  INVX1 U938 ( .A(n4292), .Y(n4329) );
  INVX1 U939 ( .A(n4293), .Y(n4326) );
  INVX1 U940 ( .A(n4040), .Y(n4080) );
  INVX1 U941 ( .A(n4292), .Y(n4328) );
  INVX1 U942 ( .A(n4039), .Y(n4081) );
  INVX1 U943 ( .A(n4292), .Y(n4327) );
  INVX1 U944 ( .A(n4295), .Y(n4319) );
  INVX1 U945 ( .A(n4043), .Y(n4071) );
  INVX1 U946 ( .A(n4043), .Y(n4070) );
  INVX1 U947 ( .A(n4295), .Y(n4318) );
  INVX1 U948 ( .A(n4041), .Y(n4076) );
  INVX1 U949 ( .A(n4294), .Y(n4322) );
  INVX1 U950 ( .A(n4041), .Y(n4075) );
  INVX1 U951 ( .A(n4294), .Y(n4323) );
  INVX1 U952 ( .A(n4042), .Y(n4072) );
  INVX1 U953 ( .A(n4295), .Y(n4320) );
  INVX1 U954 ( .A(n4042), .Y(n4073) );
  INVX1 U955 ( .A(n4042), .Y(n4074) );
  INVX1 U956 ( .A(n4294), .Y(n4321) );
  INVX1 U957 ( .A(n4045), .Y(n4065) );
  INVX1 U958 ( .A(n4048), .Y(n4064) );
  INVX1 U959 ( .A(n4296), .Y(n4317) );
  INVX1 U960 ( .A(n4043), .Y(n4069) );
  INVX1 U961 ( .A(n4044), .Y(n4068) );
  INVX1 U962 ( .A(n4296), .Y(n4316) );
  INVX1 U963 ( .A(n4296), .Y(n4315) );
  INVX1 U964 ( .A(n4044), .Y(n4067) );
  INVX1 U965 ( .A(n4044), .Y(n4066) );
  INVX1 U966 ( .A(n4046), .Y(n4058) );
  INVX1 U967 ( .A(n4047), .Y(n4057) );
  INVX1 U968 ( .A(n4045), .Y(n4063) );
  INVX1 U969 ( .A(n4045), .Y(n4062) );
  INVX1 U970 ( .A(n4046), .Y(n4059) );
  INVX1 U971 ( .A(n4045), .Y(n4061) );
  INVX1 U972 ( .A(n4046), .Y(n4060) );
  INVX1 U973 ( .A(n4047), .Y(n4056) );
  INVX1 U974 ( .A(n4047), .Y(n4055) );
  INVX1 U975 ( .A(n4048), .Y(n4052) );
  INVX1 U976 ( .A(n4048), .Y(n4054) );
  INVX1 U977 ( .A(n4048), .Y(n4053) );
  INVX1 U978 ( .A(n7639), .Y(n7654) );
  INVX1 U979 ( .A(n7639), .Y(n7655) );
  INVX1 U980 ( .A(n7639), .Y(n7656) );
  INVX1 U981 ( .A(n7640), .Y(n7649) );
  INVX1 U982 ( .A(n7641), .Y(n7648) );
  INVX1 U983 ( .A(n7641), .Y(n7647) );
  INVX1 U984 ( .A(n7620), .Y(n7653) );
  INVX1 U985 ( .A(n7620), .Y(n7652) );
  INVX1 U986 ( .A(n7640), .Y(n7650) );
  INVX1 U987 ( .A(n7640), .Y(n7651) );
  INVX1 U988 ( .A(n7640), .Y(n7643) );
  INVX1 U989 ( .A(n7394), .Y(n7396) );
  INVX1 U990 ( .A(n7393), .Y(n7397) );
  INVX1 U991 ( .A(n7641), .Y(n7642) );
  INVX1 U992 ( .A(n7641), .Y(n7646) );
  INVX1 U993 ( .A(n7641), .Y(n7645) );
  INVX1 U994 ( .A(n7639), .Y(n7644) );
  INVX1 U995 ( .A(n4032), .Y(n4104) );
  INVX1 U996 ( .A(n4286), .Y(n4348) );
  INVX1 U997 ( .A(n7380), .Y(n7382) );
  INVX1 U998 ( .A(n7380), .Y(n7381) );
  INVX1 U999 ( .A(n7626), .Y(n7628) );
  INVX1 U1000 ( .A(n7379), .Y(n7383) );
  INVX1 U1001 ( .A(n7627), .Y(n7629) );
  INVX1 U1002 ( .A(n7379), .Y(n7384) );
  INVX1 U1003 ( .A(n7627), .Y(n7630) );
  INVX1 U1004 ( .A(n7377), .Y(n7387) );
  INVX1 U1005 ( .A(n7378), .Y(n7385) );
  INVX1 U1006 ( .A(n7626), .Y(n7631) );
  INVX1 U1007 ( .A(n7378), .Y(n7386) );
  INVX1 U1008 ( .A(n7626), .Y(n7632) );
  INVX1 U1009 ( .A(n7625), .Y(n7633) );
  INVX1 U1010 ( .A(n7624), .Y(n7635) );
  INVX1 U1011 ( .A(n7376), .Y(n7389) );
  INVX1 U1012 ( .A(n7377), .Y(n7388) );
  INVX1 U1013 ( .A(n7625), .Y(n7634) );
  INVX1 U1014 ( .A(n7376), .Y(n7390) );
  INVX1 U1015 ( .A(n7623), .Y(n7637) );
  INVX1 U1016 ( .A(n7375), .Y(n7391) );
  INVX1 U1017 ( .A(n7624), .Y(n7636) );
  INVX1 U1018 ( .A(n7375), .Y(n7392) );
  INVX1 U1019 ( .A(n7374), .Y(n7394) );
  INVX1 U1020 ( .A(n7623), .Y(n7638) );
  INVX1 U1021 ( .A(n7374), .Y(n7393) );
  INVX1 U1022 ( .A(n7374), .Y(n7395) );
  CLKINVX3 U1023 ( .A(n4510), .Y(n4558) );
  CLKINVX3 U1024 ( .A(n4510), .Y(n4559) );
  CLKINVX3 U1025 ( .A(n7854), .Y(n7898) );
  CLKINVX3 U1026 ( .A(n7847), .Y(n7902) );
  CLKINVX3 U1027 ( .A(n7854), .Y(n7899) );
  CLKINVX3 U1028 ( .A(n7853), .Y(n7901) );
  CLKINVX3 U1029 ( .A(n7853), .Y(n7900) );
  INVX1 U1030 ( .A(n4507), .Y(n4523) );
  INVX1 U1031 ( .A(n4506), .Y(n4522) );
  INVX1 U1032 ( .A(n4506), .Y(n4521) );
  INVX1 U1033 ( .A(n4506), .Y(n4520) );
  INVX1 U1034 ( .A(n4506), .Y(n4519) );
  INVX1 U1035 ( .A(n4507), .Y(n4518) );
  INVX1 U1036 ( .A(n4508), .Y(n4516) );
  INVX1 U1037 ( .A(n4507), .Y(n4517) );
  INVX1 U1038 ( .A(n4509), .Y(n4513) );
  INVX1 U1039 ( .A(n4508), .Y(n4515) );
  INVX1 U1040 ( .A(n4508), .Y(n4514) );
  INVX1 U1041 ( .A(n4509), .Y(n4511) );
  INVX1 U1042 ( .A(n4509), .Y(n4512) );
  INVX1 U1043 ( .A(n7849), .Y(n7862) );
  INVX1 U1044 ( .A(n7849), .Y(n7864) );
  INVX1 U1045 ( .A(n7849), .Y(n7863) );
  INVX1 U1046 ( .A(n7850), .Y(n7861) );
  INVX1 U1047 ( .A(n7850), .Y(n7860) );
  INVX1 U1048 ( .A(n7851), .Y(n7857) );
  INVX1 U1049 ( .A(n7850), .Y(n7859) );
  INVX1 U1050 ( .A(n7851), .Y(n7858) );
  INVX1 U1051 ( .A(n7852), .Y(n7855) );
  INVX1 U1052 ( .A(n7851), .Y(n7856) );
  INVX1 U1053 ( .A(n4506), .Y(n4524) );
  INVX1 U1054 ( .A(n7849), .Y(n7865) );
  INVX1 U1055 ( .A(n4563), .Y(n4586) );
  INVX1 U1056 ( .A(n4563), .Y(n4585) );
  INVX1 U1057 ( .A(n4564), .Y(n4582) );
  INVX1 U1058 ( .A(n4563), .Y(n4584) );
  INVX1 U1059 ( .A(n4564), .Y(n4583) );
  INVX1 U1060 ( .A(n4564), .Y(n4581) );
  INVX1 U1061 ( .A(n4564), .Y(n4580) );
  INVX1 U1062 ( .A(n4565), .Y(n4578) );
  INVX1 U1063 ( .A(n4564), .Y(n4579) );
  INVX1 U1064 ( .A(n4566), .Y(n4575) );
  INVX1 U1065 ( .A(n4565), .Y(n4577) );
  INVX1 U1066 ( .A(n4566), .Y(n4576) );
  INVX1 U1067 ( .A(n4567), .Y(n4574) );
  INVX1 U1068 ( .A(n4567), .Y(n4573) );
  INVX1 U1069 ( .A(n4568), .Y(n4572) );
  INVX1 U1070 ( .A(n4569), .Y(n4570) );
  INVX1 U1071 ( .A(n4568), .Y(n4571) );
  INVX1 U1072 ( .A(n7906), .Y(n7929) );
  INVX1 U1073 ( .A(n7906), .Y(n7927) );
  INVX1 U1074 ( .A(n7906), .Y(n7928) );
  INVX1 U1075 ( .A(n7907), .Y(n7924) );
  INVX1 U1076 ( .A(n7906), .Y(n7926) );
  INVX1 U1077 ( .A(n7907), .Y(n7925) );
  INVX1 U1078 ( .A(n7907), .Y(n7923) );
  INVX1 U1079 ( .A(n7907), .Y(n7922) );
  INVX1 U1080 ( .A(n7908), .Y(n7920) );
  INVX1 U1081 ( .A(n7907), .Y(n7921) );
  INVX1 U1082 ( .A(n7909), .Y(n7917) );
  INVX1 U1083 ( .A(n7908), .Y(n7919) );
  INVX1 U1084 ( .A(n7909), .Y(n7918) );
  INVX1 U1085 ( .A(n7908), .Y(n7916) );
  INVX1 U1086 ( .A(n7909), .Y(n7915) );
  INVX1 U1087 ( .A(n7910), .Y(n7914) );
  INVX1 U1088 ( .A(n7911), .Y(n7912) );
  INVX1 U1089 ( .A(n7910), .Y(n7913) );
  BUFX3 U1090 ( .A(n8694), .Y(n8050) );
  BUFX3 U1091 ( .A(n8722), .Y(n8106) );
  BUFX3 U1092 ( .A(n8694), .Y(n8049) );
  BUFX3 U1093 ( .A(n8722), .Y(n8105) );
  BUFX3 U1094 ( .A(n8665), .Y(n7994) );
  BUFX4 U1095 ( .A(n8750), .Y(n8161) );
  BUFX3 U1096 ( .A(n8773), .Y(n8203) );
  BUFX3 U1097 ( .A(n8802), .Y(n8261) );
  BUFX3 U1098 ( .A(n8831), .Y(n8319) );
  BUFX3 U1099 ( .A(n8694), .Y(n8051) );
  BUFX3 U1100 ( .A(n8722), .Y(n8107) );
  BUFX3 U1101 ( .A(n8860), .Y(n8377) );
  INVX1 U1102 ( .A(n4297), .Y(n4312) );
  INVX1 U1103 ( .A(n4298), .Y(n4311) );
  INVX1 U1104 ( .A(n4297), .Y(n4313) );
  INVX1 U1105 ( .A(n4297), .Y(n4314) );
  INVX1 U1106 ( .A(n4299), .Y(n4307) );
  INVX1 U1107 ( .A(n4299), .Y(n4306) );
  INVX1 U1108 ( .A(n4298), .Y(n4310) );
  INVX1 U1109 ( .A(n4298), .Y(n4309) );
  INVX1 U1110 ( .A(n4298), .Y(n4308) );
  INVX1 U1111 ( .A(n4047), .Y(n4051) );
  INVX1 U1112 ( .A(n4046), .Y(n4049) );
  INVX1 U1113 ( .A(n4044), .Y(n4050) );
  INVX1 U1114 ( .A(n4300), .Y(n4301) );
  INVX1 U1115 ( .A(n4299), .Y(n4305) );
  INVX1 U1116 ( .A(n4300), .Y(n4302) );
  INVX1 U1117 ( .A(n4300), .Y(n4304) );
  INVX1 U1118 ( .A(n4300), .Y(n4303) );
  INVX1 U1119 ( .A(n8648), .Y(n7374) );
  INVX1 U1120 ( .A(n4031), .Y(n4033) );
  INVX1 U1121 ( .A(n4031), .Y(n4032) );
  INVX1 U1122 ( .A(n4285), .Y(n4286) );
  INVX1 U1123 ( .A(n4030), .Y(n4034) );
  INVX1 U1124 ( .A(n4284), .Y(n4287) );
  INVX1 U1125 ( .A(n4030), .Y(n4035) );
  INVX1 U1126 ( .A(n4284), .Y(n4288) );
  INVX1 U1127 ( .A(n4029), .Y(n4038) );
  INVX1 U1128 ( .A(n4029), .Y(n4036) );
  INVX1 U1129 ( .A(n4283), .Y(n4289) );
  INVX1 U1130 ( .A(n4029), .Y(n4037) );
  INVX1 U1131 ( .A(n4283), .Y(n4290) );
  INVX1 U1132 ( .A(n4282), .Y(n4291) );
  INVX1 U1133 ( .A(n4281), .Y(n4293) );
  INVX1 U1134 ( .A(n4028), .Y(n4040) );
  INVX1 U1135 ( .A(n4029), .Y(n4039) );
  INVX1 U1136 ( .A(n4282), .Y(n4292) );
  INVX1 U1137 ( .A(n4028), .Y(n4041) );
  INVX1 U1138 ( .A(n4280), .Y(n4295) );
  INVX1 U1139 ( .A(n4031), .Y(n4042) );
  INVX1 U1140 ( .A(n4281), .Y(n4294) );
  INVX1 U1141 ( .A(n4028), .Y(n4043) );
  INVX1 U1142 ( .A(n4280), .Y(n4296) );
  INVX1 U1143 ( .A(n4027), .Y(n4044) );
  INVX1 U1144 ( .A(n4027), .Y(n4045) );
  INVX1 U1145 ( .A(n4027), .Y(n4046) );
  INVX1 U1146 ( .A(n4027), .Y(n4047) );
  INVX1 U1147 ( .A(n4027), .Y(n4048) );
  INVX1 U1148 ( .A(n7622), .Y(n7639) );
  INVX1 U1149 ( .A(n7622), .Y(n7640) );
  INVX1 U1150 ( .A(n7622), .Y(n7641) );
  INVX1 U1151 ( .A(n7620), .Y(n7627) );
  INVX1 U1152 ( .A(n7620), .Y(n7626) );
  INVX1 U1153 ( .A(n7621), .Y(n7625) );
  INVX1 U1154 ( .A(n7621), .Y(n7624) );
  INVX1 U1155 ( .A(n7621), .Y(n7623) );
  INVX1 U1156 ( .A(n7371), .Y(n7380) );
  INVX1 U1157 ( .A(n7371), .Y(n7379) );
  INVX1 U1158 ( .A(n7372), .Y(n7378) );
  INVX1 U1159 ( .A(n7372), .Y(n7377) );
  INVX1 U1160 ( .A(n7373), .Y(n7376) );
  INVX1 U1161 ( .A(n7373), .Y(n7375) );
  CLKINVX3 U1162 ( .A(n4636), .Y(n4637) );
  CLKINVX3 U1163 ( .A(n4636), .Y(n4638) );
  CLKINVX3 U1164 ( .A(n8653), .Y(n4639) );
  CLKINVX3 U1165 ( .A(n8653), .Y(n4640) );
  CLKINVX3 U1166 ( .A(n8653), .Y(n4641) );
  CLKINVX3 U1167 ( .A(n4636), .Y(n4642) );
  CLKINVX3 U1168 ( .A(n8653), .Y(n4643) );
  CLKINVX3 U1169 ( .A(n4636), .Y(n4644) );
  CLKINVX3 U1170 ( .A(n7979), .Y(n7981) );
  CLKINVX3 U1171 ( .A(n8643), .Y(n7982) );
  CLKINVX3 U1172 ( .A(n7979), .Y(n7983) );
  CLKINVX3 U1173 ( .A(n8643), .Y(n7984) );
  CLKINVX3 U1174 ( .A(n8643), .Y(n7985) );
  CLKINVX3 U1175 ( .A(n7979), .Y(n7986) );
  CLKINVX3 U1176 ( .A(n8643), .Y(n7987) );
  CLKINVX3 U1177 ( .A(n7979), .Y(n7988) );
  CLKINVX3 U1178 ( .A(n4627), .Y(n4628) );
  CLKINVX3 U1179 ( .A(n4627), .Y(n4629) );
  CLKINVX3 U1180 ( .A(n4627), .Y(n4630) );
  CLKINVX3 U1181 ( .A(n4627), .Y(n4631) );
  CLKINVX3 U1182 ( .A(n8654), .Y(n4632) );
  CLKINVX3 U1183 ( .A(n8654), .Y(n4633) );
  CLKINVX3 U1184 ( .A(n8654), .Y(n4634) );
  CLKINVX3 U1185 ( .A(n8654), .Y(n4635) );
  CLKINVX3 U1186 ( .A(n8645), .Y(n7972) );
  CLKINVX3 U1187 ( .A(n7970), .Y(n7973) );
  CLKINVX3 U1188 ( .A(n7970), .Y(n7974) );
  CLKINVX3 U1189 ( .A(n7970), .Y(n7975) );
  CLKINVX3 U1190 ( .A(n7970), .Y(n7976) );
  CLKINVX3 U1191 ( .A(n8645), .Y(n7977) );
  CLKINVX3 U1192 ( .A(n8645), .Y(n7971) );
  INVX1 U1193 ( .A(n8656), .Y(n4563) );
  INVX1 U1194 ( .A(n4625), .Y(n4564) );
  INVX1 U1195 ( .A(n4562), .Y(n4565) );
  INVX1 U1196 ( .A(n4562), .Y(n4566) );
  INVX1 U1197 ( .A(n4562), .Y(n4567) );
  INVX1 U1198 ( .A(n7905), .Y(n7906) );
  INVX1 U1199 ( .A(n7905), .Y(n7907) );
  INVX1 U1200 ( .A(n7904), .Y(n7908) );
  INVX1 U1201 ( .A(n7904), .Y(n7909) );
  INVX1 U1202 ( .A(n4561), .Y(n4569) );
  INVX1 U1203 ( .A(n4561), .Y(n4568) );
  INVX1 U1204 ( .A(n7904), .Y(n7911) );
  INVX1 U1205 ( .A(n7904), .Y(n7910) );
  INVX1 U1206 ( .A(n4505), .Y(n4506) );
  INVX1 U1207 ( .A(n4505), .Y(n4507) );
  INVX1 U1208 ( .A(n4504), .Y(n4508) );
  INVX1 U1209 ( .A(n4504), .Y(n4509) );
  INVX1 U1210 ( .A(n7848), .Y(n7849) );
  INVX1 U1211 ( .A(n7847), .Y(n7850) );
  INVX1 U1212 ( .A(n7847), .Y(n7851) );
  INVX1 U1213 ( .A(n8647), .Y(n7852) );
  INVX1 U1214 ( .A(n4507), .Y(n4510) );
  INVX1 U1215 ( .A(n7852), .Y(n7854) );
  INVX1 U1216 ( .A(n7852), .Y(n7853) );
  AND2X2 U1217 ( .A(n8504), .B(n8611), .Y(n10) );
  AND2X2 U1218 ( .A(n8504), .B(n8608), .Y(n11) );
  AND2X2 U1219 ( .A(n8504), .B(n8606), .Y(n12) );
  AND2X2 U1220 ( .A(n8504), .B(n8603), .Y(n13) );
  AND2X2 U1221 ( .A(n8504), .B(n8599), .Y(n14) );
  AND2X2 U1222 ( .A(n8504), .B(n8596), .Y(n15) );
  AND2X2 U1223 ( .A(n8504), .B(n8593), .Y(n16) );
  AND2X2 U1224 ( .A(n8504), .B(n8590), .Y(n17) );
  AND2X2 U1225 ( .A(n8504), .B(n8588), .Y(n18) );
  AND2X2 U1226 ( .A(n8504), .B(n8584), .Y(n19) );
  AND2X2 U1227 ( .A(n8504), .B(n8582), .Y(n20) );
  AND2X2 U1228 ( .A(n8504), .B(n8579), .Y(n21) );
  AND2X2 U1229 ( .A(n8501), .B(n8611), .Y(n22) );
  AND2X2 U1230 ( .A(n8501), .B(n8608), .Y(n23) );
  AND2X2 U1231 ( .A(n8501), .B(n8606), .Y(n24) );
  AND2X2 U1232 ( .A(n8501), .B(n8603), .Y(n25) );
  AND2X2 U1233 ( .A(n8501), .B(n8599), .Y(n26) );
  AND2X2 U1234 ( .A(n8501), .B(n8596), .Y(n27) );
  AND2X2 U1235 ( .A(n8501), .B(n8593), .Y(n28) );
  AND2X2 U1236 ( .A(n8501), .B(n8590), .Y(n29) );
  AND2X2 U1237 ( .A(n8501), .B(n8588), .Y(n30) );
  AND2X2 U1238 ( .A(n8501), .B(n8584), .Y(n31) );
  AND2X2 U1239 ( .A(n8501), .B(n8582), .Y(n32) );
  AND2X2 U1240 ( .A(n8501), .B(n8579), .Y(n33) );
  AND2X2 U1241 ( .A(n8498), .B(n8611), .Y(n34) );
  AND2X2 U1242 ( .A(n8498), .B(n8608), .Y(n35) );
  AND2X2 U1243 ( .A(n8498), .B(n8606), .Y(n36) );
  AND2X2 U1244 ( .A(n8498), .B(n8603), .Y(n37) );
  AND2X2 U1245 ( .A(n8498), .B(n8599), .Y(n38) );
  AND2X2 U1246 ( .A(n8498), .B(n8596), .Y(n39) );
  AND2X2 U1247 ( .A(n8498), .B(n8593), .Y(n40) );
  AND2X2 U1248 ( .A(n8498), .B(n8590), .Y(n41) );
  AND2X2 U1249 ( .A(n8498), .B(n8588), .Y(n42) );
  AND2X2 U1250 ( .A(n8498), .B(n8584), .Y(n43) );
  AND2X2 U1251 ( .A(n8498), .B(n8582), .Y(n44) );
  AND2X2 U1252 ( .A(n8498), .B(n8579), .Y(n45) );
  AND2X2 U1253 ( .A(n8495), .B(n8611), .Y(n46) );
  AND2X2 U1254 ( .A(n8495), .B(n8608), .Y(n47) );
  AND2X2 U1255 ( .A(n8495), .B(n8606), .Y(n48) );
  AND2X2 U1256 ( .A(n8495), .B(n8603), .Y(n49) );
  AND2X2 U1257 ( .A(n8495), .B(n8599), .Y(n50) );
  AND2X2 U1258 ( .A(n8495), .B(n8596), .Y(n51) );
  AND2X2 U1259 ( .A(n8495), .B(n8593), .Y(n52) );
  AND2X2 U1260 ( .A(n8495), .B(n8590), .Y(n53) );
  AND2X2 U1261 ( .A(n8495), .B(n8588), .Y(n55) );
  AND2X2 U1262 ( .A(n8495), .B(n8584), .Y(n56) );
  AND2X2 U1263 ( .A(n8495), .B(n8582), .Y(n57) );
  AND2X2 U1264 ( .A(n8495), .B(n8579), .Y(n58) );
  AND2X2 U1265 ( .A(n8492), .B(n8611), .Y(n59) );
  AND2X2 U1266 ( .A(n8492), .B(n8608), .Y(n60) );
  AND2X2 U1267 ( .A(n8492), .B(n8606), .Y(n61) );
  AND2X2 U1268 ( .A(n8492), .B(n8603), .Y(n62) );
  AND2X2 U1269 ( .A(n8492), .B(n8599), .Y(n63) );
  AND2X2 U1270 ( .A(n8492), .B(n8596), .Y(n64) );
  AND2X2 U1271 ( .A(n8492), .B(n8593), .Y(n65) );
  AND2X2 U1272 ( .A(n8492), .B(n8590), .Y(n66) );
  AND2X2 U1273 ( .A(n8492), .B(n8588), .Y(n67) );
  AND2X2 U1274 ( .A(n8492), .B(n8584), .Y(n68) );
  AND2X2 U1275 ( .A(n8492), .B(n8582), .Y(n69) );
  AND2X2 U1276 ( .A(n8492), .B(n8579), .Y(n70) );
  AND2X2 U1277 ( .A(n8489), .B(n8611), .Y(n71) );
  AND2X2 U1278 ( .A(n8489), .B(n8608), .Y(n72) );
  AND2X2 U1279 ( .A(n8489), .B(n8606), .Y(n73) );
  AND2X2 U1280 ( .A(n8489), .B(n8603), .Y(n74) );
  AND2X2 U1281 ( .A(n8489), .B(n8599), .Y(n75) );
  AND2X2 U1282 ( .A(n8489), .B(n8596), .Y(n76) );
  AND2X2 U1283 ( .A(n8489), .B(n8593), .Y(n77) );
  AND2X2 U1284 ( .A(n8489), .B(n8590), .Y(n78) );
  AND2X2 U1285 ( .A(n8489), .B(n8588), .Y(n79) );
  AND2X2 U1286 ( .A(n8489), .B(n8584), .Y(n80) );
  AND2X2 U1287 ( .A(n8489), .B(n8582), .Y(n81) );
  AND2X2 U1288 ( .A(n8489), .B(n8579), .Y(n82) );
  AND2X2 U1289 ( .A(n8486), .B(n8611), .Y(n83) );
  AND2X2 U1290 ( .A(n8486), .B(n8608), .Y(n84) );
  AND2X2 U1291 ( .A(n8486), .B(n8606), .Y(n85) );
  AND2X2 U1292 ( .A(n8486), .B(n8603), .Y(n86) );
  AND2X2 U1293 ( .A(n8486), .B(n8599), .Y(n87) );
  AND2X2 U1294 ( .A(n8486), .B(n8596), .Y(n88) );
  AND2X2 U1295 ( .A(n8486), .B(n8593), .Y(n89) );
  AND2X2 U1296 ( .A(n8486), .B(n8590), .Y(n90) );
  AND2X2 U1297 ( .A(n8486), .B(n8588), .Y(n91) );
  AND2X2 U1298 ( .A(n8486), .B(n8584), .Y(n92) );
  AND2X2 U1299 ( .A(n8486), .B(n8582), .Y(n93) );
  AND2X2 U1300 ( .A(n8486), .B(n8579), .Y(n94) );
  AND2X2 U1301 ( .A(n8483), .B(n8611), .Y(n95) );
  AND2X2 U1302 ( .A(n8483), .B(n8608), .Y(n96) );
  AND2X2 U1303 ( .A(n8483), .B(n8606), .Y(n97) );
  AND2X2 U1304 ( .A(n8483), .B(n8603), .Y(n98) );
  AND2X2 U1305 ( .A(n8483), .B(n8599), .Y(n99) );
  AND2X2 U1306 ( .A(n8483), .B(n8596), .Y(n100) );
  AND2X2 U1307 ( .A(n8483), .B(n8593), .Y(n101) );
  AND2X2 U1308 ( .A(n8483), .B(n8590), .Y(n102) );
  AND2X2 U1309 ( .A(n8483), .B(n8588), .Y(n103) );
  AND2X2 U1310 ( .A(n8483), .B(n8584), .Y(n104) );
  AND2X2 U1311 ( .A(n8483), .B(n8582), .Y(n105) );
  AND2X2 U1312 ( .A(n8483), .B(n8579), .Y(n106) );
  AND2X2 U1313 ( .A(n8480), .B(n8611), .Y(n107) );
  AND2X2 U1314 ( .A(n8480), .B(n8608), .Y(n108) );
  AND2X2 U1315 ( .A(n8480), .B(n8606), .Y(n109) );
  AND2X2 U1316 ( .A(n8480), .B(n8603), .Y(n110) );
  AND2X2 U1317 ( .A(n8480), .B(n8599), .Y(n111) );
  AND2X2 U1318 ( .A(n8480), .B(n8596), .Y(n112) );
  AND2X2 U1319 ( .A(n8480), .B(n8593), .Y(n113) );
  AND2X2 U1320 ( .A(n8480), .B(n8590), .Y(n114) );
  AND2X2 U1321 ( .A(n8480), .B(n8588), .Y(n115) );
  AND2X2 U1322 ( .A(n8480), .B(n8584), .Y(n116) );
  AND2X2 U1323 ( .A(n8480), .B(n8582), .Y(n117) );
  AND2X2 U1324 ( .A(n8480), .B(n8579), .Y(n118) );
  AND2X2 U1325 ( .A(n8477), .B(n8611), .Y(n119) );
  AND2X2 U1326 ( .A(n8477), .B(n8608), .Y(n120) );
  AND2X2 U1327 ( .A(n8477), .B(n8606), .Y(n121) );
  AND2X2 U1328 ( .A(n8477), .B(n8603), .Y(n122) );
  AND2X2 U1329 ( .A(n8477), .B(n8599), .Y(n123) );
  AND2X2 U1330 ( .A(n8477), .B(n8596), .Y(n124) );
  AND2X2 U1331 ( .A(n8477), .B(n8593), .Y(n125) );
  AND2X2 U1332 ( .A(n8477), .B(n8590), .Y(n126) );
  AND2X2 U1333 ( .A(n8477), .B(n8588), .Y(n127) );
  AND2X2 U1334 ( .A(n8477), .B(n8584), .Y(n128) );
  AND2X2 U1335 ( .A(n8477), .B(n8582), .Y(n129) );
  AND2X2 U1336 ( .A(n8477), .B(n8579), .Y(n130) );
  AND2X2 U1337 ( .A(n8474), .B(n8611), .Y(n131) );
  AND2X2 U1338 ( .A(n8474), .B(n8608), .Y(n132) );
  AND2X2 U1339 ( .A(n8474), .B(n8606), .Y(n133) );
  AND2X2 U1340 ( .A(n8474), .B(n8603), .Y(n134) );
  AND2X2 U1341 ( .A(n8474), .B(n8599), .Y(n135) );
  AND2X2 U1342 ( .A(n8474), .B(n8596), .Y(n136) );
  AND2X2 U1343 ( .A(n8474), .B(n8593), .Y(n137) );
  AND2X2 U1344 ( .A(n8474), .B(n8590), .Y(n138) );
  AND2X2 U1345 ( .A(n8474), .B(n8588), .Y(n139) );
  AND2X2 U1346 ( .A(n8474), .B(n8584), .Y(n140) );
  AND2X2 U1347 ( .A(n8474), .B(n8582), .Y(n141) );
  AND2X2 U1348 ( .A(n8474), .B(n8579), .Y(n142) );
  AND2X2 U1349 ( .A(n8471), .B(n8611), .Y(n143) );
  AND2X2 U1350 ( .A(n8471), .B(n8608), .Y(n144) );
  AND2X2 U1351 ( .A(n8471), .B(n8606), .Y(n145) );
  AND2X2 U1352 ( .A(n8471), .B(n8603), .Y(n146) );
  AND2X2 U1353 ( .A(n8471), .B(n8599), .Y(n147) );
  AND2X2 U1354 ( .A(n8471), .B(n8596), .Y(n148) );
  AND2X2 U1355 ( .A(n8471), .B(n8593), .Y(n149) );
  AND2X2 U1356 ( .A(n8471), .B(n8590), .Y(n150) );
  AND2X2 U1357 ( .A(n8471), .B(n8588), .Y(n151) );
  AND2X2 U1358 ( .A(n8471), .B(n8584), .Y(n152) );
  AND2X2 U1359 ( .A(n8471), .B(n8582), .Y(n153) );
  AND2X2 U1360 ( .A(n8471), .B(n8579), .Y(n154) );
  AND2X2 U1361 ( .A(n8468), .B(n8611), .Y(n155) );
  AND2X2 U1362 ( .A(n8468), .B(n8608), .Y(n156) );
  AND2X2 U1363 ( .A(n8468), .B(n8606), .Y(n157) );
  AND2X2 U1364 ( .A(n8468), .B(n8603), .Y(n158) );
  AND2X2 U1365 ( .A(n8468), .B(n8599), .Y(n159) );
  AND2X2 U1366 ( .A(n8468), .B(n8596), .Y(n160) );
  AND2X2 U1367 ( .A(n8468), .B(n8593), .Y(n161) );
  AND2X2 U1368 ( .A(n8468), .B(n8590), .Y(n162) );
  AND2X2 U1369 ( .A(n8468), .B(n8588), .Y(n163) );
  AND2X2 U1370 ( .A(n8468), .B(n8584), .Y(n164) );
  AND2X2 U1371 ( .A(n8468), .B(n8582), .Y(n165) );
  AND2X2 U1372 ( .A(n8468), .B(n8579), .Y(n166) );
  AND2X2 U1373 ( .A(n8465), .B(n8612), .Y(n167) );
  AND2X2 U1374 ( .A(n8465), .B(n8609), .Y(n168) );
  AND2X2 U1375 ( .A(n8465), .B(n8606), .Y(n169) );
  AND2X2 U1376 ( .A(n8465), .B(n8603), .Y(n170) );
  AND2X2 U1377 ( .A(n8465), .B(n8600), .Y(n171) );
  AND2X2 U1378 ( .A(n8465), .B(n8597), .Y(n172) );
  AND2X2 U1379 ( .A(n8465), .B(n8594), .Y(n173) );
  AND2X2 U1380 ( .A(n8465), .B(n8591), .Y(n174) );
  AND2X2 U1381 ( .A(n8465), .B(n8588), .Y(n175) );
  AND2X2 U1382 ( .A(n8465), .B(n8585), .Y(n176) );
  AND2X2 U1383 ( .A(n8465), .B(n8582), .Y(n177) );
  AND2X2 U1384 ( .A(n8465), .B(n8579), .Y(n178) );
  AND2X2 U1385 ( .A(n8462), .B(n8612), .Y(n179) );
  AND2X2 U1386 ( .A(n8462), .B(n8609), .Y(n180) );
  AND2X2 U1387 ( .A(n8462), .B(n1290), .Y(n181) );
  AND2X2 U1388 ( .A(n8462), .B(n1292), .Y(n182) );
  AND2X2 U1389 ( .A(n8462), .B(n8600), .Y(n183) );
  AND2X2 U1390 ( .A(n8462), .B(n8597), .Y(n184) );
  AND2X2 U1391 ( .A(n8462), .B(n8594), .Y(n185) );
  AND2X2 U1392 ( .A(n8462), .B(n8591), .Y(n186) );
  AND2X2 U1393 ( .A(n8462), .B(n1302), .Y(n187) );
  AND2X2 U1394 ( .A(n8462), .B(n8585), .Y(n188) );
  AND2X2 U1395 ( .A(n8462), .B(n1306), .Y(n189) );
  AND2X2 U1396 ( .A(n8462), .B(n1308), .Y(n190) );
  AND2X2 U1397 ( .A(n8459), .B(n8612), .Y(n191) );
  AND2X2 U1398 ( .A(n8459), .B(n8609), .Y(n192) );
  AND2X2 U1399 ( .A(n8459), .B(n1290), .Y(n193) );
  AND2X2 U1400 ( .A(n8459), .B(n1292), .Y(n194) );
  AND2X2 U1401 ( .A(n8459), .B(n8600), .Y(n195) );
  AND2X2 U1402 ( .A(n8459), .B(n8597), .Y(n196) );
  AND2X2 U1403 ( .A(n8459), .B(n8594), .Y(n197) );
  AND2X2 U1404 ( .A(n8459), .B(n8591), .Y(n198) );
  AND2X2 U1405 ( .A(n8459), .B(n1302), .Y(n199) );
  AND2X2 U1406 ( .A(n8459), .B(n8585), .Y(n200) );
  AND2X2 U1407 ( .A(n8459), .B(n1306), .Y(n201) );
  AND2X2 U1408 ( .A(n8459), .B(n1308), .Y(n202) );
  AND2X2 U1409 ( .A(n8456), .B(n8612), .Y(n203) );
  AND2X2 U1410 ( .A(n8456), .B(n8609), .Y(n204) );
  AND2X2 U1411 ( .A(n8456), .B(n1290), .Y(n205) );
  AND2X2 U1412 ( .A(n8456), .B(n1292), .Y(n206) );
  AND2X2 U1413 ( .A(n8456), .B(n8600), .Y(n207) );
  AND2X2 U1414 ( .A(n8456), .B(n8597), .Y(n208) );
  AND2X2 U1415 ( .A(n8456), .B(n8594), .Y(n209) );
  AND2X2 U1416 ( .A(n8456), .B(n8591), .Y(n210) );
  AND2X2 U1417 ( .A(n8456), .B(n1302), .Y(n211) );
  AND2X2 U1418 ( .A(n8456), .B(n8585), .Y(n212) );
  AND2X2 U1419 ( .A(n8456), .B(n1306), .Y(n213) );
  AND2X2 U1420 ( .A(n8456), .B(n1308), .Y(n214) );
  AND2X2 U1421 ( .A(n8453), .B(n8612), .Y(n215) );
  AND2X2 U1422 ( .A(n8453), .B(n8609), .Y(n216) );
  AND2X2 U1423 ( .A(n8453), .B(n1290), .Y(n217) );
  AND2X2 U1424 ( .A(n8453), .B(n1292), .Y(n218) );
  AND2X2 U1425 ( .A(n8453), .B(n8600), .Y(n219) );
  AND2X2 U1426 ( .A(n8453), .B(n8597), .Y(n220) );
  AND2X2 U1427 ( .A(n8453), .B(n8594), .Y(n221) );
  AND2X2 U1428 ( .A(n8453), .B(n8591), .Y(n222) );
  AND2X2 U1429 ( .A(n8453), .B(n1302), .Y(n223) );
  AND2X2 U1430 ( .A(n8453), .B(n8585), .Y(n224) );
  AND2X2 U1431 ( .A(n8453), .B(n1306), .Y(n225) );
  AND2X2 U1432 ( .A(n8453), .B(n1308), .Y(n226) );
  AND2X2 U1433 ( .A(n8450), .B(n8612), .Y(n227) );
  AND2X2 U1434 ( .A(n8450), .B(n8609), .Y(n228) );
  AND2X2 U1435 ( .A(n8450), .B(n1290), .Y(n229) );
  AND2X2 U1436 ( .A(n8450), .B(n1292), .Y(n230) );
  AND2X2 U1437 ( .A(n8450), .B(n8600), .Y(n231) );
  AND2X2 U1438 ( .A(n8450), .B(n8597), .Y(n232) );
  AND2X2 U1439 ( .A(n8450), .B(n8594), .Y(n233) );
  AND2X2 U1440 ( .A(n8450), .B(n8591), .Y(n234) );
  AND2X2 U1441 ( .A(n8450), .B(n1302), .Y(n235) );
  AND2X2 U1442 ( .A(n8450), .B(n8585), .Y(n236) );
  AND2X2 U1443 ( .A(n8450), .B(n1306), .Y(n237) );
  AND2X2 U1444 ( .A(n8450), .B(n1308), .Y(n238) );
  AND2X2 U1445 ( .A(n1740), .B(n8636), .Y(n239) );
  AND2X2 U1446 ( .A(n1740), .B(n8630), .Y(n240) );
  AND2X2 U1447 ( .A(n1740), .B(n8627), .Y(n241) );
  AND2X2 U1448 ( .A(n1740), .B(n8624), .Y(n242) );
  AND2X2 U1449 ( .A(n1740), .B(n8621), .Y(n243) );
  AND2X2 U1450 ( .A(n1740), .B(n8618), .Y(n244) );
  AND2X2 U1451 ( .A(n1740), .B(n8615), .Y(n245) );
  AND2X2 U1452 ( .A(n1773), .B(n8636), .Y(n246) );
  AND2X2 U1453 ( .A(n1773), .B(n8630), .Y(n247) );
  AND2X2 U1454 ( .A(n1773), .B(n8627), .Y(n248) );
  AND2X2 U1455 ( .A(n1773), .B(n8624), .Y(n249) );
  AND2X2 U1456 ( .A(n1773), .B(n8621), .Y(n250) );
  AND2X2 U1457 ( .A(n1773), .B(n8618), .Y(n251) );
  AND2X2 U1458 ( .A(n1773), .B(n8615), .Y(n252) );
  AND2X2 U1459 ( .A(n1806), .B(n8636), .Y(n253) );
  AND2X2 U1460 ( .A(n1806), .B(n8630), .Y(n254) );
  AND2X2 U1461 ( .A(n1806), .B(n8627), .Y(n255) );
  AND2X2 U1462 ( .A(n1806), .B(n8624), .Y(n256) );
  AND2X2 U1463 ( .A(n1806), .B(n8621), .Y(n257) );
  AND2X2 U1464 ( .A(n1806), .B(n8618), .Y(n258) );
  AND2X2 U1465 ( .A(n1806), .B(n8615), .Y(n259) );
  AND2X2 U1466 ( .A(n1839), .B(n8636), .Y(n260) );
  AND2X2 U1467 ( .A(n1839), .B(n8630), .Y(n261) );
  AND2X2 U1468 ( .A(n1839), .B(n8627), .Y(n262) );
  AND2X2 U1469 ( .A(n1839), .B(n8624), .Y(n263) );
  AND2X2 U1470 ( .A(n1839), .B(n8621), .Y(n264) );
  AND2X2 U1471 ( .A(n1839), .B(n8618), .Y(n265) );
  AND2X2 U1472 ( .A(n1839), .B(n8615), .Y(n266) );
  AND2X2 U1473 ( .A(n1873), .B(n8636), .Y(n267) );
  AND2X2 U1474 ( .A(n1873), .B(n8630), .Y(n268) );
  AND2X2 U1475 ( .A(n1873), .B(n8627), .Y(n269) );
  AND2X2 U1476 ( .A(n1873), .B(n8624), .Y(n270) );
  AND2X2 U1477 ( .A(n1873), .B(n8621), .Y(n271) );
  AND2X2 U1478 ( .A(n1873), .B(n8618), .Y(n272) );
  AND2X2 U1479 ( .A(n1873), .B(n8615), .Y(n273) );
  AND2X2 U1480 ( .A(n1906), .B(n8636), .Y(n274) );
  AND2X2 U1481 ( .A(n1906), .B(n8630), .Y(n275) );
  AND2X2 U1482 ( .A(n1906), .B(n8627), .Y(n276) );
  AND2X2 U1483 ( .A(n1906), .B(n8624), .Y(n277) );
  AND2X2 U1484 ( .A(n1906), .B(n8621), .Y(n278) );
  AND2X2 U1485 ( .A(n1906), .B(n8618), .Y(n279) );
  AND2X2 U1486 ( .A(n1906), .B(n8615), .Y(n280) );
  AND2X2 U1487 ( .A(n1939), .B(n8636), .Y(n281) );
  AND2X2 U1488 ( .A(n1939), .B(n8630), .Y(n282) );
  AND2X2 U1489 ( .A(n1939), .B(n8627), .Y(n283) );
  AND2X2 U1490 ( .A(n1939), .B(n8624), .Y(n284) );
  AND2X2 U1491 ( .A(n1939), .B(n8621), .Y(n285) );
  AND2X2 U1492 ( .A(n1939), .B(n8618), .Y(n286) );
  AND2X2 U1493 ( .A(n1939), .B(n8615), .Y(n287) );
  AND2X2 U1494 ( .A(n1972), .B(n8636), .Y(n288) );
  AND2X2 U1495 ( .A(n1972), .B(n8630), .Y(n289) );
  AND2X2 U1496 ( .A(n1972), .B(n8627), .Y(n290) );
  AND2X2 U1497 ( .A(n1972), .B(n8624), .Y(n291) );
  AND2X2 U1498 ( .A(n1972), .B(n8621), .Y(n292) );
  AND2X2 U1499 ( .A(n1972), .B(n8618), .Y(n293) );
  AND2X2 U1500 ( .A(n1972), .B(n8615), .Y(n294) );
  AND2X2 U1501 ( .A(n2005), .B(n8636), .Y(n295) );
  AND2X2 U1502 ( .A(n2005), .B(n8630), .Y(n296) );
  AND2X2 U1503 ( .A(n2005), .B(n8627), .Y(n297) );
  AND2X2 U1504 ( .A(n2005), .B(n8624), .Y(n298) );
  AND2X2 U1505 ( .A(n2005), .B(n8621), .Y(n299) );
  AND2X2 U1506 ( .A(n2005), .B(n8618), .Y(n300) );
  AND2X2 U1507 ( .A(n2005), .B(n8615), .Y(n301) );
  AND2X2 U1508 ( .A(n2038), .B(n8636), .Y(n302) );
  AND2X2 U1509 ( .A(n2038), .B(n8630), .Y(n303) );
  AND2X2 U1510 ( .A(n2038), .B(n8627), .Y(n304) );
  AND2X2 U1511 ( .A(n2038), .B(n8624), .Y(n305) );
  AND2X2 U1512 ( .A(n2038), .B(n8621), .Y(n306) );
  AND2X2 U1513 ( .A(n2038), .B(n8618), .Y(n307) );
  AND2X2 U1514 ( .A(n2038), .B(n8615), .Y(n308) );
  AND2X2 U1515 ( .A(n2071), .B(n8636), .Y(n309) );
  AND2X2 U1516 ( .A(n2071), .B(n8630), .Y(n310) );
  AND2X2 U1517 ( .A(n2071), .B(n8627), .Y(n311) );
  AND2X2 U1518 ( .A(n2071), .B(n8624), .Y(n312) );
  AND2X2 U1519 ( .A(n2071), .B(n8621), .Y(n313) );
  AND2X2 U1520 ( .A(n2071), .B(n8618), .Y(n314) );
  AND2X2 U1521 ( .A(n2071), .B(n8615), .Y(n315) );
  AND2X2 U1522 ( .A(n2104), .B(n8636), .Y(n316) );
  AND2X2 U1523 ( .A(n2104), .B(n8630), .Y(n317) );
  AND2X2 U1524 ( .A(n2104), .B(n8627), .Y(n318) );
  AND2X2 U1525 ( .A(n2104), .B(n8624), .Y(n319) );
  AND2X2 U1526 ( .A(n2104), .B(n8621), .Y(n320) );
  AND2X2 U1527 ( .A(n2104), .B(n8618), .Y(n321) );
  AND2X2 U1528 ( .A(n2104), .B(n8615), .Y(n322) );
  AND2X2 U1529 ( .A(n2138), .B(n8636), .Y(n323) );
  AND2X2 U1530 ( .A(n2138), .B(n8630), .Y(n324) );
  AND2X2 U1531 ( .A(n2138), .B(n8627), .Y(n325) );
  AND2X2 U1532 ( .A(n2138), .B(n8624), .Y(n326) );
  AND2X2 U1533 ( .A(n2138), .B(n8621), .Y(n327) );
  AND2X2 U1534 ( .A(n2138), .B(n8618), .Y(n328) );
  AND2X2 U1535 ( .A(n2138), .B(n8615), .Y(n329) );
  AND2X2 U1536 ( .A(n1573), .B(n8638), .Y(n330) );
  AND2X2 U1537 ( .A(n1608), .B(n8638), .Y(n331) );
  AND2X2 U1538 ( .A(n1641), .B(n8638), .Y(n332) );
  AND2X2 U1539 ( .A(n1674), .B(n8638), .Y(n333) );
  AND2X2 U1540 ( .A(n1707), .B(n8638), .Y(n334) );
  AND2X2 U1541 ( .A(n1740), .B(n8638), .Y(n335) );
  AND2X2 U1542 ( .A(n1773), .B(n8638), .Y(n336) );
  AND2X2 U1543 ( .A(n1806), .B(n8638), .Y(n337) );
  AND2X2 U1544 ( .A(n1839), .B(n8638), .Y(n338) );
  AND2X2 U1545 ( .A(n1873), .B(n8638), .Y(n339) );
  AND2X2 U1546 ( .A(n1906), .B(n8638), .Y(n340) );
  AND2X2 U1547 ( .A(n1939), .B(n8638), .Y(n341) );
  AND2X2 U1548 ( .A(n1334), .B(n8639), .Y(n342) );
  AND2X2 U1549 ( .A(n1369), .B(n8639), .Y(n343) );
  AND2X2 U1550 ( .A(n1403), .B(n8639), .Y(n344) );
  AND2X2 U1551 ( .A(n2171), .B(n8636), .Y(n345) );
  AND2X2 U1552 ( .A(n2171), .B(n8630), .Y(n346) );
  AND2X2 U1553 ( .A(n2171), .B(n8627), .Y(n347) );
  AND2X2 U1554 ( .A(n2171), .B(n8624), .Y(n348) );
  AND2X2 U1555 ( .A(n2171), .B(n8621), .Y(n349) );
  AND2X2 U1556 ( .A(n2171), .B(n8618), .Y(n350) );
  AND2X2 U1557 ( .A(n2171), .B(n8615), .Y(n351) );
  AND2X2 U1558 ( .A(n2204), .B(n1271), .Y(n352) );
  AND2X2 U1559 ( .A(n2204), .B(n1274), .Y(n353) );
  AND2X2 U1560 ( .A(n2204), .B(n1276), .Y(n354) );
  AND2X2 U1561 ( .A(n2204), .B(n1278), .Y(n355) );
  AND2X2 U1562 ( .A(n2204), .B(n1280), .Y(n356) );
  AND2X2 U1563 ( .A(n2204), .B(n1282), .Y(n357) );
  AND2X2 U1564 ( .A(n2204), .B(n1284), .Y(n358) );
  AND2X2 U1565 ( .A(n2237), .B(n1271), .Y(n359) );
  AND2X2 U1566 ( .A(n2237), .B(n1274), .Y(n360) );
  AND2X2 U1567 ( .A(n2237), .B(n1276), .Y(n361) );
  AND2X2 U1568 ( .A(n2237), .B(n1278), .Y(n362) );
  AND2X2 U1569 ( .A(n2237), .B(n1280), .Y(n363) );
  AND2X2 U1570 ( .A(n2237), .B(n1282), .Y(n364) );
  AND2X2 U1571 ( .A(n2237), .B(n1284), .Y(n365) );
  AND2X2 U1572 ( .A(n2270), .B(n1271), .Y(n366) );
  AND2X2 U1573 ( .A(n2270), .B(n1274), .Y(n367) );
  AND2X2 U1574 ( .A(n2270), .B(n1276), .Y(n368) );
  AND2X2 U1575 ( .A(n2270), .B(n1278), .Y(n369) );
  AND2X2 U1576 ( .A(n2270), .B(n1280), .Y(n370) );
  AND2X2 U1577 ( .A(n2270), .B(n1282), .Y(n371) );
  AND2X2 U1578 ( .A(n2270), .B(n1284), .Y(n372) );
  AND2X2 U1579 ( .A(n2303), .B(n1271), .Y(n373) );
  AND2X2 U1580 ( .A(n2303), .B(n1274), .Y(n374) );
  AND2X2 U1581 ( .A(n2303), .B(n1276), .Y(n375) );
  AND2X2 U1582 ( .A(n2303), .B(n1278), .Y(n376) );
  AND2X2 U1583 ( .A(n2303), .B(n1280), .Y(n377) );
  AND2X2 U1584 ( .A(n2303), .B(n1282), .Y(n378) );
  AND2X2 U1585 ( .A(n2303), .B(n1284), .Y(n379) );
  AND2X2 U1586 ( .A(n2336), .B(n1271), .Y(n380) );
  AND2X2 U1587 ( .A(n2336), .B(n1274), .Y(n381) );
  AND2X2 U1588 ( .A(n2336), .B(n1276), .Y(n382) );
  AND2X2 U1589 ( .A(n2336), .B(n1278), .Y(n383) );
  AND2X2 U1590 ( .A(n2336), .B(n1280), .Y(n384) );
  AND2X2 U1591 ( .A(n2336), .B(n1282), .Y(n385) );
  AND2X2 U1592 ( .A(n2336), .B(n1284), .Y(n386) );
  CLKINVX3 U1593 ( .A(n8634), .Y(n8633) );
  AND2X2 U1594 ( .A(n1437), .B(n8639), .Y(n387) );
  AND2X2 U1595 ( .A(n1471), .B(n8639), .Y(n388) );
  AND2X2 U1596 ( .A(n1505), .B(n8639), .Y(n389) );
  AND2X2 U1597 ( .A(n1539), .B(n8639), .Y(n390) );
  BUFX4 U1598 ( .A(n8758), .Y(n8187) );
  BUFX4 U1599 ( .A(n8758), .Y(n8186) );
  BUFX4 U1600 ( .A(n8758), .Y(n8185) );
  BUFX4 U1601 ( .A(n8759), .Y(n8190) );
  BUFX4 U1602 ( .A(n8759), .Y(n8189) );
  BUFX4 U1603 ( .A(n8759), .Y(n8188) );
  BUFX4 U1604 ( .A(n8752), .Y(n8169) );
  BUFX4 U1605 ( .A(n8752), .Y(n8168) );
  BUFX4 U1606 ( .A(n8752), .Y(n8167) );
  BUFX4 U1607 ( .A(n8751), .Y(n8163) );
  BUFX4 U1608 ( .A(n8751), .Y(n8162) );
  BUFX4 U1609 ( .A(n8162), .Y(n8165) );
  BUFX4 U1610 ( .A(n8762), .Y(n8164) );
  BUFX4 U1611 ( .A(n8763), .Y(n8166) );
  BUFX4 U1612 ( .A(n8756), .Y(n8181) );
  BUFX4 U1613 ( .A(n8756), .Y(n8180) );
  BUFX4 U1614 ( .A(n8756), .Y(n8179) );
  BUFX4 U1615 ( .A(n8757), .Y(n8183) );
  BUFX4 U1616 ( .A(n8757), .Y(n8182) );
  BUFX4 U1617 ( .A(n8753), .Y(n8172) );
  BUFX4 U1618 ( .A(n8753), .Y(n8171) );
  BUFX4 U1619 ( .A(n8753), .Y(n8170) );
  BUFX4 U1620 ( .A(n8754), .Y(n8175) );
  BUFX4 U1621 ( .A(n8754), .Y(n8174) );
  BUFX4 U1622 ( .A(n8754), .Y(n8173) );
  BUFX4 U1623 ( .A(n8755), .Y(n8176) );
  BUFX4 U1624 ( .A(n8755), .Y(n8178) );
  BUFX4 U1625 ( .A(n8755), .Y(n8177) );
  BUFX4 U1626 ( .A(n8757), .Y(n8184) );
  BUFX3 U1627 ( .A(n8782), .Y(n8240) );
  BUFX3 U1628 ( .A(n8811), .Y(n8298) );
  BUFX3 U1629 ( .A(n8840), .Y(n8356) );
  BUFX3 U1630 ( .A(n8869), .Y(n8414) );
  BUFX3 U1631 ( .A(n8782), .Y(n8239) );
  BUFX3 U1632 ( .A(n8811), .Y(n8297) );
  BUFX3 U1633 ( .A(n8840), .Y(n8355) );
  BUFX3 U1634 ( .A(n8869), .Y(n8413) );
  BUFX3 U1635 ( .A(n8674), .Y(n8029) );
  BUFX3 U1636 ( .A(n8706), .Y(n8089) );
  BUFX3 U1637 ( .A(n8734), .Y(n8145) );
  BUFX3 U1638 ( .A(n8674), .Y(n8030) );
  BUFX3 U1639 ( .A(n8706), .Y(n8090) );
  BUFX3 U1640 ( .A(n8734), .Y(n8146) );
  BUFX3 U1641 ( .A(n8674), .Y(n8028) );
  BUFX3 U1642 ( .A(n8706), .Y(n8088) );
  BUFX3 U1643 ( .A(n8734), .Y(n8144) );
  BUFX3 U1644 ( .A(n8783), .Y(n8243) );
  BUFX3 U1645 ( .A(n8812), .Y(n8301) );
  BUFX3 U1646 ( .A(n8841), .Y(n8359) );
  BUFX3 U1647 ( .A(n8870), .Y(n8417) );
  BUFX3 U1648 ( .A(n8783), .Y(n8242) );
  BUFX3 U1649 ( .A(n8812), .Y(n8300) );
  BUFX3 U1650 ( .A(n8841), .Y(n8358) );
  BUFX3 U1651 ( .A(n8870), .Y(n8416) );
  BUFX3 U1652 ( .A(n8675), .Y(n8033) );
  BUFX3 U1653 ( .A(n8707), .Y(n8093) );
  BUFX3 U1654 ( .A(n8735), .Y(n8149) );
  BUFX3 U1655 ( .A(n8675), .Y(n8032) );
  BUFX3 U1656 ( .A(n8707), .Y(n8092) );
  BUFX3 U1657 ( .A(n8735), .Y(n8148) );
  BUFX3 U1658 ( .A(n8675), .Y(n8031) );
  BUFX3 U1659 ( .A(n8707), .Y(n8091) );
  BUFX3 U1660 ( .A(n8735), .Y(n8147) );
  BUFX3 U1661 ( .A(n8780), .Y(n8234) );
  BUFX3 U1662 ( .A(n8809), .Y(n8292) );
  BUFX3 U1663 ( .A(n8838), .Y(n8350) );
  BUFX3 U1664 ( .A(n8867), .Y(n8408) );
  BUFX3 U1665 ( .A(n8780), .Y(n8233) );
  BUFX3 U1666 ( .A(n8809), .Y(n8291) );
  BUFX3 U1667 ( .A(n8838), .Y(n8349) );
  BUFX3 U1668 ( .A(n8867), .Y(n8407) );
  BUFX3 U1669 ( .A(n8672), .Y(n8024) );
  BUFX3 U1670 ( .A(n8672), .Y(n8023) );
  BUFX3 U1671 ( .A(n8704), .Y(n8084) );
  BUFX3 U1672 ( .A(n8732), .Y(n8140) );
  BUFX3 U1673 ( .A(n8672), .Y(n8022) );
  BUFX3 U1674 ( .A(n8704), .Y(n8083) );
  BUFX3 U1675 ( .A(n8732), .Y(n8139) );
  BUFX3 U1676 ( .A(n8704), .Y(n8082) );
  BUFX3 U1677 ( .A(n8732), .Y(n8138) );
  BUFX3 U1678 ( .A(n8673), .Y(n8026) );
  BUFX3 U1679 ( .A(n8673), .Y(n8025) );
  BUFX3 U1680 ( .A(n8705), .Y(n8086) );
  BUFX3 U1681 ( .A(n8733), .Y(n8142) );
  BUFX3 U1682 ( .A(n8781), .Y(n8236) );
  BUFX3 U1683 ( .A(n8810), .Y(n8294) );
  BUFX3 U1684 ( .A(n8839), .Y(n8352) );
  BUFX3 U1685 ( .A(n8868), .Y(n8410) );
  BUFX3 U1686 ( .A(n8673), .Y(n8027) );
  BUFX3 U1687 ( .A(n8705), .Y(n8085) );
  BUFX3 U1688 ( .A(n8733), .Y(n8141) );
  BUFX3 U1689 ( .A(n8705), .Y(n8087) );
  BUFX3 U1690 ( .A(n8733), .Y(n8143) );
  BUFX3 U1691 ( .A(n8781), .Y(n8237) );
  BUFX3 U1692 ( .A(n8810), .Y(n8295) );
  BUFX3 U1693 ( .A(n8839), .Y(n8353) );
  BUFX3 U1694 ( .A(n8868), .Y(n8411) );
  BUFX3 U1695 ( .A(n8679), .Y(n8043) );
  BUFX3 U1696 ( .A(n8679), .Y(n8045) );
  BUFX3 U1697 ( .A(n8710), .Y(n8102) );
  BUFX3 U1698 ( .A(n8738), .Y(n8158) );
  BUFX3 U1699 ( .A(n8679), .Y(n8044) );
  BUFX3 U1700 ( .A(n8710), .Y(n8104) );
  BUFX3 U1701 ( .A(n8738), .Y(n8160) );
  BUFX3 U1702 ( .A(n8710), .Y(n8103) );
  BUFX3 U1703 ( .A(n8738), .Y(n8159) );
  BUFX3 U1704 ( .A(n8788), .Y(n8257) );
  BUFX3 U1705 ( .A(n8817), .Y(n8315) );
  BUFX3 U1706 ( .A(n8846), .Y(n8373) );
  BUFX3 U1707 ( .A(n8875), .Y(n8431) );
  BUFX3 U1708 ( .A(n8788), .Y(n8256) );
  BUFX3 U1709 ( .A(n8817), .Y(n8314) );
  BUFX3 U1710 ( .A(n8846), .Y(n8372) );
  BUFX3 U1711 ( .A(n8875), .Y(n8430) );
  BUFX3 U1712 ( .A(n8680), .Y(n8048) );
  BUFX3 U1713 ( .A(n8680), .Y(n8047) );
  BUFX3 U1714 ( .A(n8680), .Y(n8046) );
  BUFX3 U1715 ( .A(n8784), .Y(n8246) );
  BUFX3 U1716 ( .A(n8813), .Y(n8304) );
  BUFX3 U1717 ( .A(n8842), .Y(n8362) );
  BUFX3 U1718 ( .A(n8871), .Y(n8420) );
  BUFX3 U1719 ( .A(n8784), .Y(n8245) );
  BUFX3 U1720 ( .A(n8813), .Y(n8303) );
  BUFX3 U1721 ( .A(n8842), .Y(n8361) );
  BUFX3 U1722 ( .A(n8871), .Y(n8419) );
  BUFX3 U1723 ( .A(n8676), .Y(n8036) );
  BUFX3 U1724 ( .A(n8676), .Y(n8035) );
  BUFX3 U1725 ( .A(n8676), .Y(n8034) );
  BUFX3 U1726 ( .A(n8708), .Y(n8095) );
  BUFX3 U1727 ( .A(n8736), .Y(n8151) );
  BUFX3 U1728 ( .A(n8708), .Y(n8094) );
  BUFX3 U1729 ( .A(n8736), .Y(n8150) );
  BUFX3 U1730 ( .A(n8785), .Y(n8249) );
  BUFX3 U1731 ( .A(n8814), .Y(n8307) );
  BUFX3 U1732 ( .A(n8843), .Y(n8365) );
  BUFX3 U1733 ( .A(n8872), .Y(n8423) );
  BUFX3 U1734 ( .A(n8785), .Y(n8248) );
  BUFX3 U1735 ( .A(n8814), .Y(n8306) );
  BUFX3 U1736 ( .A(n8843), .Y(n8364) );
  BUFX3 U1737 ( .A(n8872), .Y(n8422) );
  BUFX3 U1738 ( .A(n8677), .Y(n8039) );
  BUFX3 U1739 ( .A(n8677), .Y(n8038) );
  BUFX3 U1740 ( .A(n8709), .Y(n8098) );
  BUFX3 U1741 ( .A(n8737), .Y(n8154) );
  BUFX3 U1742 ( .A(n8677), .Y(n8037) );
  BUFX3 U1743 ( .A(n8709), .Y(n8097) );
  BUFX3 U1744 ( .A(n8737), .Y(n8153) );
  BUFX3 U1745 ( .A(n8709), .Y(n8096) );
  BUFX3 U1746 ( .A(n8737), .Y(n8152) );
  BUFX3 U1747 ( .A(n8786), .Y(n8252) );
  BUFX3 U1748 ( .A(n8815), .Y(n8310) );
  BUFX3 U1749 ( .A(n8844), .Y(n8368) );
  BUFX3 U1750 ( .A(n8873), .Y(n8426) );
  BUFX3 U1751 ( .A(n8786), .Y(n8251) );
  BUFX3 U1752 ( .A(n8815), .Y(n8309) );
  BUFX3 U1753 ( .A(n8844), .Y(n8367) );
  BUFX3 U1754 ( .A(n8873), .Y(n8425) );
  BUFX3 U1755 ( .A(n8678), .Y(n8040) );
  BUFX3 U1756 ( .A(n8678), .Y(n8042) );
  BUFX3 U1757 ( .A(n8700), .Y(n8099) );
  BUFX3 U1758 ( .A(n8728), .Y(n8155) );
  BUFX3 U1759 ( .A(n8678), .Y(n8041) );
  BUFX3 U1760 ( .A(n8701), .Y(n8101) );
  BUFX3 U1761 ( .A(n8729), .Y(n8157) );
  BUFX3 U1762 ( .A(n8787), .Y(n8255) );
  BUFX3 U1763 ( .A(n8816), .Y(n8313) );
  BUFX3 U1764 ( .A(n8845), .Y(n8371) );
  BUFX3 U1765 ( .A(n8874), .Y(n8429) );
  BUFX3 U1766 ( .A(n8696), .Y(n8100) );
  BUFX3 U1767 ( .A(n8724), .Y(n8156) );
  BUFX3 U1768 ( .A(n8787), .Y(n8254) );
  BUFX3 U1769 ( .A(n8816), .Y(n8312) );
  BUFX3 U1770 ( .A(n8845), .Y(n8370) );
  BUFX3 U1771 ( .A(n8874), .Y(n8428) );
  BUFX3 U1772 ( .A(n8663), .Y(n8000) );
  BUFX3 U1773 ( .A(data_in[0]), .Y(n7999) );
  BUFX3 U1774 ( .A(n8781), .Y(n8210) );
  BUFX3 U1775 ( .A(n8810), .Y(n8268) );
  BUFX3 U1776 ( .A(n8839), .Y(n8326) );
  BUFX3 U1777 ( .A(n8868), .Y(n8384) );
  BUFX3 U1778 ( .A(data_in[0]), .Y(n7998) );
  BUFX3 U1779 ( .A(n8696), .Y(n8060) );
  BUFX3 U1780 ( .A(n8724), .Y(n8116) );
  BUFX3 U1781 ( .A(n8696), .Y(n8059) );
  BUFX3 U1782 ( .A(n8724), .Y(n8115) );
  BUFX3 U1783 ( .A(n8696), .Y(n8058) );
  BUFX3 U1784 ( .A(n8724), .Y(n8114) );
  BUFX3 U1785 ( .A(n8774), .Y(n8213) );
  BUFX3 U1786 ( .A(n8803), .Y(n8271) );
  BUFX3 U1787 ( .A(n8832), .Y(n8329) );
  BUFX3 U1788 ( .A(n8861), .Y(n8387) );
  BUFX3 U1789 ( .A(n8774), .Y(n8212) );
  BUFX3 U1790 ( .A(n8803), .Y(n8270) );
  BUFX3 U1791 ( .A(n8832), .Y(n8328) );
  BUFX3 U1792 ( .A(n8861), .Y(n8386) );
  BUFX3 U1793 ( .A(n8689), .Y(n8003) );
  BUFX3 U1794 ( .A(n7994), .Y(n8002) );
  BUFX3 U1795 ( .A(n7994), .Y(n8001) );
  BUFX3 U1796 ( .A(n8697), .Y(n8063) );
  BUFX3 U1797 ( .A(n8725), .Y(n8119) );
  BUFX3 U1798 ( .A(n8697), .Y(n8062) );
  BUFX3 U1799 ( .A(n8725), .Y(n8118) );
  BUFX3 U1800 ( .A(n8697), .Y(n8061) );
  BUFX3 U1801 ( .A(n8725), .Y(n8117) );
  BUFX3 U1802 ( .A(n8785), .Y(n8205) );
  BUFX3 U1803 ( .A(n8814), .Y(n8263) );
  BUFX3 U1804 ( .A(n8843), .Y(n8321) );
  BUFX3 U1805 ( .A(n8872), .Y(n8379) );
  BUFX3 U1806 ( .A(n8705), .Y(n8054) );
  BUFX3 U1807 ( .A(n8733), .Y(n8110) );
  BUFX3 U1808 ( .A(n8786), .Y(n8204) );
  BUFX3 U1809 ( .A(n8815), .Y(n8262) );
  BUFX3 U1810 ( .A(n8844), .Y(n8320) );
  BUFX3 U1811 ( .A(n8873), .Y(n8378) );
  BUFX3 U1812 ( .A(n8674), .Y(n7995) );
  BUFX3 U1813 ( .A(n8710), .Y(n8053) );
  BUFX3 U1814 ( .A(n8738), .Y(n8109) );
  BUFX3 U1815 ( .A(n8698), .Y(n8052) );
  BUFX3 U1816 ( .A(n8726), .Y(n8108) );
  BUFX3 U1817 ( .A(n8695), .Y(n8055) );
  BUFX3 U1818 ( .A(n8723), .Y(n8111) );
  BUFX3 U1819 ( .A(n8784), .Y(n8207) );
  BUFX3 U1820 ( .A(n8813), .Y(n8265) );
  BUFX3 U1821 ( .A(n8842), .Y(n8323) );
  BUFX3 U1822 ( .A(n8871), .Y(n8381) );
  BUFX3 U1823 ( .A(n8679), .Y(n7997) );
  BUFX3 U1824 ( .A(n8695), .Y(n8057) );
  BUFX3 U1825 ( .A(n8723), .Y(n8113) );
  BUFX3 U1826 ( .A(n8678), .Y(n7996) );
  BUFX3 U1827 ( .A(n8695), .Y(n8056) );
  BUFX3 U1828 ( .A(n8723), .Y(n8112) );
  BUFX3 U1829 ( .A(n8782), .Y(n8208) );
  BUFX3 U1830 ( .A(n8811), .Y(n8266) );
  BUFX3 U1831 ( .A(n8840), .Y(n8324) );
  BUFX3 U1832 ( .A(n8869), .Y(n8382) );
  BUFX3 U1833 ( .A(n8786), .Y(n8225) );
  BUFX3 U1834 ( .A(n8815), .Y(n8283) );
  BUFX3 U1835 ( .A(n8844), .Y(n8341) );
  BUFX3 U1836 ( .A(n8873), .Y(n8399) );
  BUFX3 U1837 ( .A(n8774), .Y(n8224) );
  BUFX3 U1838 ( .A(n8803), .Y(n8282) );
  BUFX3 U1839 ( .A(n8832), .Y(n8340) );
  BUFX3 U1840 ( .A(n8861), .Y(n8398) );
  BUFX3 U1841 ( .A(n8669), .Y(n8014) );
  BUFX3 U1842 ( .A(n8701), .Y(n8075) );
  BUFX3 U1843 ( .A(n8729), .Y(n8131) );
  BUFX3 U1844 ( .A(n8669), .Y(n8015) );
  BUFX3 U1845 ( .A(n8669), .Y(n8013) );
  BUFX3 U1846 ( .A(n8701), .Y(n8074) );
  BUFX3 U1847 ( .A(n8729), .Y(n8130) );
  BUFX3 U1848 ( .A(n8701), .Y(n8073) );
  BUFX3 U1849 ( .A(n8729), .Y(n8129) );
  BUFX3 U1850 ( .A(n8778), .Y(n8228) );
  BUFX3 U1851 ( .A(n8807), .Y(n8286) );
  BUFX3 U1852 ( .A(n8836), .Y(n8344) );
  BUFX3 U1853 ( .A(n8865), .Y(n8402) );
  BUFX3 U1854 ( .A(n8778), .Y(n8227) );
  BUFX3 U1855 ( .A(n8807), .Y(n8285) );
  BUFX3 U1856 ( .A(n8836), .Y(n8343) );
  BUFX3 U1857 ( .A(n8865), .Y(n8401) );
  BUFX3 U1858 ( .A(n8670), .Y(n8018) );
  BUFX3 U1859 ( .A(n8670), .Y(n8017) );
  BUFX3 U1860 ( .A(n8702), .Y(n8078) );
  BUFX3 U1861 ( .A(n8730), .Y(n8134) );
  BUFX3 U1862 ( .A(n8670), .Y(n8016) );
  BUFX3 U1863 ( .A(n8702), .Y(n8077) );
  BUFX3 U1864 ( .A(n8730), .Y(n8133) );
  BUFX3 U1865 ( .A(n8702), .Y(n8076) );
  BUFX3 U1866 ( .A(n8730), .Y(n8132) );
  BUFX3 U1867 ( .A(n8671), .Y(n8021) );
  BUFX3 U1868 ( .A(n8703), .Y(n8079) );
  BUFX3 U1869 ( .A(n8731), .Y(n8135) );
  BUFX3 U1870 ( .A(n8779), .Y(n8231) );
  BUFX3 U1871 ( .A(n8808), .Y(n8289) );
  BUFX3 U1872 ( .A(n8837), .Y(n8347) );
  BUFX3 U1873 ( .A(n8866), .Y(n8405) );
  BUFX3 U1874 ( .A(n8671), .Y(n8020) );
  BUFX3 U1875 ( .A(n8703), .Y(n8081) );
  BUFX3 U1876 ( .A(n8731), .Y(n8137) );
  BUFX3 U1877 ( .A(n8779), .Y(n8230) );
  BUFX3 U1878 ( .A(n8808), .Y(n8288) );
  BUFX3 U1879 ( .A(n8837), .Y(n8346) );
  BUFX3 U1880 ( .A(n8866), .Y(n8404) );
  BUFX3 U1881 ( .A(n8775), .Y(n8216) );
  BUFX3 U1882 ( .A(n8804), .Y(n8274) );
  BUFX3 U1883 ( .A(n8833), .Y(n8332) );
  BUFX3 U1884 ( .A(n8862), .Y(n8390) );
  BUFX3 U1885 ( .A(n8775), .Y(n8215) );
  BUFX3 U1886 ( .A(n8804), .Y(n8273) );
  BUFX3 U1887 ( .A(n8833), .Y(n8331) );
  BUFX3 U1888 ( .A(n8862), .Y(n8389) );
  BUFX3 U1889 ( .A(n8666), .Y(n8006) );
  BUFX3 U1890 ( .A(n8666), .Y(n8005) );
  BUFX3 U1891 ( .A(n8698), .Y(n8066) );
  BUFX3 U1892 ( .A(n8726), .Y(n8122) );
  BUFX3 U1893 ( .A(n8666), .Y(n8004) );
  BUFX3 U1894 ( .A(n8698), .Y(n8065) );
  BUFX3 U1895 ( .A(n8726), .Y(n8121) );
  BUFX3 U1896 ( .A(n8698), .Y(n8064) );
  BUFX3 U1897 ( .A(n8726), .Y(n8120) );
  BUFX3 U1898 ( .A(n8776), .Y(n8219) );
  BUFX3 U1899 ( .A(n8805), .Y(n8277) );
  BUFX3 U1900 ( .A(n8834), .Y(n8335) );
  BUFX3 U1901 ( .A(n8863), .Y(n8393) );
  BUFX3 U1902 ( .A(n8776), .Y(n8218) );
  BUFX3 U1903 ( .A(n8805), .Y(n8276) );
  BUFX3 U1904 ( .A(n8834), .Y(n8334) );
  BUFX3 U1905 ( .A(n8863), .Y(n8392) );
  BUFX3 U1906 ( .A(n8667), .Y(n8009) );
  BUFX3 U1907 ( .A(n8667), .Y(n8008) );
  BUFX3 U1908 ( .A(n8699), .Y(n8069) );
  BUFX3 U1909 ( .A(n8727), .Y(n8125) );
  BUFX3 U1910 ( .A(n8667), .Y(n8007) );
  BUFX3 U1911 ( .A(n8699), .Y(n8068) );
  BUFX3 U1912 ( .A(n8727), .Y(n8124) );
  BUFX3 U1913 ( .A(n8699), .Y(n8067) );
  BUFX3 U1914 ( .A(n8727), .Y(n8123) );
  BUFX3 U1915 ( .A(n8668), .Y(n8011) );
  BUFX3 U1916 ( .A(n8700), .Y(n8072) );
  BUFX3 U1917 ( .A(n8728), .Y(n8128) );
  BUFX3 U1918 ( .A(n8777), .Y(n8221) );
  BUFX3 U1919 ( .A(n8806), .Y(n8279) );
  BUFX3 U1920 ( .A(n8835), .Y(n8337) );
  BUFX3 U1921 ( .A(n8864), .Y(n8395) );
  BUFX3 U1922 ( .A(n8668), .Y(n8010) );
  BUFX3 U1923 ( .A(n8700), .Y(n8071) );
  BUFX3 U1924 ( .A(n8728), .Y(n8127) );
  BUFX3 U1925 ( .A(n8668), .Y(n8012) );
  BUFX3 U1926 ( .A(n8700), .Y(n8070) );
  BUFX3 U1927 ( .A(n8728), .Y(n8126) );
  BUFX3 U1928 ( .A(n8777), .Y(n8222) );
  BUFX3 U1929 ( .A(n8806), .Y(n8280) );
  BUFX3 U1930 ( .A(n8835), .Y(n8338) );
  BUFX3 U1931 ( .A(n8864), .Y(n8396) );
  BUFX3 U1932 ( .A(n8671), .Y(n8019) );
  BUFX3 U1933 ( .A(n8703), .Y(n8080) );
  BUFX3 U1934 ( .A(n8731), .Y(n8136) );
  BUFX3 U1935 ( .A(n8782), .Y(n8241) );
  BUFX3 U1936 ( .A(n8811), .Y(n8299) );
  BUFX3 U1937 ( .A(n8840), .Y(n8357) );
  BUFX3 U1938 ( .A(n8869), .Y(n8415) );
  BUFX3 U1939 ( .A(n8783), .Y(n8244) );
  BUFX3 U1940 ( .A(n8812), .Y(n8302) );
  BUFX3 U1941 ( .A(n8841), .Y(n8360) );
  BUFX3 U1942 ( .A(n8870), .Y(n8418) );
  BUFX3 U1943 ( .A(n8780), .Y(n8235) );
  BUFX3 U1944 ( .A(n8809), .Y(n8293) );
  BUFX3 U1945 ( .A(n8838), .Y(n8351) );
  BUFX3 U1946 ( .A(n8867), .Y(n8409) );
  BUFX3 U1947 ( .A(n8781), .Y(n8238) );
  BUFX3 U1948 ( .A(n8810), .Y(n8296) );
  BUFX3 U1949 ( .A(n8839), .Y(n8354) );
  BUFX3 U1950 ( .A(n8868), .Y(n8412) );
  BUFX3 U1951 ( .A(n8788), .Y(n8258) );
  BUFX3 U1952 ( .A(n8817), .Y(n8316) );
  BUFX3 U1953 ( .A(n8846), .Y(n8374) );
  BUFX3 U1954 ( .A(n8875), .Y(n8432) );
  BUFX3 U1955 ( .A(n8784), .Y(n8247) );
  BUFX3 U1956 ( .A(n8813), .Y(n8305) );
  BUFX3 U1957 ( .A(n8842), .Y(n8363) );
  BUFX3 U1958 ( .A(n8871), .Y(n8421) );
  BUFX3 U1959 ( .A(n8785), .Y(n8250) );
  BUFX3 U1960 ( .A(n8814), .Y(n8308) );
  BUFX3 U1961 ( .A(n8843), .Y(n8366) );
  BUFX3 U1962 ( .A(n8872), .Y(n8424) );
  BUFX3 U1963 ( .A(n8786), .Y(n8253) );
  BUFX3 U1964 ( .A(n8815), .Y(n8311) );
  BUFX3 U1965 ( .A(n8844), .Y(n8369) );
  BUFX3 U1966 ( .A(n8873), .Y(n8427) );
  BUFX3 U1967 ( .A(n8778), .Y(n8211) );
  BUFX3 U1968 ( .A(n8807), .Y(n8269) );
  BUFX3 U1969 ( .A(n8836), .Y(n8327) );
  BUFX3 U1970 ( .A(n8865), .Y(n8385) );
  BUFX3 U1971 ( .A(n8774), .Y(n8214) );
  BUFX3 U1972 ( .A(n8803), .Y(n8272) );
  BUFX3 U1973 ( .A(n8832), .Y(n8330) );
  BUFX3 U1974 ( .A(n8861), .Y(n8388) );
  BUFX3 U1975 ( .A(n8787), .Y(n8206) );
  BUFX3 U1976 ( .A(n8816), .Y(n8264) );
  BUFX3 U1977 ( .A(n8845), .Y(n8322) );
  BUFX3 U1978 ( .A(n8874), .Y(n8380) );
  BUFX3 U1979 ( .A(n8788), .Y(n8209) );
  BUFX3 U1980 ( .A(n8817), .Y(n8267) );
  BUFX3 U1981 ( .A(n8846), .Y(n8325) );
  BUFX3 U1982 ( .A(n8875), .Y(n8383) );
  BUFX3 U1983 ( .A(n8787), .Y(n8226) );
  BUFX3 U1984 ( .A(n8816), .Y(n8284) );
  BUFX3 U1985 ( .A(n8845), .Y(n8342) );
  BUFX3 U1986 ( .A(n8874), .Y(n8400) );
  BUFX3 U1987 ( .A(n8778), .Y(n8229) );
  BUFX3 U1988 ( .A(n8807), .Y(n8287) );
  BUFX3 U1989 ( .A(n8836), .Y(n8345) );
  BUFX3 U1990 ( .A(n8865), .Y(n8403) );
  BUFX3 U1991 ( .A(n8775), .Y(n8217) );
  BUFX3 U1992 ( .A(n8804), .Y(n8275) );
  BUFX3 U1993 ( .A(n8833), .Y(n8333) );
  BUFX3 U1994 ( .A(n8862), .Y(n8391) );
  BUFX3 U1995 ( .A(n8776), .Y(n8220) );
  BUFX3 U1996 ( .A(n8805), .Y(n8278) );
  BUFX3 U1997 ( .A(n8834), .Y(n8336) );
  BUFX3 U1998 ( .A(n8863), .Y(n8394) );
  BUFX3 U1999 ( .A(n8777), .Y(n8223) );
  BUFX3 U2000 ( .A(n8806), .Y(n8281) );
  BUFX3 U2001 ( .A(n8835), .Y(n8339) );
  BUFX3 U2002 ( .A(n8864), .Y(n8397) );
  BUFX3 U2003 ( .A(n8779), .Y(n8232) );
  BUFX3 U2004 ( .A(n8808), .Y(n8290) );
  BUFX3 U2005 ( .A(n8837), .Y(n8348) );
  BUFX3 U2006 ( .A(n8866), .Y(n8406) );
  BUFX3 U2007 ( .A(n8783), .Y(n8260) );
  BUFX3 U2008 ( .A(n8812), .Y(n8318) );
  BUFX3 U2009 ( .A(n8841), .Y(n8376) );
  BUFX3 U2010 ( .A(n8870), .Y(n8434) );
  BUFX3 U2011 ( .A(n8780), .Y(n8259) );
  BUFX3 U2012 ( .A(n8809), .Y(n8317) );
  BUFX3 U2013 ( .A(n8838), .Y(n8375) );
  BUFX3 U2014 ( .A(n8867), .Y(n8433) );
  INVX1 U2015 ( .A(n8681), .Y(n8665) );
  INVX1 U2016 ( .A(n8711), .Y(n8694) );
  INVX1 U2017 ( .A(n8739), .Y(n8722) );
  INVX1 U2018 ( .A(n8764), .Y(n8750) );
  INVX1 U2019 ( .A(n8789), .Y(n8773) );
  INVX1 U2020 ( .A(n8818), .Y(n8802) );
  INVX1 U2021 ( .A(n8847), .Y(n8831) );
  INVX1 U2022 ( .A(n8876), .Y(n8860) );
  CLKINVX3 U2023 ( .A(n8641), .Y(n7993) );
  CLKINVX3 U2024 ( .A(n8641), .Y(n7992) );
  CLKINVX3 U2025 ( .A(n8650), .Y(n4649) );
  CLKINVX3 U2026 ( .A(n7989), .Y(n7990) );
  CLKINVX3 U2027 ( .A(n8650), .Y(n4648) );
  INVX1 U2028 ( .A(n7370), .Y(n7371) );
  INVX1 U2029 ( .A(n7370), .Y(n7372) );
  INVX1 U2030 ( .A(n7370), .Y(n7373) );
  INVX1 U2031 ( .A(n7622), .Y(n7620) );
  INVX1 U2032 ( .A(n7649), .Y(n7621) );
  INVX1 U2033 ( .A(n4279), .Y(n4297) );
  INVX1 U2034 ( .A(n4279), .Y(n4298) );
  INVX1 U2035 ( .A(n4285), .Y(n4299) );
  INVX1 U2036 ( .A(n4279), .Y(n4300) );
  INVX1 U2037 ( .A(n4276), .Y(n4285) );
  INVX1 U2038 ( .A(n4276), .Y(n4284) );
  INVX1 U2039 ( .A(n4276), .Y(n4283) );
  INVX1 U2040 ( .A(n4277), .Y(n4282) );
  INVX1 U2041 ( .A(n4277), .Y(n4281) );
  INVX1 U2042 ( .A(n4277), .Y(n4280) );
  INVX1 U2043 ( .A(N79), .Y(n7622) );
  INVX1 U2044 ( .A(n4026), .Y(n4031) );
  INVX1 U2045 ( .A(n4026), .Y(n4030) );
  INVX1 U2046 ( .A(N68), .Y(n4029) );
  INVX1 U2047 ( .A(n4026), .Y(n4028) );
  INVX1 U2048 ( .A(N68), .Y(n4027) );
  CLKINVX3 U2049 ( .A(n4636), .Y(n4645) );
  INVX1 U2050 ( .A(N73), .Y(n4636) );
  INVX1 U2051 ( .A(n4626), .Y(n4562) );
  INVX1 U2052 ( .A(n7969), .Y(n7905) );
  INVX1 U2053 ( .A(n4626), .Y(n4561) );
  INVX1 U2054 ( .A(n7968), .Y(n7904) );
  INVX1 U2055 ( .A(N72), .Y(n4627) );
  INVX1 U2056 ( .A(n7978), .Y(n7970) );
  INVX1 U2057 ( .A(N70), .Y(n4505) );
  INVX1 U2058 ( .A(n4560), .Y(n4504) );
  INVX1 U2059 ( .A(n7903), .Y(n7848) );
  INVX1 U2060 ( .A(n7903), .Y(n7847) );
  AND2X2 U2061 ( .A(n8635), .B(n1272), .Y(n391) );
  AND2X2 U2062 ( .A(n8629), .B(n1272), .Y(n392) );
  AND2X2 U2063 ( .A(n8626), .B(n1272), .Y(n393) );
  AND2X2 U2064 ( .A(n8612), .B(n8633), .Y(n394) );
  AND2X2 U2065 ( .A(n8609), .B(n8633), .Y(n395) );
  AND2X2 U2066 ( .A(n8605), .B(n8633), .Y(n396) );
  AND2X2 U2067 ( .A(n8602), .B(n8633), .Y(n397) );
  AND2X2 U2068 ( .A(n8600), .B(n8633), .Y(n398) );
  AND2X2 U2069 ( .A(n8597), .B(n8633), .Y(n399) );
  AND2X2 U2070 ( .A(n8594), .B(n8633), .Y(n400) );
  AND2X2 U2071 ( .A(n8591), .B(n8633), .Y(n401) );
  AND2X2 U2072 ( .A(n8587), .B(n8633), .Y(n402) );
  AND2X2 U2073 ( .A(n8585), .B(n8633), .Y(n403) );
  AND2X2 U2074 ( .A(n8581), .B(n8633), .Y(n404) );
  AND2X2 U2075 ( .A(n8578), .B(n8633), .Y(n405) );
  AND2X2 U2076 ( .A(n8575), .B(n8632), .Y(n406) );
  AND2X2 U2077 ( .A(n8572), .B(n8632), .Y(n407) );
  AND2X2 U2078 ( .A(n8569), .B(n8632), .Y(n408) );
  AND2X2 U2079 ( .A(n8566), .B(n8632), .Y(n409) );
  AND2X2 U2080 ( .A(n8563), .B(n8632), .Y(n410) );
  AND2X2 U2081 ( .A(n8561), .B(n8632), .Y(n411) );
  AND2X2 U2082 ( .A(n8557), .B(n8632), .Y(n412) );
  AND2X2 U2083 ( .A(n8554), .B(n8632), .Y(n413) );
  AND2X2 U2084 ( .A(n8551), .B(n8632), .Y(n414) );
  AND2X2 U2085 ( .A(n8548), .B(n8632), .Y(n415) );
  AND2X2 U2086 ( .A(n8545), .B(n8632), .Y(n416) );
  AND2X2 U2087 ( .A(n8542), .B(n8632), .Y(n417) );
  AND2X2 U2088 ( .A(n8540), .B(n8612), .Y(n418) );
  AND2X2 U2089 ( .A(n8540), .B(n8609), .Y(n419) );
  AND2X2 U2090 ( .A(n8540), .B(n8605), .Y(n420) );
  AND2X2 U2091 ( .A(n8540), .B(n8602), .Y(n421) );
  AND2X2 U2092 ( .A(n8540), .B(n8600), .Y(n422) );
  AND2X2 U2093 ( .A(n8540), .B(n8597), .Y(n423) );
  AND2X2 U2094 ( .A(n8540), .B(n8594), .Y(n424) );
  AND2X2 U2095 ( .A(n8540), .B(n8591), .Y(n425) );
  AND2X2 U2096 ( .A(n8540), .B(n8587), .Y(n426) );
  AND2X2 U2097 ( .A(n8540), .B(n8585), .Y(n427) );
  AND2X2 U2098 ( .A(n8540), .B(n8581), .Y(n428) );
  AND2X2 U2099 ( .A(n8540), .B(n8578), .Y(n429) );
  AND2X2 U2100 ( .A(n8539), .B(n8575), .Y(n430) );
  AND2X2 U2101 ( .A(n8539), .B(n8572), .Y(n431) );
  AND2X2 U2102 ( .A(n8539), .B(n8569), .Y(n432) );
  AND2X2 U2103 ( .A(n8539), .B(n8566), .Y(n433) );
  AND2X2 U2104 ( .A(n8539), .B(n8563), .Y(n434) );
  AND2X2 U2105 ( .A(n8539), .B(n8561), .Y(n435) );
  AND2X2 U2106 ( .A(n8539), .B(n8557), .Y(n436) );
  AND2X2 U2107 ( .A(n8539), .B(n8554), .Y(n437) );
  AND2X2 U2108 ( .A(n8539), .B(n8551), .Y(n438) );
  AND2X2 U2109 ( .A(n8539), .B(n8548), .Y(n439) );
  AND2X2 U2110 ( .A(n8539), .B(n8545), .Y(n440) );
  AND2X2 U2111 ( .A(n8539), .B(n8542), .Y(n441) );
  AND2X2 U2112 ( .A(n8537), .B(n8612), .Y(n442) );
  AND2X2 U2113 ( .A(n8537), .B(n8609), .Y(n443) );
  AND2X2 U2114 ( .A(n8537), .B(n8605), .Y(n444) );
  AND2X2 U2115 ( .A(n8537), .B(n8602), .Y(n445) );
  AND2X2 U2116 ( .A(n8537), .B(n8600), .Y(n446) );
  AND2X2 U2117 ( .A(n8537), .B(n8597), .Y(n447) );
  AND2X2 U2118 ( .A(n8537), .B(n8594), .Y(n448) );
  AND2X2 U2119 ( .A(n8537), .B(n8591), .Y(n449) );
  AND2X2 U2120 ( .A(n8537), .B(n8587), .Y(n450) );
  AND2X2 U2121 ( .A(n8537), .B(n8585), .Y(n451) );
  AND2X2 U2122 ( .A(n8537), .B(n8581), .Y(n452) );
  AND2X2 U2123 ( .A(n8537), .B(n8578), .Y(n453) );
  AND2X2 U2124 ( .A(n8536), .B(n8575), .Y(n454) );
  AND2X2 U2125 ( .A(n8536), .B(n8572), .Y(n455) );
  AND2X2 U2126 ( .A(n8536), .B(n8569), .Y(n456) );
  AND2X2 U2127 ( .A(n8536), .B(n8566), .Y(n457) );
  AND2X2 U2128 ( .A(n8536), .B(n8563), .Y(n458) );
  AND2X2 U2129 ( .A(n8536), .B(n8561), .Y(n459) );
  AND2X2 U2130 ( .A(n8536), .B(n8557), .Y(n460) );
  AND2X2 U2131 ( .A(n8536), .B(n8554), .Y(n461) );
  AND2X2 U2132 ( .A(n8536), .B(n8551), .Y(n462) );
  AND2X2 U2133 ( .A(n8536), .B(n8548), .Y(n463) );
  AND2X2 U2134 ( .A(n8536), .B(n8545), .Y(n464) );
  AND2X2 U2135 ( .A(n8536), .B(n8542), .Y(n465) );
  AND2X2 U2136 ( .A(n8534), .B(n8612), .Y(n466) );
  AND2X2 U2137 ( .A(n8534), .B(n8609), .Y(n467) );
  AND2X2 U2138 ( .A(n8534), .B(n8605), .Y(n468) );
  AND2X2 U2139 ( .A(n8534), .B(n8602), .Y(n469) );
  AND2X2 U2140 ( .A(n8534), .B(n8600), .Y(n470) );
  AND2X2 U2141 ( .A(n8534), .B(n8597), .Y(n471) );
  AND2X2 U2142 ( .A(n8534), .B(n8594), .Y(n472) );
  AND2X2 U2143 ( .A(n8534), .B(n8591), .Y(n473) );
  AND2X2 U2144 ( .A(n8534), .B(n8587), .Y(n474) );
  AND2X2 U2145 ( .A(n8534), .B(n8585), .Y(n475) );
  AND2X2 U2146 ( .A(n8534), .B(n8581), .Y(n476) );
  AND2X2 U2147 ( .A(n8534), .B(n8578), .Y(n477) );
  AND2X2 U2148 ( .A(n8533), .B(n8575), .Y(n478) );
  AND2X2 U2149 ( .A(n8533), .B(n8572), .Y(n479) );
  AND2X2 U2150 ( .A(n8533), .B(n8569), .Y(n480) );
  AND2X2 U2151 ( .A(n8533), .B(n8566), .Y(n481) );
  AND2X2 U2152 ( .A(n8533), .B(n8563), .Y(n482) );
  AND2X2 U2153 ( .A(n8533), .B(n8561), .Y(n483) );
  AND2X2 U2154 ( .A(n8533), .B(n8557), .Y(n484) );
  AND2X2 U2155 ( .A(n8533), .B(n8554), .Y(n485) );
  AND2X2 U2156 ( .A(n8533), .B(n8551), .Y(n486) );
  AND2X2 U2157 ( .A(n8533), .B(n8548), .Y(n487) );
  AND2X2 U2158 ( .A(n8533), .B(n8545), .Y(n488) );
  AND2X2 U2159 ( .A(n8533), .B(n8542), .Y(n489) );
  AND2X2 U2160 ( .A(n8531), .B(n8612), .Y(n490) );
  AND2X2 U2161 ( .A(n8531), .B(n8609), .Y(n491) );
  AND2X2 U2162 ( .A(n8531), .B(n8605), .Y(n492) );
  AND2X2 U2163 ( .A(n8531), .B(n8602), .Y(n493) );
  AND2X2 U2164 ( .A(n8531), .B(n8600), .Y(n494) );
  AND2X2 U2165 ( .A(n8531), .B(n8597), .Y(n495) );
  AND2X2 U2166 ( .A(n8531), .B(n8594), .Y(n496) );
  AND2X2 U2167 ( .A(n8531), .B(n8591), .Y(n497) );
  AND2X2 U2168 ( .A(n8531), .B(n8587), .Y(n498) );
  AND2X2 U2169 ( .A(n8531), .B(n8585), .Y(n499) );
  AND2X2 U2170 ( .A(n8531), .B(n8581), .Y(n500) );
  AND2X2 U2171 ( .A(n8531), .B(n8578), .Y(n501) );
  AND2X2 U2172 ( .A(n8530), .B(n8575), .Y(n502) );
  AND2X2 U2173 ( .A(n8530), .B(n8572), .Y(n503) );
  AND2X2 U2174 ( .A(n8530), .B(n8569), .Y(n504) );
  AND2X2 U2175 ( .A(n8530), .B(n8566), .Y(n505) );
  AND2X2 U2176 ( .A(n8530), .B(n8563), .Y(n506) );
  AND2X2 U2177 ( .A(n8530), .B(n8561), .Y(n507) );
  AND2X2 U2178 ( .A(n8530), .B(n8557), .Y(n508) );
  AND2X2 U2179 ( .A(n8530), .B(n8554), .Y(n509) );
  AND2X2 U2180 ( .A(n8530), .B(n8551), .Y(n510) );
  AND2X2 U2181 ( .A(n8530), .B(n8548), .Y(n511) );
  AND2X2 U2182 ( .A(n8530), .B(n8545), .Y(n512) );
  AND2X2 U2183 ( .A(n8530), .B(n8542), .Y(n513) );
  AND2X2 U2184 ( .A(n8528), .B(n8612), .Y(n514) );
  AND2X2 U2185 ( .A(n8528), .B(n8609), .Y(n515) );
  AND2X2 U2186 ( .A(n8528), .B(n8605), .Y(n516) );
  AND2X2 U2187 ( .A(n8528), .B(n8602), .Y(n517) );
  AND2X2 U2188 ( .A(n8528), .B(n8600), .Y(n518) );
  AND2X2 U2189 ( .A(n8528), .B(n8597), .Y(n519) );
  AND2X2 U2190 ( .A(n8528), .B(n8594), .Y(n520) );
  AND2X2 U2191 ( .A(n8528), .B(n8591), .Y(n521) );
  AND2X2 U2192 ( .A(n8528), .B(n8587), .Y(n522) );
  AND2X2 U2193 ( .A(n8528), .B(n8585), .Y(n523) );
  AND2X2 U2194 ( .A(n8528), .B(n8581), .Y(n524) );
  AND2X2 U2195 ( .A(n8528), .B(n8578), .Y(n525) );
  AND2X2 U2196 ( .A(n8527), .B(n8575), .Y(n526) );
  AND2X2 U2197 ( .A(n8527), .B(n8572), .Y(n527) );
  AND2X2 U2198 ( .A(n8527), .B(n8569), .Y(n528) );
  AND2X2 U2199 ( .A(n8527), .B(n8566), .Y(n529) );
  AND2X2 U2200 ( .A(n8527), .B(n8563), .Y(n530) );
  AND2X2 U2201 ( .A(n8527), .B(n8561), .Y(n531) );
  AND2X2 U2202 ( .A(n8527), .B(n8557), .Y(n532) );
  AND2X2 U2203 ( .A(n8527), .B(n8554), .Y(n533) );
  AND2X2 U2204 ( .A(n8527), .B(n8551), .Y(n534) );
  AND2X2 U2205 ( .A(n8527), .B(n8548), .Y(n535) );
  AND2X2 U2206 ( .A(n8527), .B(n8545), .Y(n536) );
  AND2X2 U2207 ( .A(n8527), .B(n8542), .Y(n537) );
  AND2X2 U2208 ( .A(n8525), .B(n8612), .Y(n538) );
  AND2X2 U2209 ( .A(n8525), .B(n8609), .Y(n539) );
  AND2X2 U2210 ( .A(n8525), .B(n8605), .Y(n540) );
  AND2X2 U2211 ( .A(n8525), .B(n8602), .Y(n541) );
  AND2X2 U2212 ( .A(n8525), .B(n8600), .Y(n542) );
  AND2X2 U2213 ( .A(n8525), .B(n8597), .Y(n543) );
  AND2X2 U2214 ( .A(n8525), .B(n8594), .Y(n544) );
  AND2X2 U2215 ( .A(n8525), .B(n8591), .Y(n545) );
  AND2X2 U2216 ( .A(n8525), .B(n8587), .Y(n546) );
  AND2X2 U2217 ( .A(n8525), .B(n8585), .Y(n547) );
  AND2X2 U2218 ( .A(n8525), .B(n8581), .Y(n548) );
  AND2X2 U2219 ( .A(n8525), .B(n8578), .Y(n549) );
  AND2X2 U2220 ( .A(n8524), .B(n8575), .Y(n550) );
  AND2X2 U2221 ( .A(n8524), .B(n8572), .Y(n551) );
  AND2X2 U2222 ( .A(n8524), .B(n8569), .Y(n552) );
  AND2X2 U2223 ( .A(n8524), .B(n8566), .Y(n553) );
  AND2X2 U2224 ( .A(n8524), .B(n8563), .Y(n554) );
  AND2X2 U2225 ( .A(n8524), .B(n8561), .Y(n555) );
  AND2X2 U2226 ( .A(n8524), .B(n8557), .Y(n556) );
  AND2X2 U2227 ( .A(n8524), .B(n8554), .Y(n557) );
  AND2X2 U2228 ( .A(n8524), .B(n8551), .Y(n558) );
  AND2X2 U2229 ( .A(n8524), .B(n8548), .Y(n559) );
  AND2X2 U2230 ( .A(n8524), .B(n8545), .Y(n560) );
  AND2X2 U2231 ( .A(n8524), .B(n8542), .Y(n561) );
  AND2X2 U2232 ( .A(n8522), .B(n1286), .Y(n562) );
  AND2X2 U2233 ( .A(n8522), .B(n1288), .Y(n563) );
  AND2X2 U2234 ( .A(n8522), .B(n8605), .Y(n564) );
  AND2X2 U2235 ( .A(n8522), .B(n8602), .Y(n565) );
  AND2X2 U2236 ( .A(n8522), .B(n1294), .Y(n566) );
  AND2X2 U2237 ( .A(n8522), .B(n1296), .Y(n567) );
  AND2X2 U2238 ( .A(n8522), .B(n1298), .Y(n568) );
  AND2X2 U2239 ( .A(n8522), .B(n1300), .Y(n569) );
  AND2X2 U2240 ( .A(n8522), .B(n8587), .Y(n570) );
  AND2X2 U2241 ( .A(n8522), .B(n1304), .Y(n571) );
  AND2X2 U2242 ( .A(n8522), .B(n8581), .Y(n572) );
  AND2X2 U2243 ( .A(n8522), .B(n8578), .Y(n573) );
  AND2X2 U2244 ( .A(n8521), .B(n8575), .Y(n574) );
  AND2X2 U2245 ( .A(n8521), .B(n8572), .Y(n575) );
  AND2X2 U2246 ( .A(n8521), .B(n8569), .Y(n576) );
  AND2X2 U2247 ( .A(n8521), .B(n8566), .Y(n577) );
  AND2X2 U2248 ( .A(n8521), .B(n8563), .Y(n578) );
  AND2X2 U2249 ( .A(n8521), .B(n1320), .Y(n579) );
  AND2X2 U2250 ( .A(n8521), .B(n8557), .Y(n580) );
  AND2X2 U2251 ( .A(n8521), .B(n8554), .Y(n581) );
  AND2X2 U2252 ( .A(n8521), .B(n8551), .Y(n582) );
  AND2X2 U2253 ( .A(n8521), .B(n8548), .Y(n583) );
  AND2X2 U2254 ( .A(n8521), .B(n8545), .Y(n584) );
  AND2X2 U2255 ( .A(n8521), .B(n8542), .Y(n585) );
  AND2X2 U2256 ( .A(n8519), .B(n1286), .Y(n586) );
  AND2X2 U2257 ( .A(n8519), .B(n1288), .Y(n587) );
  AND2X2 U2258 ( .A(n8519), .B(n8605), .Y(n588) );
  AND2X2 U2259 ( .A(n8519), .B(n8602), .Y(n589) );
  AND2X2 U2260 ( .A(n8519), .B(n1294), .Y(n590) );
  AND2X2 U2261 ( .A(n8519), .B(n1296), .Y(n591) );
  AND2X2 U2262 ( .A(n8519), .B(n1298), .Y(n592) );
  AND2X2 U2263 ( .A(n8519), .B(n1300), .Y(n593) );
  AND2X2 U2264 ( .A(n8519), .B(n8587), .Y(n594) );
  AND2X2 U2265 ( .A(n8519), .B(n1304), .Y(n595) );
  AND2X2 U2266 ( .A(n8519), .B(n8581), .Y(n596) );
  AND2X2 U2267 ( .A(n8519), .B(n8578), .Y(n597) );
  AND2X2 U2268 ( .A(n8518), .B(n8575), .Y(n598) );
  AND2X2 U2269 ( .A(n8518), .B(n8572), .Y(n599) );
  AND2X2 U2270 ( .A(n8518), .B(n8569), .Y(n600) );
  AND2X2 U2271 ( .A(n8518), .B(n8566), .Y(n601) );
  AND2X2 U2272 ( .A(n8518), .B(n8563), .Y(n602) );
  AND2X2 U2273 ( .A(n8518), .B(n1320), .Y(n603) );
  AND2X2 U2274 ( .A(n8518), .B(n8557), .Y(n604) );
  AND2X2 U2275 ( .A(n8518), .B(n8554), .Y(n605) );
  AND2X2 U2276 ( .A(n8518), .B(n8551), .Y(n606) );
  AND2X2 U2277 ( .A(n8518), .B(n8548), .Y(n607) );
  AND2X2 U2278 ( .A(n8518), .B(n8545), .Y(n608) );
  AND2X2 U2279 ( .A(n8518), .B(n8542), .Y(n609) );
  AND2X2 U2280 ( .A(n8516), .B(n1286), .Y(n610) );
  AND2X2 U2281 ( .A(n8516), .B(n1288), .Y(n611) );
  AND2X2 U2282 ( .A(n8516), .B(n8605), .Y(n612) );
  AND2X2 U2283 ( .A(n8516), .B(n8602), .Y(n613) );
  AND2X2 U2284 ( .A(n8516), .B(n1294), .Y(n614) );
  AND2X2 U2285 ( .A(n8516), .B(n1296), .Y(n615) );
  AND2X2 U2286 ( .A(n8516), .B(n1298), .Y(n616) );
  AND2X2 U2287 ( .A(n8516), .B(n1300), .Y(n617) );
  AND2X2 U2288 ( .A(n8516), .B(n8587), .Y(n618) );
  AND2X2 U2289 ( .A(n8516), .B(n1304), .Y(n619) );
  AND2X2 U2290 ( .A(n8516), .B(n8581), .Y(n620) );
  AND2X2 U2291 ( .A(n8516), .B(n8578), .Y(n621) );
  AND2X2 U2292 ( .A(n8515), .B(n8575), .Y(n622) );
  AND2X2 U2293 ( .A(n8515), .B(n8572), .Y(n623) );
  AND2X2 U2294 ( .A(n8515), .B(n8569), .Y(n624) );
  AND2X2 U2295 ( .A(n8515), .B(n8566), .Y(n625) );
  AND2X2 U2296 ( .A(n8515), .B(n8563), .Y(n626) );
  AND2X2 U2297 ( .A(n8515), .B(n1320), .Y(n627) );
  AND2X2 U2298 ( .A(n8515), .B(n8557), .Y(n628) );
  AND2X2 U2299 ( .A(n8515), .B(n8554), .Y(n629) );
  AND2X2 U2300 ( .A(n8515), .B(n8551), .Y(n630) );
  AND2X2 U2301 ( .A(n8515), .B(n8548), .Y(n631) );
  AND2X2 U2302 ( .A(n8515), .B(n8545), .Y(n632) );
  AND2X2 U2303 ( .A(n8515), .B(n8542), .Y(n633) );
  AND2X2 U2304 ( .A(n8513), .B(n1286), .Y(n634) );
  AND2X2 U2305 ( .A(n8513), .B(n1288), .Y(n635) );
  AND2X2 U2306 ( .A(n8513), .B(n8605), .Y(n636) );
  AND2X2 U2307 ( .A(n8513), .B(n8602), .Y(n637) );
  AND2X2 U2308 ( .A(n8513), .B(n1294), .Y(n638) );
  AND2X2 U2309 ( .A(n8513), .B(n1296), .Y(n639) );
  AND2X2 U2310 ( .A(n8513), .B(n1298), .Y(n640) );
  AND2X2 U2311 ( .A(n8513), .B(n1300), .Y(n641) );
  AND2X2 U2312 ( .A(n8513), .B(n8587), .Y(n642) );
  AND2X2 U2313 ( .A(n8513), .B(n1304), .Y(n643) );
  AND2X2 U2314 ( .A(n8513), .B(n8581), .Y(n644) );
  AND2X2 U2315 ( .A(n8513), .B(n8578), .Y(n645) );
  AND2X2 U2316 ( .A(n8512), .B(n8575), .Y(n646) );
  AND2X2 U2317 ( .A(n8512), .B(n8572), .Y(n647) );
  AND2X2 U2318 ( .A(n8512), .B(n8569), .Y(n648) );
  AND2X2 U2319 ( .A(n8512), .B(n8566), .Y(n649) );
  AND2X2 U2320 ( .A(n8512), .B(n8563), .Y(n650) );
  AND2X2 U2321 ( .A(n8512), .B(n1320), .Y(n651) );
  AND2X2 U2322 ( .A(n8512), .B(n8557), .Y(n652) );
  AND2X2 U2323 ( .A(n8512), .B(n8554), .Y(n653) );
  AND2X2 U2324 ( .A(n8512), .B(n8551), .Y(n654) );
  AND2X2 U2325 ( .A(n8512), .B(n8548), .Y(n655) );
  AND2X2 U2326 ( .A(n8512), .B(n8545), .Y(n656) );
  AND2X2 U2327 ( .A(n8512), .B(n8542), .Y(n657) );
  AND2X2 U2328 ( .A(n8510), .B(n1286), .Y(n658) );
  AND2X2 U2329 ( .A(n8510), .B(n1288), .Y(n659) );
  AND2X2 U2330 ( .A(n8510), .B(n8605), .Y(n660) );
  AND2X2 U2331 ( .A(n8510), .B(n8602), .Y(n661) );
  AND2X2 U2332 ( .A(n8510), .B(n1294), .Y(n662) );
  AND2X2 U2333 ( .A(n8510), .B(n1296), .Y(n663) );
  AND2X2 U2334 ( .A(n8510), .B(n1298), .Y(n664) );
  AND2X2 U2335 ( .A(n8510), .B(n1300), .Y(n665) );
  AND2X2 U2336 ( .A(n8510), .B(n8587), .Y(n666) );
  AND2X2 U2337 ( .A(n8510), .B(n1304), .Y(n667) );
  AND2X2 U2338 ( .A(n8510), .B(n8581), .Y(n668) );
  AND2X2 U2339 ( .A(n8510), .B(n8578), .Y(n669) );
  AND2X2 U2340 ( .A(n8509), .B(n8575), .Y(n670) );
  AND2X2 U2341 ( .A(n8509), .B(n8572), .Y(n671) );
  AND2X2 U2342 ( .A(n8509), .B(n8569), .Y(n672) );
  AND2X2 U2343 ( .A(n8509), .B(n8566), .Y(n673) );
  AND2X2 U2344 ( .A(n8509), .B(n8563), .Y(n674) );
  AND2X2 U2345 ( .A(n8509), .B(n1320), .Y(n675) );
  AND2X2 U2346 ( .A(n8509), .B(n8557), .Y(n676) );
  AND2X2 U2347 ( .A(n8509), .B(n8554), .Y(n677) );
  AND2X2 U2348 ( .A(n8509), .B(n8551), .Y(n678) );
  AND2X2 U2349 ( .A(n8509), .B(n8548), .Y(n679) );
  AND2X2 U2350 ( .A(n8509), .B(n8545), .Y(n680) );
  AND2X2 U2351 ( .A(n8509), .B(n8542), .Y(n681) );
  AND2X2 U2352 ( .A(n8507), .B(n1286), .Y(n682) );
  AND2X2 U2353 ( .A(n8507), .B(n1288), .Y(n683) );
  AND2X2 U2354 ( .A(n8507), .B(n8605), .Y(n684) );
  AND2X2 U2355 ( .A(n8507), .B(n8602), .Y(n685) );
  AND2X2 U2356 ( .A(n8507), .B(n1294), .Y(n686) );
  AND2X2 U2357 ( .A(n8507), .B(n1296), .Y(n687) );
  AND2X2 U2358 ( .A(n8507), .B(n1298), .Y(n688) );
  AND2X2 U2359 ( .A(n8507), .B(n1300), .Y(n689) );
  AND2X2 U2360 ( .A(n8507), .B(n8587), .Y(n690) );
  AND2X2 U2361 ( .A(n8507), .B(n1304), .Y(n691) );
  AND2X2 U2362 ( .A(n8507), .B(n8581), .Y(n692) );
  AND2X2 U2363 ( .A(n8507), .B(n8578), .Y(n693) );
  AND2X2 U2364 ( .A(n8506), .B(n8575), .Y(n694) );
  AND2X2 U2365 ( .A(n8506), .B(n8572), .Y(n695) );
  AND2X2 U2366 ( .A(n8506), .B(n8569), .Y(n696) );
  AND2X2 U2367 ( .A(n8506), .B(n8566), .Y(n697) );
  AND2X2 U2368 ( .A(n8506), .B(n8563), .Y(n698) );
  AND2X2 U2369 ( .A(n8506), .B(n1320), .Y(n699) );
  AND2X2 U2370 ( .A(n8506), .B(n8557), .Y(n700) );
  AND2X2 U2371 ( .A(n8506), .B(n8554), .Y(n701) );
  AND2X2 U2372 ( .A(n8506), .B(n8551), .Y(n702) );
  AND2X2 U2373 ( .A(n8506), .B(n8548), .Y(n703) );
  AND2X2 U2374 ( .A(n8506), .B(n8545), .Y(n704) );
  AND2X2 U2375 ( .A(n8506), .B(n8542), .Y(n705) );
  AND2X2 U2376 ( .A(n8503), .B(n8576), .Y(n706) );
  AND2X2 U2377 ( .A(n8503), .B(n8573), .Y(n707) );
  AND2X2 U2378 ( .A(n8503), .B(n8570), .Y(n708) );
  AND2X2 U2379 ( .A(n8503), .B(n8567), .Y(n709) );
  AND2X2 U2380 ( .A(n8503), .B(n8564), .Y(n710) );
  AND2X2 U2381 ( .A(n8503), .B(n8560), .Y(n711) );
  AND2X2 U2382 ( .A(n8503), .B(n8558), .Y(n712) );
  AND2X2 U2383 ( .A(n8503), .B(n8555), .Y(n713) );
  AND2X2 U2384 ( .A(n8503), .B(n8552), .Y(n714) );
  AND2X2 U2385 ( .A(n8503), .B(n8549), .Y(n715) );
  AND2X2 U2386 ( .A(n8503), .B(n8546), .Y(n716) );
  AND2X2 U2387 ( .A(n8503), .B(n8543), .Y(n717) );
  AND2X2 U2388 ( .A(n8500), .B(n8576), .Y(n718) );
  AND2X2 U2389 ( .A(n8500), .B(n8573), .Y(n719) );
  AND2X2 U2390 ( .A(n8500), .B(n8570), .Y(n720) );
  AND2X2 U2391 ( .A(n8500), .B(n8567), .Y(n721) );
  AND2X2 U2392 ( .A(n8500), .B(n8564), .Y(n722) );
  AND2X2 U2393 ( .A(n8500), .B(n8560), .Y(n723) );
  AND2X2 U2394 ( .A(n8500), .B(n8558), .Y(n724) );
  AND2X2 U2395 ( .A(n8500), .B(n8555), .Y(n725) );
  AND2X2 U2396 ( .A(n8500), .B(n8552), .Y(n726) );
  AND2X2 U2397 ( .A(n8500), .B(n8549), .Y(n727) );
  AND2X2 U2398 ( .A(n8500), .B(n8546), .Y(n728) );
  AND2X2 U2399 ( .A(n8500), .B(n8543), .Y(n729) );
  AND2X2 U2400 ( .A(n8497), .B(n8576), .Y(n730) );
  AND2X2 U2401 ( .A(n8497), .B(n8573), .Y(n731) );
  AND2X2 U2402 ( .A(n8497), .B(n8570), .Y(n732) );
  AND2X2 U2403 ( .A(n8497), .B(n8567), .Y(n733) );
  AND2X2 U2404 ( .A(n8497), .B(n8564), .Y(n734) );
  AND2X2 U2405 ( .A(n8497), .B(n8560), .Y(n735) );
  AND2X2 U2406 ( .A(n8497), .B(n8558), .Y(n736) );
  AND2X2 U2407 ( .A(n8497), .B(n8555), .Y(n737) );
  AND2X2 U2408 ( .A(n8497), .B(n8552), .Y(n738) );
  AND2X2 U2409 ( .A(n8497), .B(n8549), .Y(n739) );
  AND2X2 U2410 ( .A(n8497), .B(n8546), .Y(n740) );
  AND2X2 U2411 ( .A(n8497), .B(n8543), .Y(n741) );
  AND2X2 U2412 ( .A(n8494), .B(n8576), .Y(n742) );
  AND2X2 U2413 ( .A(n8494), .B(n8573), .Y(n743) );
  AND2X2 U2414 ( .A(n8494), .B(n8570), .Y(n744) );
  AND2X2 U2415 ( .A(n8494), .B(n8567), .Y(n745) );
  AND2X2 U2416 ( .A(n8494), .B(n8564), .Y(n746) );
  AND2X2 U2417 ( .A(n8494), .B(n8560), .Y(n747) );
  AND2X2 U2418 ( .A(n8494), .B(n8558), .Y(n748) );
  AND2X2 U2419 ( .A(n8494), .B(n8555), .Y(n749) );
  AND2X2 U2420 ( .A(n8494), .B(n8552), .Y(n750) );
  AND2X2 U2421 ( .A(n8494), .B(n8549), .Y(n751) );
  AND2X2 U2422 ( .A(n8494), .B(n8546), .Y(n752) );
  AND2X2 U2423 ( .A(n8494), .B(n8543), .Y(n753) );
  AND2X2 U2424 ( .A(n8491), .B(n8576), .Y(n754) );
  AND2X2 U2425 ( .A(n8491), .B(n8573), .Y(n755) );
  AND2X2 U2426 ( .A(n8491), .B(n8570), .Y(n756) );
  AND2X2 U2427 ( .A(n8491), .B(n8567), .Y(n757) );
  AND2X2 U2428 ( .A(n8491), .B(n8564), .Y(n758) );
  AND2X2 U2429 ( .A(n8491), .B(n8560), .Y(n759) );
  AND2X2 U2430 ( .A(n8491), .B(n8558), .Y(n760) );
  AND2X2 U2431 ( .A(n8491), .B(n8555), .Y(n761) );
  AND2X2 U2432 ( .A(n8491), .B(n8552), .Y(n762) );
  AND2X2 U2433 ( .A(n8491), .B(n8549), .Y(n763) );
  AND2X2 U2434 ( .A(n8491), .B(n8546), .Y(n764) );
  AND2X2 U2435 ( .A(n8491), .B(n8543), .Y(n765) );
  AND2X2 U2436 ( .A(n8488), .B(n8576), .Y(n766) );
  AND2X2 U2437 ( .A(n8488), .B(n8573), .Y(n767) );
  AND2X2 U2438 ( .A(n8488), .B(n8570), .Y(n768) );
  AND2X2 U2439 ( .A(n8488), .B(n8567), .Y(n769) );
  AND2X2 U2440 ( .A(n8488), .B(n8564), .Y(n770) );
  AND2X2 U2441 ( .A(n8488), .B(n8560), .Y(n771) );
  AND2X2 U2442 ( .A(n8488), .B(n8558), .Y(n772) );
  AND2X2 U2443 ( .A(n8488), .B(n8555), .Y(n773) );
  AND2X2 U2444 ( .A(n8488), .B(n8552), .Y(n774) );
  AND2X2 U2445 ( .A(n8488), .B(n8549), .Y(n775) );
  AND2X2 U2446 ( .A(n8488), .B(n8546), .Y(n776) );
  AND2X2 U2447 ( .A(n8488), .B(n8543), .Y(n777) );
  AND2X2 U2448 ( .A(n8485), .B(n8576), .Y(n778) );
  AND2X2 U2449 ( .A(n8485), .B(n8573), .Y(n779) );
  AND2X2 U2450 ( .A(n8485), .B(n8570), .Y(n780) );
  AND2X2 U2451 ( .A(n8485), .B(n8567), .Y(n781) );
  AND2X2 U2452 ( .A(n8485), .B(n8564), .Y(n782) );
  AND2X2 U2453 ( .A(n8485), .B(n8560), .Y(n783) );
  AND2X2 U2454 ( .A(n8485), .B(n8558), .Y(n784) );
  AND2X2 U2455 ( .A(n8485), .B(n8555), .Y(n785) );
  AND2X2 U2456 ( .A(n8485), .B(n8552), .Y(n786) );
  AND2X2 U2457 ( .A(n8485), .B(n8549), .Y(n787) );
  AND2X2 U2458 ( .A(n8485), .B(n8546), .Y(n788) );
  AND2X2 U2459 ( .A(n8485), .B(n8543), .Y(n789) );
  AND2X2 U2460 ( .A(n8482), .B(n8576), .Y(n790) );
  AND2X2 U2461 ( .A(n8482), .B(n8573), .Y(n791) );
  AND2X2 U2462 ( .A(n8482), .B(n8570), .Y(n792) );
  AND2X2 U2463 ( .A(n8482), .B(n8567), .Y(n793) );
  AND2X2 U2464 ( .A(n8482), .B(n8564), .Y(n794) );
  AND2X2 U2465 ( .A(n8482), .B(n8560), .Y(n795) );
  AND2X2 U2466 ( .A(n8482), .B(n8558), .Y(n796) );
  AND2X2 U2467 ( .A(n8482), .B(n8555), .Y(n797) );
  AND2X2 U2468 ( .A(n8482), .B(n8552), .Y(n798) );
  AND2X2 U2469 ( .A(n8482), .B(n8549), .Y(n799) );
  AND2X2 U2470 ( .A(n8482), .B(n8546), .Y(n800) );
  AND2X2 U2471 ( .A(n8482), .B(n8543), .Y(n801) );
  AND2X2 U2472 ( .A(n8479), .B(n8576), .Y(n802) );
  AND2X2 U2473 ( .A(n8479), .B(n8573), .Y(n803) );
  AND2X2 U2474 ( .A(n8479), .B(n8570), .Y(n804) );
  AND2X2 U2475 ( .A(n8479), .B(n8567), .Y(n805) );
  AND2X2 U2476 ( .A(n8479), .B(n8564), .Y(n806) );
  AND2X2 U2477 ( .A(n8479), .B(n8560), .Y(n807) );
  AND2X2 U2478 ( .A(n8479), .B(n8558), .Y(n808) );
  AND2X2 U2479 ( .A(n8479), .B(n8555), .Y(n809) );
  AND2X2 U2480 ( .A(n8479), .B(n8552), .Y(n810) );
  AND2X2 U2481 ( .A(n8479), .B(n8549), .Y(n811) );
  AND2X2 U2482 ( .A(n8479), .B(n8546), .Y(n812) );
  AND2X2 U2483 ( .A(n8479), .B(n8543), .Y(n813) );
  AND2X2 U2484 ( .A(n8476), .B(n8576), .Y(n814) );
  AND2X2 U2485 ( .A(n8476), .B(n8573), .Y(n815) );
  AND2X2 U2486 ( .A(n8476), .B(n8570), .Y(n816) );
  AND2X2 U2487 ( .A(n8476), .B(n8567), .Y(n817) );
  AND2X2 U2488 ( .A(n8476), .B(n8564), .Y(n818) );
  AND2X2 U2489 ( .A(n8476), .B(n8560), .Y(n819) );
  AND2X2 U2490 ( .A(n8476), .B(n8558), .Y(n820) );
  AND2X2 U2491 ( .A(n8476), .B(n8555), .Y(n821) );
  AND2X2 U2492 ( .A(n8476), .B(n8552), .Y(n822) );
  AND2X2 U2493 ( .A(n8476), .B(n8549), .Y(n823) );
  AND2X2 U2494 ( .A(n8476), .B(n8546), .Y(n824) );
  AND2X2 U2495 ( .A(n8476), .B(n8543), .Y(n825) );
  AND2X2 U2496 ( .A(n8473), .B(n8576), .Y(n826) );
  AND2X2 U2497 ( .A(n8473), .B(n8573), .Y(n827) );
  AND2X2 U2498 ( .A(n8473), .B(n8570), .Y(n828) );
  AND2X2 U2499 ( .A(n8473), .B(n8567), .Y(n829) );
  AND2X2 U2500 ( .A(n8473), .B(n8564), .Y(n830) );
  AND2X2 U2501 ( .A(n8473), .B(n8560), .Y(n831) );
  AND2X2 U2502 ( .A(n8473), .B(n8558), .Y(n832) );
  AND2X2 U2503 ( .A(n8473), .B(n8555), .Y(n833) );
  AND2X2 U2504 ( .A(n8473), .B(n8552), .Y(n834) );
  AND2X2 U2505 ( .A(n8473), .B(n8549), .Y(n835) );
  AND2X2 U2506 ( .A(n8473), .B(n8546), .Y(n836) );
  AND2X2 U2507 ( .A(n8473), .B(n8543), .Y(n837) );
  AND2X2 U2508 ( .A(n8470), .B(n8576), .Y(n838) );
  AND2X2 U2509 ( .A(n8470), .B(n8573), .Y(n839) );
  AND2X2 U2510 ( .A(n8470), .B(n8570), .Y(n840) );
  AND2X2 U2511 ( .A(n8470), .B(n8567), .Y(n841) );
  AND2X2 U2512 ( .A(n8470), .B(n8564), .Y(n842) );
  AND2X2 U2513 ( .A(n8470), .B(n8560), .Y(n843) );
  AND2X2 U2514 ( .A(n8470), .B(n8558), .Y(n844) );
  AND2X2 U2515 ( .A(n8470), .B(n8555), .Y(n845) );
  AND2X2 U2516 ( .A(n8470), .B(n8552), .Y(n846) );
  AND2X2 U2517 ( .A(n8470), .B(n8549), .Y(n847) );
  AND2X2 U2518 ( .A(n8470), .B(n8546), .Y(n848) );
  AND2X2 U2519 ( .A(n8470), .B(n8543), .Y(n849) );
  AND2X2 U2520 ( .A(n8467), .B(n8576), .Y(n850) );
  AND2X2 U2521 ( .A(n8467), .B(n8573), .Y(n851) );
  AND2X2 U2522 ( .A(n8467), .B(n8570), .Y(n852) );
  AND2X2 U2523 ( .A(n8467), .B(n8567), .Y(n853) );
  AND2X2 U2524 ( .A(n8467), .B(n8564), .Y(n854) );
  AND2X2 U2525 ( .A(n8467), .B(n8560), .Y(n855) );
  AND2X2 U2526 ( .A(n8467), .B(n8558), .Y(n856) );
  AND2X2 U2527 ( .A(n8467), .B(n8555), .Y(n857) );
  AND2X2 U2528 ( .A(n8467), .B(n8552), .Y(n858) );
  AND2X2 U2529 ( .A(n8467), .B(n8549), .Y(n859) );
  AND2X2 U2530 ( .A(n8467), .B(n8546), .Y(n860) );
  AND2X2 U2531 ( .A(n8467), .B(n8543), .Y(n861) );
  AND2X2 U2532 ( .A(n8464), .B(n8576), .Y(n862) );
  AND2X2 U2533 ( .A(n8464), .B(n8573), .Y(n863) );
  AND2X2 U2534 ( .A(n8464), .B(n8570), .Y(n864) );
  AND2X2 U2535 ( .A(n8464), .B(n8567), .Y(n865) );
  AND2X2 U2536 ( .A(n8464), .B(n8564), .Y(n866) );
  AND2X2 U2537 ( .A(n8464), .B(n8561), .Y(n867) );
  AND2X2 U2538 ( .A(n8464), .B(n8558), .Y(n868) );
  AND2X2 U2539 ( .A(n8464), .B(n8555), .Y(n869) );
  AND2X2 U2540 ( .A(n8464), .B(n8552), .Y(n870) );
  AND2X2 U2541 ( .A(n8464), .B(n8549), .Y(n871) );
  AND2X2 U2542 ( .A(n8464), .B(n8546), .Y(n872) );
  AND2X2 U2543 ( .A(n8464), .B(n8543), .Y(n873) );
  AND2X2 U2544 ( .A(n8461), .B(n1310), .Y(n874) );
  AND2X2 U2545 ( .A(n8461), .B(n1312), .Y(n875) );
  AND2X2 U2546 ( .A(n8461), .B(n1314), .Y(n876) );
  AND2X2 U2547 ( .A(n8461), .B(n1316), .Y(n877) );
  AND2X2 U2548 ( .A(n8461), .B(n1318), .Y(n878) );
  AND2X2 U2549 ( .A(n8461), .B(n8561), .Y(n879) );
  AND2X2 U2550 ( .A(n8461), .B(n1322), .Y(n880) );
  AND2X2 U2551 ( .A(n8461), .B(n1324), .Y(n881) );
  AND2X2 U2552 ( .A(n8461), .B(n1326), .Y(n882) );
  AND2X2 U2553 ( .A(n8461), .B(n1328), .Y(n883) );
  AND2X2 U2554 ( .A(n8461), .B(n1330), .Y(n884) );
  AND2X2 U2555 ( .A(n8461), .B(n1332), .Y(n885) );
  AND2X2 U2556 ( .A(n8458), .B(n1310), .Y(n886) );
  AND2X2 U2557 ( .A(n8458), .B(n1312), .Y(n887) );
  AND2X2 U2558 ( .A(n8458), .B(n1314), .Y(n888) );
  AND2X2 U2559 ( .A(n8458), .B(n1316), .Y(n889) );
  AND2X2 U2560 ( .A(n8458), .B(n1318), .Y(n890) );
  AND2X2 U2561 ( .A(n8458), .B(n8561), .Y(n891) );
  AND2X2 U2562 ( .A(n8458), .B(n1322), .Y(n892) );
  AND2X2 U2563 ( .A(n8458), .B(n1324), .Y(n893) );
  AND2X2 U2564 ( .A(n8458), .B(n1326), .Y(n894) );
  AND2X2 U2565 ( .A(n8458), .B(n1328), .Y(n895) );
  AND2X2 U2566 ( .A(n8458), .B(n1330), .Y(n896) );
  AND2X2 U2567 ( .A(n8458), .B(n1332), .Y(n897) );
  AND2X2 U2568 ( .A(n8455), .B(n1310), .Y(n898) );
  AND2X2 U2569 ( .A(n8455), .B(n1312), .Y(n899) );
  AND2X2 U2570 ( .A(n8455), .B(n1314), .Y(n900) );
  AND2X2 U2571 ( .A(n8455), .B(n1316), .Y(n901) );
  AND2X2 U2572 ( .A(n8455), .B(n1318), .Y(n902) );
  AND2X2 U2573 ( .A(n8455), .B(n8561), .Y(n903) );
  AND2X2 U2574 ( .A(n8455), .B(n1322), .Y(n904) );
  AND2X2 U2575 ( .A(n8455), .B(n1324), .Y(n905) );
  AND2X2 U2576 ( .A(n8455), .B(n1326), .Y(n906) );
  AND2X2 U2577 ( .A(n8455), .B(n1328), .Y(n907) );
  AND2X2 U2578 ( .A(n8455), .B(n1330), .Y(n908) );
  AND2X2 U2579 ( .A(n8455), .B(n1332), .Y(n909) );
  AND2X2 U2580 ( .A(n8452), .B(n1310), .Y(n910) );
  AND2X2 U2581 ( .A(n8452), .B(n1312), .Y(n911) );
  AND2X2 U2582 ( .A(n8452), .B(n1314), .Y(n912) );
  AND2X2 U2583 ( .A(n8452), .B(n1316), .Y(n913) );
  AND2X2 U2584 ( .A(n8452), .B(n1318), .Y(n914) );
  AND2X2 U2585 ( .A(n8452), .B(n8561), .Y(n915) );
  AND2X2 U2586 ( .A(n8452), .B(n1322), .Y(n916) );
  AND2X2 U2587 ( .A(n8452), .B(n1324), .Y(n917) );
  AND2X2 U2588 ( .A(n8452), .B(n1326), .Y(n918) );
  AND2X2 U2589 ( .A(n8452), .B(n1328), .Y(n919) );
  AND2X2 U2590 ( .A(n8452), .B(n1330), .Y(n920) );
  AND2X2 U2591 ( .A(n8452), .B(n1332), .Y(n921) );
  AND2X2 U2592 ( .A(n8449), .B(n1310), .Y(n922) );
  AND2X2 U2593 ( .A(n8449), .B(n1312), .Y(n923) );
  AND2X2 U2594 ( .A(n8449), .B(n1314), .Y(n924) );
  AND2X2 U2595 ( .A(n8449), .B(n1316), .Y(n925) );
  AND2X2 U2596 ( .A(n8449), .B(n1318), .Y(n926) );
  AND2X2 U2597 ( .A(n8449), .B(n8561), .Y(n927) );
  AND2X2 U2598 ( .A(n8449), .B(n1322), .Y(n928) );
  AND2X2 U2599 ( .A(n8449), .B(n1324), .Y(n929) );
  AND2X2 U2600 ( .A(n8449), .B(n1326), .Y(n930) );
  AND2X2 U2601 ( .A(n8449), .B(n1328), .Y(n931) );
  AND2X2 U2602 ( .A(n8449), .B(n1330), .Y(n932) );
  AND2X2 U2603 ( .A(n8449), .B(n1332), .Y(n933) );
  AND2X2 U2604 ( .A(n1334), .B(n8635), .Y(n934) );
  AND2X2 U2605 ( .A(n1334), .B(n8629), .Y(n935) );
  AND2X2 U2606 ( .A(n1334), .B(n8626), .Y(n936) );
  AND2X2 U2607 ( .A(n1334), .B(n8623), .Y(n937) );
  AND2X2 U2608 ( .A(n1334), .B(n8620), .Y(n938) );
  AND2X2 U2609 ( .A(n1334), .B(n8617), .Y(n939) );
  AND2X2 U2610 ( .A(n1334), .B(n8614), .Y(n940) );
  AND2X2 U2611 ( .A(n1369), .B(n8635), .Y(n941) );
  AND2X2 U2612 ( .A(n1369), .B(n8629), .Y(n942) );
  AND2X2 U2613 ( .A(n1369), .B(n8626), .Y(n943) );
  AND2X2 U2614 ( .A(n1369), .B(n8623), .Y(n944) );
  AND2X2 U2615 ( .A(n1369), .B(n8620), .Y(n945) );
  AND2X2 U2616 ( .A(n1369), .B(n8617), .Y(n946) );
  AND2X2 U2617 ( .A(n1369), .B(n8614), .Y(n947) );
  AND2X2 U2618 ( .A(n1403), .B(n8635), .Y(n948) );
  AND2X2 U2619 ( .A(n1403), .B(n8629), .Y(n949) );
  AND2X2 U2620 ( .A(n1403), .B(n8626), .Y(n950) );
  AND2X2 U2621 ( .A(n1403), .B(n8623), .Y(n951) );
  AND2X2 U2622 ( .A(n1403), .B(n8620), .Y(n952) );
  AND2X2 U2623 ( .A(n1403), .B(n8617), .Y(n953) );
  AND2X2 U2624 ( .A(n1403), .B(n8614), .Y(n954) );
  AND2X2 U2625 ( .A(n1437), .B(n8635), .Y(n955) );
  AND2X2 U2626 ( .A(n1437), .B(n8629), .Y(n956) );
  AND2X2 U2627 ( .A(n1437), .B(n8626), .Y(n957) );
  AND2X2 U2628 ( .A(n1471), .B(n8635), .Y(n958) );
  AND2X2 U2629 ( .A(n1471), .B(n8629), .Y(n959) );
  AND2X2 U2630 ( .A(n1471), .B(n8626), .Y(n960) );
  AND2X2 U2631 ( .A(n1505), .B(n8635), .Y(n961) );
  AND2X2 U2632 ( .A(n1505), .B(n8629), .Y(n962) );
  AND2X2 U2633 ( .A(n1505), .B(n8626), .Y(n963) );
  AND2X2 U2634 ( .A(n1539), .B(n8635), .Y(n964) );
  AND2X2 U2635 ( .A(n1539), .B(n8629), .Y(n965) );
  AND2X2 U2636 ( .A(n1539), .B(n8626), .Y(n966) );
  AND2X2 U2637 ( .A(n1573), .B(n8635), .Y(n967) );
  AND2X2 U2638 ( .A(n1573), .B(n8629), .Y(n968) );
  AND2X2 U2639 ( .A(n1573), .B(n8626), .Y(n969) );
  AND2X2 U2640 ( .A(n1573), .B(n8623), .Y(n970) );
  AND2X2 U2641 ( .A(n1573), .B(n8620), .Y(n971) );
  AND2X2 U2642 ( .A(n1573), .B(n8617), .Y(n972) );
  AND2X2 U2643 ( .A(n1573), .B(n8614), .Y(n973) );
  AND2X2 U2644 ( .A(n1608), .B(n8635), .Y(n974) );
  AND2X2 U2645 ( .A(n1608), .B(n8629), .Y(n975) );
  AND2X2 U2646 ( .A(n1608), .B(n8626), .Y(n976) );
  AND2X2 U2647 ( .A(n1608), .B(n8623), .Y(n977) );
  AND2X2 U2648 ( .A(n1608), .B(n8620), .Y(n978) );
  AND2X2 U2649 ( .A(n1608), .B(n8617), .Y(n979) );
  AND2X2 U2650 ( .A(n1608), .B(n8614), .Y(n980) );
  AND2X2 U2651 ( .A(n1641), .B(n8635), .Y(n981) );
  AND2X2 U2652 ( .A(n1641), .B(n8629), .Y(n982) );
  AND2X2 U2653 ( .A(n1641), .B(n8626), .Y(n983) );
  AND2X2 U2654 ( .A(n1641), .B(n8623), .Y(n984) );
  AND2X2 U2655 ( .A(n1641), .B(n8620), .Y(n985) );
  AND2X2 U2656 ( .A(n1641), .B(n8617), .Y(n986) );
  AND2X2 U2657 ( .A(n1641), .B(n8614), .Y(n987) );
  AND2X2 U2658 ( .A(n1674), .B(n8635), .Y(n988) );
  AND2X2 U2659 ( .A(n1674), .B(n8629), .Y(n989) );
  AND2X2 U2660 ( .A(n1674), .B(n8626), .Y(n990) );
  AND2X2 U2661 ( .A(n1674), .B(n8623), .Y(n991) );
  AND2X2 U2662 ( .A(n1674), .B(n8620), .Y(n992) );
  AND2X2 U2663 ( .A(n1674), .B(n8617), .Y(n993) );
  AND2X2 U2664 ( .A(n1674), .B(n8614), .Y(n994) );
  AND2X2 U2665 ( .A(n1707), .B(n8635), .Y(n995) );
  AND2X2 U2666 ( .A(n1707), .B(n8629), .Y(n996) );
  AND2X2 U2667 ( .A(n1707), .B(n8626), .Y(n997) );
  AND2X2 U2668 ( .A(n1707), .B(n8623), .Y(n998) );
  AND2X2 U2669 ( .A(n1707), .B(n8620), .Y(n999) );
  AND2X2 U2670 ( .A(n1707), .B(n8617), .Y(n1000) );
  AND2X2 U2671 ( .A(n1707), .B(n8614), .Y(n1001) );
  AND2X2 U2672 ( .A(n1972), .B(n8638), .Y(n1002) );
  AND2X2 U2673 ( .A(n2005), .B(n8638), .Y(n1003) );
  AND2X2 U2674 ( .A(n2038), .B(n8638), .Y(n1004) );
  AND2X2 U2675 ( .A(n2071), .B(n8638), .Y(n1005) );
  AND2X2 U2676 ( .A(n2104), .B(n8638), .Y(n1006) );
  AND2X2 U2677 ( .A(n2138), .B(n1268), .Y(n1007) );
  AND2X2 U2678 ( .A(n2171), .B(n1268), .Y(n1008) );
  AND2X2 U2679 ( .A(n2204), .B(n1268), .Y(n1009) );
  AND2X2 U2680 ( .A(n2237), .B(n1268), .Y(n1010) );
  AND2X2 U2681 ( .A(n2270), .B(n1268), .Y(n1011) );
  AND2X2 U2682 ( .A(n2303), .B(n1268), .Y(n1012) );
  AND2X2 U2683 ( .A(n2336), .B(n1268), .Y(n1013) );
  CLKINVX3 U2684 ( .A(n8637), .Y(n8636) );
  CLKINVX3 U2685 ( .A(n8631), .Y(n8630) );
  CLKINVX3 U2686 ( .A(n8628), .Y(n8627) );
  CLKINVX3 U2687 ( .A(n8613), .Y(n8611) );
  CLKINVX3 U2688 ( .A(n8610), .Y(n8608) );
  CLKINVX3 U2689 ( .A(n8607), .Y(n8606) );
  CLKINVX3 U2690 ( .A(n8604), .Y(n8603) );
  CLKINVX3 U2691 ( .A(n8601), .Y(n8599) );
  CLKINVX3 U2692 ( .A(n8598), .Y(n8596) );
  CLKINVX3 U2693 ( .A(n8595), .Y(n8593) );
  CLKINVX3 U2694 ( .A(n8592), .Y(n8590) );
  CLKINVX3 U2695 ( .A(n8589), .Y(n8588) );
  CLKINVX3 U2696 ( .A(n8586), .Y(n8584) );
  CLKINVX3 U2697 ( .A(n8583), .Y(n8582) );
  CLKINVX3 U2698 ( .A(n8580), .Y(n8579) );
  CLKINVX3 U2699 ( .A(n8577), .Y(n8576) );
  CLKINVX3 U2700 ( .A(n8574), .Y(n8573) );
  CLKINVX3 U2701 ( .A(n8571), .Y(n8570) );
  CLKINVX3 U2702 ( .A(n8568), .Y(n8567) );
  CLKINVX3 U2703 ( .A(n8565), .Y(n8564) );
  CLKINVX3 U2704 ( .A(n8562), .Y(n8560) );
  CLKINVX3 U2705 ( .A(n8559), .Y(n8558) );
  CLKINVX3 U2706 ( .A(n8556), .Y(n8555) );
  CLKINVX3 U2707 ( .A(n8553), .Y(n8552) );
  CLKINVX3 U2708 ( .A(n8550), .Y(n8549) );
  CLKINVX3 U2709 ( .A(n8547), .Y(n8546) );
  CLKINVX3 U2710 ( .A(n8544), .Y(n8543) );
  CLKINVX3 U2711 ( .A(n8541), .Y(n8540) );
  CLKINVX3 U2712 ( .A(n8538), .Y(n8537) );
  CLKINVX3 U2713 ( .A(n8535), .Y(n8534) );
  CLKINVX3 U2714 ( .A(n8520), .Y(n8519) );
  CLKINVX3 U2715 ( .A(n8517), .Y(n8516) );
  CLKINVX3 U2716 ( .A(n8514), .Y(n8513) );
  CLKINVX3 U2717 ( .A(n8511), .Y(n8510) );
  CLKINVX3 U2718 ( .A(n8508), .Y(n8507) );
  CLKINVX3 U2719 ( .A(n8505), .Y(n8504) );
  CLKINVX3 U2720 ( .A(n8502), .Y(n8501) );
  CLKINVX3 U2721 ( .A(n8499), .Y(n8498) );
  CLKINVX3 U2722 ( .A(n8496), .Y(n8495) );
  CLKINVX3 U2723 ( .A(n8493), .Y(n8492) );
  CLKINVX3 U2724 ( .A(n8490), .Y(n8489) );
  CLKINVX3 U2725 ( .A(n8487), .Y(n8486) );
  CLKINVX3 U2726 ( .A(n8484), .Y(n8483) );
  CLKINVX3 U2727 ( .A(n8481), .Y(n8480) );
  CLKINVX3 U2728 ( .A(n8478), .Y(n8477) );
  CLKINVX3 U2729 ( .A(n8475), .Y(n8474) );
  CLKINVX3 U2730 ( .A(n8472), .Y(n8471) );
  CLKINVX3 U2731 ( .A(n8469), .Y(n8468) );
  CLKINVX3 U2732 ( .A(n8466), .Y(n8465) );
  CLKINVX3 U2733 ( .A(n8463), .Y(n8462) );
  CLKINVX3 U2734 ( .A(n8460), .Y(n8459) );
  CLKINVX3 U2735 ( .A(n8457), .Y(n8456) );
  CLKINVX3 U2736 ( .A(n8454), .Y(n8453) );
  CLKINVX3 U2737 ( .A(n8451), .Y(n8450) );
  CLKINVX3 U2738 ( .A(n8634), .Y(n8632) );
  INVX1 U2739 ( .A(n1272), .Y(n8634) );
  CLKINVX3 U2740 ( .A(n8640), .Y(n8639) );
  CLKINVX3 U2741 ( .A(n8613), .Y(n8612) );
  CLKINVX3 U2742 ( .A(n8610), .Y(n8609) );
  CLKINVX3 U2743 ( .A(n8601), .Y(n8600) );
  CLKINVX3 U2744 ( .A(n8598), .Y(n8597) );
  CLKINVX3 U2745 ( .A(n8595), .Y(n8594) );
  CLKINVX3 U2746 ( .A(n8592), .Y(n8591) );
  CLKINVX3 U2747 ( .A(n8586), .Y(n8585) );
  CLKINVX3 U2748 ( .A(n8562), .Y(n8561) );
  AND2X2 U2749 ( .A(n8623), .B(n1272), .Y(n1014) );
  AND2X2 U2750 ( .A(n8620), .B(n1272), .Y(n1015) );
  AND2X2 U2751 ( .A(n8617), .B(n1272), .Y(n1016) );
  AND2X2 U2752 ( .A(n8614), .B(n1272), .Y(n1017) );
  AND2X2 U2753 ( .A(n1437), .B(n8623), .Y(n1018) );
  AND2X2 U2754 ( .A(n1437), .B(n8620), .Y(n1019) );
  AND2X2 U2755 ( .A(n1437), .B(n8617), .Y(n1020) );
  AND2X2 U2756 ( .A(n1437), .B(n8614), .Y(n1021) );
  AND2X2 U2757 ( .A(n1471), .B(n8623), .Y(n1022) );
  AND2X2 U2758 ( .A(n1471), .B(n8620), .Y(n1023) );
  AND2X2 U2759 ( .A(n1471), .B(n8617), .Y(n1024) );
  AND2X2 U2760 ( .A(n1471), .B(n8614), .Y(n1025) );
  AND2X2 U2761 ( .A(n1505), .B(n8623), .Y(n1026) );
  AND2X2 U2762 ( .A(n1505), .B(n8620), .Y(n1027) );
  AND2X2 U2763 ( .A(n1505), .B(n8617), .Y(n1028) );
  AND2X2 U2764 ( .A(n1505), .B(n8614), .Y(n1029) );
  AND2X2 U2765 ( .A(n1539), .B(n8623), .Y(n1030) );
  AND2X2 U2766 ( .A(n1539), .B(n8620), .Y(n1031) );
  AND2X2 U2767 ( .A(n1539), .B(n8617), .Y(n1032) );
  AND2X2 U2768 ( .A(n1539), .B(n8614), .Y(n1033) );
  CLKINVX3 U2769 ( .A(n8625), .Y(n8624) );
  CLKINVX3 U2770 ( .A(n8622), .Y(n8621) );
  CLKINVX3 U2771 ( .A(n8619), .Y(n8618) );
  CLKINVX3 U2772 ( .A(n8616), .Y(n8615) );
  CLKINVX3 U2773 ( .A(n8532), .Y(n8531) );
  CLKINVX3 U2774 ( .A(n8529), .Y(n8528) );
  CLKINVX3 U2775 ( .A(n8526), .Y(n8525) );
  CLKINVX3 U2776 ( .A(n8523), .Y(n8522) );
  CLKINVX3 U2777 ( .A(n8640), .Y(n8638) );
  BUFX4 U2778 ( .A(n8760), .Y(n8193) );
  BUFX4 U2779 ( .A(n8760), .Y(n8192) );
  BUFX4 U2780 ( .A(n8760), .Y(n8191) );
  BUFX4 U2781 ( .A(n8761), .Y(n8196) );
  BUFX4 U2782 ( .A(n8761), .Y(n8195) );
  BUFX4 U2783 ( .A(n8761), .Y(n8194) );
  BUFX4 U2784 ( .A(n8762), .Y(n8199) );
  BUFX4 U2785 ( .A(n8762), .Y(n8198) );
  BUFX4 U2786 ( .A(n8762), .Y(n8197) );
  BUFX4 U2787 ( .A(n8763), .Y(n8201) );
  BUFX4 U2788 ( .A(n8763), .Y(n8200) );
  BUFX4 U2789 ( .A(n8763), .Y(n8202) );
  INVX1 U2790 ( .A(n8793), .Y(n8782) );
  INVX1 U2791 ( .A(n8822), .Y(n8811) );
  INVX1 U2792 ( .A(n8851), .Y(n8840) );
  INVX1 U2793 ( .A(n8880), .Y(n8869) );
  INVX1 U2794 ( .A(n8684), .Y(n8674) );
  INVX1 U2795 ( .A(n8714), .Y(n8706) );
  INVX1 U2796 ( .A(n8742), .Y(n8734) );
  INVX1 U2797 ( .A(n8793), .Y(n8783) );
  INVX1 U2798 ( .A(n8822), .Y(n8812) );
  INVX1 U2799 ( .A(n8851), .Y(n8841) );
  INVX1 U2800 ( .A(n8880), .Y(n8870) );
  INVX1 U2801 ( .A(n8684), .Y(n8675) );
  INVX1 U2802 ( .A(n8714), .Y(n8707) );
  INVX1 U2803 ( .A(n8742), .Y(n8735) );
  INVX1 U2804 ( .A(n8792), .Y(n8780) );
  INVX1 U2805 ( .A(n8821), .Y(n8809) );
  INVX1 U2806 ( .A(n8850), .Y(n8838) );
  INVX1 U2807 ( .A(n8879), .Y(n8867) );
  INVX1 U2808 ( .A(n8683), .Y(n8672) );
  INVX1 U2809 ( .A(n8713), .Y(n8704) );
  INVX1 U2810 ( .A(n8741), .Y(n8732) );
  INVX1 U2811 ( .A(n8766), .Y(n8758) );
  INVX1 U2812 ( .A(n8683), .Y(n8673) );
  INVX1 U2813 ( .A(n8713), .Y(n8705) );
  INVX1 U2814 ( .A(n8741), .Y(n8733) );
  INVX1 U2815 ( .A(n8766), .Y(n8759) );
  INVX1 U2816 ( .A(n8792), .Y(n8781) );
  INVX1 U2817 ( .A(n8821), .Y(n8810) );
  INVX1 U2818 ( .A(n8850), .Y(n8839) );
  INVX1 U2819 ( .A(n8879), .Y(n8868) );
  INVX1 U2820 ( .A(n8686), .Y(n8679) );
  INVX1 U2821 ( .A(n8714), .Y(n8710) );
  INVX1 U2822 ( .A(n8742), .Y(n8738) );
  INVX1 U2823 ( .A(n8794), .Y(n8788) );
  INVX1 U2824 ( .A(n8823), .Y(n8817) );
  INVX1 U2825 ( .A(n8852), .Y(n8846) );
  INVX1 U2826 ( .A(n8881), .Y(n8875) );
  INVX1 U2827 ( .A(n8685), .Y(n8680) );
  INVX1 U2828 ( .A(n8794), .Y(n8784) );
  INVX1 U2829 ( .A(n8823), .Y(n8813) );
  INVX1 U2830 ( .A(n8852), .Y(n8842) );
  INVX1 U2831 ( .A(n8881), .Y(n8871) );
  INVX1 U2832 ( .A(n8685), .Y(n8676) );
  INVX1 U2833 ( .A(n8715), .Y(n8708) );
  INVX1 U2834 ( .A(n8743), .Y(n8736) );
  INVX1 U2835 ( .A(n8794), .Y(n8785) );
  INVX1 U2836 ( .A(n8823), .Y(n8814) );
  INVX1 U2837 ( .A(n8852), .Y(n8843) );
  INVX1 U2838 ( .A(n8881), .Y(n8872) );
  INVX1 U2839 ( .A(n8685), .Y(n8677) );
  INVX1 U2840 ( .A(n8715), .Y(n8709) );
  INVX1 U2841 ( .A(n8743), .Y(n8737) );
  INVX1 U2842 ( .A(n8795), .Y(n8786) );
  INVX1 U2843 ( .A(n8824), .Y(n8815) );
  INVX1 U2844 ( .A(n8853), .Y(n8844) );
  INVX1 U2845 ( .A(n8882), .Y(n8873) );
  INVX1 U2846 ( .A(n8686), .Y(n8678) );
  INVX1 U2847 ( .A(n8795), .Y(n8787) );
  INVX1 U2848 ( .A(n8824), .Y(n8816) );
  INVX1 U2849 ( .A(n8853), .Y(n8845) );
  INVX1 U2850 ( .A(n8882), .Y(n8874) );
  INVX1 U2851 ( .A(n8712), .Y(n8696) );
  INVX1 U2852 ( .A(n8740), .Y(n8724) );
  INVX1 U2853 ( .A(n8767), .Y(n8752) );
  INVX1 U2854 ( .A(n8794), .Y(n8774) );
  INVX1 U2855 ( .A(n8823), .Y(n8803) );
  INVX1 U2856 ( .A(n8852), .Y(n8832) );
  INVX1 U2857 ( .A(n8881), .Y(n8861) );
  INVX1 U2858 ( .A(n8712), .Y(n8697) );
  INVX1 U2859 ( .A(n8740), .Y(n8725) );
  INVX1 U2860 ( .A(n8765), .Y(n8751) );
  INVX1 U2861 ( .A(n8712), .Y(n8695) );
  INVX1 U2862 ( .A(n8740), .Y(n8723) );
  INVX1 U2863 ( .A(n8684), .Y(n8669) );
  INVX1 U2864 ( .A(n8712), .Y(n8701) );
  INVX1 U2865 ( .A(n8740), .Y(n8729) );
  INVX1 U2866 ( .A(n8791), .Y(n8778) );
  INVX1 U2867 ( .A(n8820), .Y(n8807) );
  INVX1 U2868 ( .A(n8849), .Y(n8836) );
  INVX1 U2869 ( .A(n8878), .Y(n8865) );
  INVX1 U2870 ( .A(n8766), .Y(n8756) );
  INVX1 U2871 ( .A(n8682), .Y(n8670) );
  INVX1 U2872 ( .A(n8714), .Y(n8702) );
  INVX1 U2873 ( .A(n8742), .Y(n8730) );
  INVX1 U2874 ( .A(n8790), .Y(n8775) );
  INVX1 U2875 ( .A(n8819), .Y(n8804) );
  INVX1 U2876 ( .A(n8848), .Y(n8833) );
  INVX1 U2877 ( .A(n8877), .Y(n8862) );
  INVX1 U2878 ( .A(n8683), .Y(n8666) );
  INVX1 U2879 ( .A(n8714), .Y(n8698) );
  INVX1 U2880 ( .A(n8742), .Y(n8726) );
  INVX1 U2881 ( .A(n8765), .Y(n8753) );
  INVX1 U2882 ( .A(n8790), .Y(n8776) );
  INVX1 U2883 ( .A(n8819), .Y(n8805) );
  INVX1 U2884 ( .A(n8848), .Y(n8834) );
  INVX1 U2885 ( .A(n8877), .Y(n8863) );
  INVX1 U2886 ( .A(n8682), .Y(n8667) );
  INVX1 U2887 ( .A(n8713), .Y(n8699) );
  INVX1 U2888 ( .A(n8741), .Y(n8727) );
  INVX1 U2889 ( .A(n8766), .Y(n8754) );
  INVX1 U2890 ( .A(n8686), .Y(n8668) );
  INVX1 U2891 ( .A(n8712), .Y(n8700) );
  INVX1 U2892 ( .A(n8740), .Y(n8728) );
  INVX1 U2893 ( .A(n8766), .Y(n8755) );
  INVX1 U2894 ( .A(n8790), .Y(n8777) );
  INVX1 U2895 ( .A(n8819), .Y(n8806) );
  INVX1 U2896 ( .A(n8848), .Y(n8835) );
  INVX1 U2897 ( .A(n8877), .Y(n8864) );
  INVX1 U2898 ( .A(n8682), .Y(n8671) );
  INVX1 U2899 ( .A(n8713), .Y(n8703) );
  INVX1 U2900 ( .A(n8741), .Y(n8731) );
  INVX1 U2901 ( .A(n8767), .Y(n8757) );
  INVX1 U2902 ( .A(n8791), .Y(n8779) );
  INVX1 U2903 ( .A(n8820), .Y(n8808) );
  INVX1 U2904 ( .A(n8849), .Y(n8837) );
  INVX1 U2905 ( .A(n8878), .Y(n8866) );
  INVX1 U2906 ( .A(n8690), .Y(n8681) );
  INVX1 U2907 ( .A(n8717), .Y(n8711) );
  INVX1 U2908 ( .A(n8745), .Y(n8739) );
  INVX1 U2909 ( .A(n8769), .Y(n8764) );
  INVX1 U2910 ( .A(n8798), .Y(n8789) );
  INVX1 U2911 ( .A(n8827), .Y(n8818) );
  INVX1 U2912 ( .A(n8856), .Y(n8847) );
  INVX1 U2913 ( .A(n8885), .Y(n8876) );
  CLKINVX3 U2914 ( .A(n7989), .Y(n7991) );
  INVX1 U2915 ( .A(n7619), .Y(n7370) );
  INVX1 U2916 ( .A(n4025), .Y(n4026) );
  INVX1 U2917 ( .A(n4275), .Y(n4276) );
  INVX1 U2918 ( .A(n4275), .Y(n4277) );
  INVX1 U2919 ( .A(n4278), .Y(n4279) );
  INVX1 U2920 ( .A(N84), .Y(n7989) );
  CLKINVX3 U2921 ( .A(n8652), .Y(n4646) );
  INVX1 U2922 ( .A(n7979), .Y(n7980) );
  INVX1 U2923 ( .A(n4625), .Y(n4626) );
  INVX1 U2924 ( .A(n8657), .Y(n4560) );
  INVX1 U2925 ( .A(n8646), .Y(n7969) );
  INVX1 U2926 ( .A(n8647), .Y(n7903) );
  INVX1 U2927 ( .A(n8646), .Y(n7968) );
  INVX1 U2928 ( .A(n8645), .Y(n7978) );
  AND2X2 U2929 ( .A(n8639), .B(n1269), .Y(n1267) );
  AND2X2 U2930 ( .A(ena_in), .B(n1269), .Y(n1272) );
  CLKINVX3 U2931 ( .A(n8637), .Y(n8635) );
  INVX1 U2932 ( .A(n1271), .Y(n8637) );
  CLKINVX3 U2933 ( .A(n8631), .Y(n8629) );
  INVX1 U2934 ( .A(n1274), .Y(n8631) );
  CLKINVX3 U2935 ( .A(n8628), .Y(n8626) );
  INVX1 U2936 ( .A(n1276), .Y(n8628) );
  CLKINVX3 U2937 ( .A(n8607), .Y(n8605) );
  INVX1 U2938 ( .A(n1290), .Y(n8607) );
  CLKINVX3 U2939 ( .A(n8604), .Y(n8602) );
  INVX1 U2940 ( .A(n1292), .Y(n8604) );
  CLKINVX3 U2941 ( .A(n8589), .Y(n8587) );
  INVX1 U2942 ( .A(n1302), .Y(n8589) );
  CLKINVX3 U2943 ( .A(n8583), .Y(n8581) );
  INVX1 U2944 ( .A(n1306), .Y(n8583) );
  CLKINVX3 U2945 ( .A(n8580), .Y(n8578) );
  INVX1 U2946 ( .A(n1308), .Y(n8580) );
  CLKINVX3 U2947 ( .A(n8577), .Y(n8575) );
  INVX1 U2948 ( .A(n1310), .Y(n8577) );
  CLKINVX3 U2949 ( .A(n8574), .Y(n8572) );
  INVX1 U2950 ( .A(n1312), .Y(n8574) );
  CLKINVX3 U2951 ( .A(n8571), .Y(n8569) );
  INVX1 U2952 ( .A(n1314), .Y(n8571) );
  CLKINVX3 U2953 ( .A(n8568), .Y(n8566) );
  INVX1 U2954 ( .A(n1316), .Y(n8568) );
  CLKINVX3 U2955 ( .A(n8565), .Y(n8563) );
  INVX1 U2956 ( .A(n1318), .Y(n8565) );
  CLKINVX3 U2957 ( .A(n8559), .Y(n8557) );
  INVX1 U2958 ( .A(n1322), .Y(n8559) );
  CLKINVX3 U2959 ( .A(n8556), .Y(n8554) );
  INVX1 U2960 ( .A(n1324), .Y(n8556) );
  CLKINVX3 U2961 ( .A(n8553), .Y(n8551) );
  INVX1 U2962 ( .A(n1326), .Y(n8553) );
  CLKINVX3 U2963 ( .A(n8550), .Y(n8548) );
  INVX1 U2964 ( .A(n1328), .Y(n8550) );
  CLKINVX3 U2965 ( .A(n8547), .Y(n8545) );
  INVX1 U2966 ( .A(n1330), .Y(n8547) );
  CLKINVX3 U2967 ( .A(n8544), .Y(n8542) );
  INVX1 U2968 ( .A(n1332), .Y(n8544) );
  CLKINVX3 U2969 ( .A(n8541), .Y(n8539) );
  INVX1 U2970 ( .A(n1334), .Y(n8541) );
  CLKINVX3 U2971 ( .A(n8538), .Y(n8536) );
  INVX1 U2972 ( .A(n1369), .Y(n8538) );
  CLKINVX3 U2973 ( .A(n8535), .Y(n8533) );
  INVX1 U2974 ( .A(n1403), .Y(n8535) );
  CLKINVX3 U2975 ( .A(n8520), .Y(n8518) );
  INVX1 U2976 ( .A(n1573), .Y(n8520) );
  CLKINVX3 U2977 ( .A(n8517), .Y(n8515) );
  INVX1 U2978 ( .A(n1608), .Y(n8517) );
  CLKINVX3 U2979 ( .A(n8514), .Y(n8512) );
  INVX1 U2980 ( .A(n1641), .Y(n8514) );
  CLKINVX3 U2981 ( .A(n8511), .Y(n8509) );
  INVX1 U2982 ( .A(n1674), .Y(n8511) );
  CLKINVX3 U2983 ( .A(n8508), .Y(n8506) );
  INVX1 U2984 ( .A(n1707), .Y(n8508) );
  CLKINVX3 U2985 ( .A(n8505), .Y(n8503) );
  INVX1 U2986 ( .A(n1740), .Y(n8505) );
  CLKINVX3 U2987 ( .A(n8502), .Y(n8500) );
  INVX1 U2988 ( .A(n1773), .Y(n8502) );
  CLKINVX3 U2989 ( .A(n8499), .Y(n8497) );
  INVX1 U2990 ( .A(n1806), .Y(n8499) );
  CLKINVX3 U2991 ( .A(n8496), .Y(n8494) );
  INVX1 U2992 ( .A(n1839), .Y(n8496) );
  CLKINVX3 U2993 ( .A(n8493), .Y(n8491) );
  INVX1 U2994 ( .A(n1873), .Y(n8493) );
  CLKINVX3 U2995 ( .A(n8490), .Y(n8488) );
  INVX1 U2996 ( .A(n1906), .Y(n8490) );
  CLKINVX3 U2997 ( .A(n8487), .Y(n8485) );
  INVX1 U2998 ( .A(n1939), .Y(n8487) );
  CLKINVX3 U2999 ( .A(n8484), .Y(n8482) );
  INVX1 U3000 ( .A(n1972), .Y(n8484) );
  CLKINVX3 U3001 ( .A(n8481), .Y(n8479) );
  INVX1 U3002 ( .A(n2005), .Y(n8481) );
  CLKINVX3 U3003 ( .A(n8478), .Y(n8476) );
  INVX1 U3004 ( .A(n2038), .Y(n8478) );
  CLKINVX3 U3005 ( .A(n8475), .Y(n8473) );
  INVX1 U3006 ( .A(n2071), .Y(n8475) );
  CLKINVX3 U3007 ( .A(n8472), .Y(n8470) );
  INVX1 U3008 ( .A(n2104), .Y(n8472) );
  CLKINVX3 U3009 ( .A(n8469), .Y(n8467) );
  INVX1 U3010 ( .A(n2138), .Y(n8469) );
  CLKINVX3 U3011 ( .A(n8466), .Y(n8464) );
  INVX1 U3012 ( .A(n2171), .Y(n8466) );
  CLKINVX3 U3013 ( .A(n8463), .Y(n8461) );
  INVX1 U3014 ( .A(n2204), .Y(n8463) );
  CLKINVX3 U3015 ( .A(n8460), .Y(n8458) );
  INVX1 U3016 ( .A(n2237), .Y(n8460) );
  CLKINVX3 U3017 ( .A(n8457), .Y(n8455) );
  INVX1 U3018 ( .A(n2270), .Y(n8457) );
  CLKINVX3 U3019 ( .A(n8454), .Y(n8452) );
  INVX1 U3020 ( .A(n2303), .Y(n8454) );
  CLKINVX3 U3021 ( .A(n8451), .Y(n8449) );
  INVX1 U3022 ( .A(n2336), .Y(n8451) );
  INVX1 U3023 ( .A(n1286), .Y(n8613) );
  INVX1 U3024 ( .A(n1288), .Y(n8610) );
  INVX1 U3025 ( .A(n1294), .Y(n8601) );
  INVX1 U3026 ( .A(n1296), .Y(n8598) );
  INVX1 U3027 ( .A(n1298), .Y(n8595) );
  INVX1 U3028 ( .A(n1300), .Y(n8592) );
  INVX1 U3029 ( .A(n1304), .Y(n8586) );
  INVX1 U3030 ( .A(n1320), .Y(n8562) );
  INVX1 U3031 ( .A(n1268), .Y(n8640) );
  CLKINVX3 U3032 ( .A(n8622), .Y(n8620) );
  INVX1 U3033 ( .A(n1280), .Y(n8622) );
  CLKINVX3 U3034 ( .A(n8616), .Y(n8614) );
  INVX1 U3035 ( .A(n1284), .Y(n8616) );
  CLKINVX3 U3036 ( .A(n8532), .Y(n8530) );
  INVX1 U3037 ( .A(n1437), .Y(n8532) );
  CLKINVX3 U3038 ( .A(n8529), .Y(n8527) );
  INVX1 U3039 ( .A(n1471), .Y(n8529) );
  CLKINVX3 U3040 ( .A(n8526), .Y(n8524) );
  INVX1 U3041 ( .A(n1505), .Y(n8526) );
  CLKINVX3 U3042 ( .A(n8523), .Y(n8521) );
  INVX1 U3043 ( .A(n1539), .Y(n8523) );
  BUFX3 U3044 ( .A(n8959), .Y(n8436) );
  BUFX3 U3045 ( .A(n1034), .Y(n8438) );
  BUFX3 U3046 ( .A(n1035), .Y(n8437) );
  CLKINVX3 U3047 ( .A(n8625), .Y(n8623) );
  INVX1 U3048 ( .A(n1278), .Y(n8625) );
  CLKINVX3 U3049 ( .A(n8619), .Y(n8617) );
  INVX1 U3050 ( .A(n1282), .Y(n8619) );
  INVX1 U3051 ( .A(n1240), .Y(n8958) );
  BUFX3 U3052 ( .A(n8959), .Y(n8435) );
  INVX1 U3053 ( .A(n8767), .Y(n8760) );
  INVX1 U3054 ( .A(n8767), .Y(n8761) );
  INVX1 U3055 ( .A(n8767), .Y(n8762) );
  INVX1 U3056 ( .A(n8765), .Y(n8763) );
  INVX1 U3057 ( .A(n8797), .Y(n8793) );
  INVX1 U3058 ( .A(n8826), .Y(n8822) );
  INVX1 U3059 ( .A(n8855), .Y(n8851) );
  INVX1 U3060 ( .A(n8884), .Y(n8880) );
  INVX1 U3061 ( .A(n8688), .Y(n8684) );
  INVX1 U3062 ( .A(n8708), .Y(n8714) );
  INVX1 U3063 ( .A(n8736), .Y(n8742) );
  INVX1 U3064 ( .A(n8688), .Y(n8683) );
  INVX1 U3065 ( .A(n8709), .Y(n8713) );
  INVX1 U3066 ( .A(n8737), .Y(n8741) );
  INVX1 U3067 ( .A(n8751), .Y(n8766) );
  INVX1 U3068 ( .A(n8797), .Y(n8792) );
  INVX1 U3069 ( .A(n8826), .Y(n8821) );
  INVX1 U3070 ( .A(n8855), .Y(n8850) );
  INVX1 U3071 ( .A(n8884), .Y(n8879) );
  INVX1 U3072 ( .A(n8796), .Y(n8794) );
  INVX1 U3073 ( .A(n8825), .Y(n8823) );
  INVX1 U3074 ( .A(n8854), .Y(n8852) );
  INVX1 U3075 ( .A(n8883), .Y(n8881) );
  INVX1 U3076 ( .A(n8687), .Y(n8685) );
  INVX1 U3077 ( .A(n8716), .Y(n8715) );
  INVX1 U3078 ( .A(n8744), .Y(n8743) );
  INVX1 U3079 ( .A(n8687), .Y(n8686) );
  INVX1 U3080 ( .A(n8796), .Y(n8795) );
  INVX1 U3081 ( .A(n8825), .Y(n8824) );
  INVX1 U3082 ( .A(n8854), .Y(n8853) );
  INVX1 U3083 ( .A(n8883), .Y(n8882) );
  INVX1 U3084 ( .A(n8716), .Y(n8712) );
  INVX1 U3085 ( .A(n8744), .Y(n8740) );
  INVX1 U3086 ( .A(n8769), .Y(n8765) );
  INVX1 U3087 ( .A(n8797), .Y(n8790) );
  INVX1 U3088 ( .A(n8826), .Y(n8819) );
  INVX1 U3089 ( .A(n8855), .Y(n8848) );
  INVX1 U3090 ( .A(n8884), .Y(n8877) );
  INVX1 U3091 ( .A(n8688), .Y(n8682) );
  INVX1 U3092 ( .A(n8797), .Y(n8791) );
  INVX1 U3093 ( .A(n8826), .Y(n8820) );
  INVX1 U3094 ( .A(n8855), .Y(n8849) );
  INVX1 U3095 ( .A(n8884), .Y(n8878) );
  INVX1 U3096 ( .A(n8691), .Y(n8690) );
  INVX1 U3097 ( .A(n8718), .Y(n8717) );
  INVX1 U3098 ( .A(n8746), .Y(n8745) );
  INVX1 U3099 ( .A(n8770), .Y(n8769) );
  INVX1 U3100 ( .A(n8799), .Y(n8798) );
  INVX1 U3101 ( .A(n8828), .Y(n8827) );
  INVX1 U3102 ( .A(n8857), .Y(n8856) );
  INVX1 U3103 ( .A(n8886), .Y(n8885) );
  MX4X1 U3104 ( .A(n1548), .B(n1365), .C(n1457), .D(n1171), .S0(N77), .S1(N76), 
        .Y(N1234) );
  MX4X1 U3105 ( .A(n1364), .B(n1309), .C(n1343), .D(n1209), .S0(n4648), .S1(
        n4647), .Y(n1365) );
  MX4X1 U3106 ( .A(n1170), .B(n1086), .C(n1107), .D(n1065), .S0(n4648), .S1(
        n4646), .Y(n1171) );
  MX4X1 U3107 ( .A(n1547), .B(n1501), .C(n1524), .D(n1480), .S0(n4648), .S1(
        n8651), .Y(n1548) );
  MX4X1 U3108 ( .A(n1902), .B(n1726), .C(n1814), .D(n1638), .S0(N77), .S1(N76), 
        .Y(N1233) );
  MX4X1 U3109 ( .A(n1725), .B(n1682), .C(n1703), .D(n1660), .S0(n4648), .S1(
        N74), .Y(n1726) );
  MX4X1 U3110 ( .A(n1637), .B(n1592), .C(n1616), .D(n1569), .S0(n4648), .S1(
        N74), .Y(n1638) );
  MX4X1 U3111 ( .A(n1901), .B(n1857), .C(n1880), .D(n1835), .S0(n4648), .S1(
        N74), .Y(n1902) );
  MX4X1 U3112 ( .A(n2254), .B(n2078), .C(n2166), .D(n1990), .S0(N77), .S1(N76), 
        .Y(N1232) );
  MX4X1 U3113 ( .A(n2077), .B(n2033), .C(n2055), .D(n2012), .S0(n4649), .S1(
        n8651), .Y(n2078) );
  MX4X1 U3114 ( .A(n1989), .B(n1946), .C(n1967), .D(n1924), .S0(n4649), .S1(
        n4646), .Y(n1990) );
  MX4X1 U3115 ( .A(n2253), .B(n2210), .C(n2231), .D(n2188), .S0(n4649), .S1(
        N74), .Y(n2254) );
  MX4X1 U3116 ( .A(n2664), .B(n2494), .C(n2579), .D(n2349), .S0(N77), .S1(N76), 
        .Y(N1231) );
  MX4X1 U3117 ( .A(n2493), .B(n2451), .C(n2472), .D(n2375), .S0(n4649), .S1(
        n8651), .Y(n2494) );
  MX4X1 U3118 ( .A(n2347), .B(n2297), .C(n2319), .D(n2276), .S0(n4649), .S1(
        n8651), .Y(n2349) );
  MX4X1 U3119 ( .A(n2663), .B(n2621), .C(n2642), .D(n2600), .S0(n4649), .S1(
        N74), .Y(n2664) );
  MX4X1 U3120 ( .A(n3004), .B(n2834), .C(n2919), .D(n2749), .S0(N77), .S1(N76), 
        .Y(N1230) );
  MX4X1 U3121 ( .A(n2833), .B(n2791), .C(n2812), .D(n2770), .S0(n4649), .S1(
        n4647), .Y(n2834) );
  MX4X1 U3122 ( .A(n2748), .B(n2706), .C(n2727), .D(n2685), .S0(n4649), .S1(
        N74), .Y(n2749) );
  MX4X1 U3123 ( .A(n3003), .B(n2961), .C(n2982), .D(n2940), .S0(n4649), .S1(
        n4646), .Y(n3004) );
  MX4X1 U3124 ( .A(n3344), .B(n3174), .C(n3259), .D(n3089), .S0(N77), .S1(N76), 
        .Y(N1229) );
  MX4X1 U3125 ( .A(n3173), .B(n3131), .C(n3152), .D(n3110), .S0(n4648), .S1(
        n4646), .Y(n3174) );
  MX4X1 U3126 ( .A(n3088), .B(n3046), .C(n3067), .D(n3025), .S0(n4648), .S1(
        n4646), .Y(n3089) );
  MX4X1 U3127 ( .A(n3343), .B(n3301), .C(n3322), .D(n3280), .S0(N75), .S1(
        n4646), .Y(n3344) );
  MX4X1 U3128 ( .A(n3684), .B(n3514), .C(n3599), .D(n3429), .S0(N77), .S1(N76), 
        .Y(N1228) );
  MX4X1 U3129 ( .A(n3513), .B(n3471), .C(n3492), .D(n3450), .S0(N75), .S1(
        n4646), .Y(n3514) );
  MX4X1 U3130 ( .A(n3428), .B(n3386), .C(n3407), .D(n3365), .S0(n4648), .S1(
        n4646), .Y(n3429) );
  MX4X1 U3131 ( .A(n3683), .B(n3641), .C(n3662), .D(n3620), .S0(N75), .S1(
        n4646), .Y(n3684) );
  MX4X1 U3132 ( .A(n4024), .B(n3854), .C(n3939), .D(n3769), .S0(N77), .S1(N76), 
        .Y(N1227) );
  MX4X1 U3133 ( .A(n3853), .B(n3811), .C(n3832), .D(n3790), .S0(N75), .S1(
        n4646), .Y(n3854) );
  MX4X1 U3134 ( .A(n3768), .B(n3726), .C(n3747), .D(n3705), .S0(n4648), .S1(
        n4646), .Y(n3769) );
  MX4X1 U3135 ( .A(n4023), .B(n3981), .C(n4002), .D(n3960), .S0(N75), .S1(
        n4646), .Y(n4024) );
  INVX1 U3136 ( .A(n1259), .Y(n8923) );
  INVX1 U3137 ( .A(N85), .Y(n8641) );
  INVX1 U3138 ( .A(N68), .Y(n4025) );
  INVX1 U3139 ( .A(n4502), .Y(n4278) );
  INVX1 U3140 ( .A(n4503), .Y(n4275) );
  INVX1 U3141 ( .A(n7618), .Y(n7619) );
  INVX1 U3142 ( .A(n8648), .Y(n7618) );
  INVX1 U3143 ( .A(n8649), .Y(n8648) );
  INVX1 U3144 ( .A(N78), .Y(n8649) );
  INVX1 U3145 ( .A(N75), .Y(n8650) );
  INVX1 U3146 ( .A(N73), .Y(n8653) );
  INVX1 U3147 ( .A(n8642), .Y(n7979) );
  INVX1 U3148 ( .A(n8643), .Y(n8642) );
  INVX1 U3149 ( .A(N83), .Y(n8643) );
  INVX1 U3150 ( .A(n8655), .Y(n4625) );
  INVX1 U3151 ( .A(n8656), .Y(n8655) );
  INVX1 U3152 ( .A(N71), .Y(n8656) );
  INVX1 U3153 ( .A(N70), .Y(n8657) );
  INVX1 U3154 ( .A(N81), .Y(n8646) );
  INVX1 U3155 ( .A(N80), .Y(n8647) );
  INVX1 U3156 ( .A(n8645), .Y(n8644) );
  INVX1 U3157 ( .A(N82), .Y(n8645) );
  INVX1 U3158 ( .A(n8652), .Y(n4647) );
  INVX1 U3159 ( .A(n8652), .Y(n8651) );
  INVX1 U3160 ( .A(N74), .Y(n8652) );
  INVX1 U3161 ( .A(N72), .Y(n8654) );
  NAND2X2 U3162 ( .A(n8660), .B(n1267), .Y(n1265) );
  AND2X2 U3163 ( .A(n1605), .B(n1366), .Y(n1269) );
  AND3X2 U3164 ( .A(n8661), .B(n1605), .C(n1606), .Y(n1573) );
  AND3X2 U3165 ( .A(n1367), .B(n8660), .C(n1606), .Y(n1608) );
  AND3X2 U3166 ( .A(n1401), .B(n8660), .C(n1606), .Y(n1641) );
  AND3X2 U3167 ( .A(n1435), .B(n8660), .C(n1606), .Y(n1674) );
  AND3X2 U3168 ( .A(n1469), .B(n8660), .C(n1606), .Y(n1707) );
  AND3X2 U3169 ( .A(n1503), .B(n8660), .C(n1606), .Y(n1740) );
  AND3X2 U3170 ( .A(n1537), .B(n8660), .C(n1606), .Y(n1773) );
  AND3X2 U3171 ( .A(n1571), .B(n8660), .C(n1606), .Y(n1806) );
  AND3X2 U3172 ( .A(n8661), .B(n1605), .C(n1871), .Y(n1839) );
  AND3X2 U3173 ( .A(n1367), .B(n8660), .C(n1871), .Y(n1873) );
  AND3X2 U3174 ( .A(n1401), .B(n8660), .C(n1871), .Y(n1906) );
  AND3X2 U3175 ( .A(n1435), .B(n8661), .C(n1871), .Y(n1939) );
  AND3X2 U3176 ( .A(n1469), .B(n8661), .C(n1871), .Y(n1972) );
  AND3X2 U3177 ( .A(n1503), .B(n8661), .C(n1871), .Y(n2005) );
  AND3X2 U3178 ( .A(n1537), .B(n8661), .C(n1871), .Y(n2038) );
  AND3X2 U3179 ( .A(n1571), .B(n8661), .C(n1871), .Y(n2071) );
  AND3X2 U3180 ( .A(n8661), .B(n1605), .C(n2136), .Y(n2104) );
  AND3X2 U3181 ( .A(n1367), .B(n8661), .C(n2136), .Y(n2138) );
  AND3X2 U3182 ( .A(n1401), .B(n8661), .C(n2136), .Y(n2171) );
  AND3X2 U3183 ( .A(n1435), .B(n8661), .C(n2136), .Y(n2204) );
  AND3X2 U3184 ( .A(n1469), .B(n8661), .C(n2136), .Y(n2237) );
  AND3X2 U3185 ( .A(n1503), .B(n8661), .C(n2136), .Y(n2270) );
  AND3X2 U3186 ( .A(n1537), .B(n8661), .C(n2136), .Y(n2303) );
  AND3X2 U3187 ( .A(n1571), .B(n8660), .C(n2136), .Y(n2336) );
  AND3X2 U3188 ( .A(n8660), .B(n1366), .C(n1367), .Y(n1334) );
  AND3X2 U3189 ( .A(ena_in), .B(n1366), .C(n1401), .Y(n1369) );
  AND3X2 U3190 ( .A(ena_in), .B(n1366), .C(n1435), .Y(n1403) );
  AND2X2 U3191 ( .A(n2354), .B(n2342), .Y(n1290) );
  AND2X2 U3192 ( .A(n2363), .B(n2342), .Y(n1306) );
  AND2X2 U3193 ( .A(n2372), .B(n2342), .Y(n1322) );
  AND2X2 U3194 ( .A(n2342), .B(n8439), .Y(n1274) );
  AND2X2 U3195 ( .A(n2354), .B(n2337), .Y(n1286) );
  AND2X2 U3196 ( .A(n2354), .B(n2340), .Y(n1288) );
  AND2X2 U3197 ( .A(n2354), .B(n2344), .Y(n1292) );
  AND2X2 U3198 ( .A(n2354), .B(n2346), .Y(n1294) );
  AND2X2 U3199 ( .A(n2354), .B(n2348), .Y(n1296) );
  AND2X2 U3200 ( .A(n2354), .B(n2350), .Y(n1298) );
  AND2X2 U3201 ( .A(n2354), .B(n2352), .Y(n1300) );
  AND2X2 U3202 ( .A(n2363), .B(n2337), .Y(n1302) );
  AND2X2 U3203 ( .A(n2363), .B(n2340), .Y(n1304) );
  AND2X2 U3204 ( .A(n2363), .B(n2344), .Y(n1308) );
  AND2X2 U3205 ( .A(n2363), .B(n2346), .Y(n1310) );
  AND2X2 U3206 ( .A(n2363), .B(n2348), .Y(n1312) );
  AND2X2 U3207 ( .A(n2363), .B(n2350), .Y(n1314) );
  AND2X2 U3208 ( .A(n2363), .B(n2352), .Y(n1316) );
  AND2X2 U3209 ( .A(n2372), .B(n2337), .Y(n1318) );
  AND2X2 U3210 ( .A(n2372), .B(n2340), .Y(n1320) );
  AND2X2 U3211 ( .A(n2372), .B(n2344), .Y(n1324) );
  AND2X2 U3212 ( .A(n2372), .B(n2346), .Y(n1326) );
  AND2X2 U3213 ( .A(n2372), .B(n2348), .Y(n1328) );
  AND2X2 U3214 ( .A(n2372), .B(n2350), .Y(n1330) );
  AND2X2 U3215 ( .A(n2372), .B(n2352), .Y(n1332) );
  AND2X2 U3216 ( .A(n2337), .B(n8439), .Y(n1268) );
  AND2X2 U3217 ( .A(n2340), .B(n8439), .Y(n1271) );
  AND2X2 U3218 ( .A(n2344), .B(n8439), .Y(n1276) );
  AND2X2 U3219 ( .A(n1269), .B(n8439), .Y(n2381) );
  AND3X2 U3220 ( .A(ena_in), .B(n1366), .C(n1469), .Y(n1437) );
  AND3X2 U3221 ( .A(ena_in), .B(n1366), .C(n1503), .Y(n1471) );
  AND3X2 U3222 ( .A(n8661), .B(n1366), .C(n1537), .Y(n1505) );
  AND3X2 U3223 ( .A(ena_in), .B(n1366), .C(n1571), .Y(n1539) );
  AND2X2 U3224 ( .A(n2346), .B(n8439), .Y(n1278) );
  AND2X2 U3225 ( .A(n2348), .B(n8439), .Y(n1280) );
  AND2X2 U3226 ( .A(n2350), .B(n8439), .Y(n1282) );
  AND2X2 U3227 ( .A(n2352), .B(n8439), .Y(n1284) );
  CLKINVX3 U3228 ( .A(n8662), .Y(n8661) );
  AND3X2 U3229 ( .A(n2342), .B(n8660), .C(n2381), .Y(n1034) );
  AND3X2 U3230 ( .A(n2346), .B(n8660), .C(n2381), .Y(n1035) );
  INVX1 U3231 ( .A(n1261), .Y(n8959) );
  OAI21X1 U3232 ( .A0(n8960), .A1(n8963), .B0(n8973), .Y(n1240) );
  NOR2X1 U3233 ( .A(n8960), .B(n1187), .Y(n1257) );
  NOR2X1 U3234 ( .A(n8963), .B(n1197), .Y(n1194) );
  INVX1 U3235 ( .A(n1187), .Y(n8963) );
  INVX1 U3236 ( .A(n8664), .Y(n8687) );
  INVX1 U3237 ( .A(n8719), .Y(n8716) );
  INVX1 U3238 ( .A(n8747), .Y(n8744) );
  INVX1 U3239 ( .A(n8799), .Y(n8796) );
  INVX1 U3240 ( .A(n8828), .Y(n8825) );
  INVX1 U3241 ( .A(n8857), .Y(n8854) );
  INVX1 U3242 ( .A(n8886), .Y(n8883) );
  INVX1 U3243 ( .A(n8691), .Y(n8689) );
  INVX1 U3244 ( .A(n8691), .Y(n8688) );
  INVX1 U3245 ( .A(n8799), .Y(n8797) );
  INVX1 U3246 ( .A(n8828), .Y(n8826) );
  INVX1 U3247 ( .A(n8857), .Y(n8855) );
  INVX1 U3248 ( .A(n8886), .Y(n8884) );
  INVX1 U3249 ( .A(n8768), .Y(n8767) );
  INVX1 U3250 ( .A(n1197), .Y(n8961) );
  BUFX3 U3251 ( .A(n1185), .Y(n8448) );
  NAND3X1 U3252 ( .A(n8961), .B(n1186), .C(n1187), .Y(n1185) );
  BUFX4 U3253 ( .A(n1218), .Y(n8442) );
  NOR3X1 U3254 ( .A(N1408), .B(rst), .C(n8436), .Y(n1218) );
  INVX1 U3255 ( .A(n8663), .Y(n8691) );
  INVX1 U3256 ( .A(n8692), .Y(n8718) );
  INVX1 U3257 ( .A(n8720), .Y(n8746) );
  INVX1 U3258 ( .A(n8771), .Y(n8799) );
  INVX1 U3259 ( .A(n8800), .Y(n8828) );
  INVX1 U3260 ( .A(n8829), .Y(n8857) );
  INVX1 U3261 ( .A(n8748), .Y(n8770) );
  INVX1 U3262 ( .A(n8858), .Y(n8886) );
  AND3X2 U3263 ( .A(n1200), .B(n8915), .C(n1203), .Y(n1036) );
  AND3X2 U3264 ( .A(n1200), .B(n8915), .C(n1199), .Y(n1037) );
  AND3X2 U3265 ( .A(n1203), .B(n8915), .C(n1206), .Y(n1038) );
  AND3X2 U3266 ( .A(n1199), .B(n8915), .C(n1206), .Y(n1039) );
  MX4X1 U3267 ( .A(n4989), .B(n4819), .C(n4904), .D(n4734), .S0(N87), .S1(N86), 
        .Y(N1315) );
  MX4X1 U3268 ( .A(n4818), .B(n4776), .C(n4797), .D(n4755), .S0(n7992), .S1(
        N84), .Y(n4819) );
  MX4X1 U3269 ( .A(n4733), .B(n4691), .C(n4712), .D(n4670), .S0(n7992), .S1(
        n7991), .Y(n4734) );
  MX4X1 U3270 ( .A(n4988), .B(n4946), .C(n4967), .D(n4925), .S0(n7992), .S1(
        n7990), .Y(n4989) );
  MX4X1 U3271 ( .A(n5329), .B(n5159), .C(n5244), .D(n5074), .S0(N87), .S1(N86), 
        .Y(N1314) );
  MX4X1 U3272 ( .A(n5158), .B(n5116), .C(n5137), .D(n5095), .S0(n7992), .S1(
        N84), .Y(n5159) );
  MX4X1 U3273 ( .A(n5073), .B(n5031), .C(n5052), .D(n5010), .S0(n7992), .S1(
        n7990), .Y(n5074) );
  MX4X1 U3274 ( .A(n5328), .B(n5286), .C(n5307), .D(n5265), .S0(n7992), .S1(
        n7990), .Y(n5329) );
  MX4X1 U3275 ( .A(n5669), .B(n5499), .C(n5584), .D(n5414), .S0(N87), .S1(N86), 
        .Y(N1313) );
  MX4X1 U3276 ( .A(n5498), .B(n5456), .C(n5477), .D(n5435), .S0(n7993), .S1(
        n7990), .Y(n5499) );
  MX4X1 U3277 ( .A(n5413), .B(n5371), .C(n5392), .D(n5350), .S0(n7993), .S1(
        n7990), .Y(n5414) );
  MX4X1 U3278 ( .A(n5668), .B(n5626), .C(n5647), .D(n5605), .S0(n7993), .S1(
        n7990), .Y(n5669) );
  MX4X1 U3279 ( .A(n6009), .B(n5839), .C(n5924), .D(n5754), .S0(N87), .S1(N86), 
        .Y(N1312) );
  MX4X1 U3280 ( .A(n5838), .B(n5796), .C(n5817), .D(n5775), .S0(n7993), .S1(
        n7990), .Y(n5839) );
  MX4X1 U3281 ( .A(n5753), .B(n5711), .C(n5732), .D(n5690), .S0(n7993), .S1(
        n7990), .Y(n5754) );
  MX4X1 U3282 ( .A(n6008), .B(n5966), .C(n5987), .D(n5945), .S0(n7993), .S1(
        n7990), .Y(n6009) );
  MX4X1 U3283 ( .A(n6349), .B(n6179), .C(n6264), .D(n6094), .S0(N87), .S1(N86), 
        .Y(N1311) );
  MX4X1 U3284 ( .A(n6178), .B(n6136), .C(n6157), .D(n6115), .S0(n7993), .S1(
        n7990), .Y(n6179) );
  MX4X1 U3285 ( .A(n6093), .B(n6051), .C(n6072), .D(n6030), .S0(n7993), .S1(
        n7990), .Y(n6094) );
  MX4X1 U3286 ( .A(n6348), .B(n6306), .C(n6327), .D(n6285), .S0(n7993), .S1(
        n7991), .Y(n6349) );
  MX4X1 U3287 ( .A(n6689), .B(n6519), .C(n6604), .D(n6434), .S0(N87), .S1(N86), 
        .Y(N1310) );
  MX4X1 U3288 ( .A(n6518), .B(n6476), .C(n6497), .D(n6455), .S0(n7993), .S1(
        n7991), .Y(n6519) );
  MX4X1 U3289 ( .A(n6433), .B(n6391), .C(n6412), .D(n6370), .S0(n7992), .S1(
        n7991), .Y(n6434) );
  MX4X1 U3290 ( .A(n6688), .B(n6646), .C(n6667), .D(n6625), .S0(N85), .S1(
        n7991), .Y(n6689) );
  MX4X1 U3291 ( .A(n7029), .B(n6859), .C(n6944), .D(n6774), .S0(N87), .S1(N86), 
        .Y(N1309) );
  MX4X1 U3292 ( .A(n6858), .B(n6816), .C(n6837), .D(n6795), .S0(N85), .S1(
        n7991), .Y(n6859) );
  MX4X1 U3293 ( .A(n6773), .B(n6731), .C(n6752), .D(n6710), .S0(n7992), .S1(
        n7991), .Y(n6774) );
  MX4X1 U3294 ( .A(n7028), .B(n6986), .C(n7007), .D(n6965), .S0(N85), .S1(
        n7991), .Y(n7029) );
  MX4X1 U3295 ( .A(n7369), .B(n7199), .C(n7284), .D(n7114), .S0(N87), .S1(N86), 
        .Y(N1308) );
  MX4X1 U3296 ( .A(n7198), .B(n7156), .C(n7177), .D(n7135), .S0(N85), .S1(
        n7991), .Y(n7199) );
  MX4X1 U3297 ( .A(n7113), .B(n7071), .C(n7092), .D(n7050), .S0(n7992), .S1(
        n7991), .Y(n7114) );
  MX4X1 U3298 ( .A(n7368), .B(n7326), .C(n7347), .D(n7305), .S0(N85), .S1(
        n7991), .Y(n7369) );
  AOI21X1 U3299 ( .A0(n1257), .A1(N1195), .B0(n1261), .Y(n1259) );
  BUFX3 U3300 ( .A(n1244), .Y(n8441) );
  NOR2BXL U3301 ( .AN(n1257), .B(N1195), .Y(n1244) );
  MX4X1 U3302 ( .A(n5583), .B(n5541), .C(n5562), .D(n5520), .S0(n7993), .S1(
        n7990), .Y(n5584) );
  MX4X1 U3303 ( .A(n5540), .B(n5530), .C(n5535), .D(n5525), .S0(n8642), .S1(
        n7974), .Y(n5541) );
  MX4X1 U3304 ( .A(n5519), .B(n5509), .C(n5514), .D(n5504), .S0(n7983), .S1(
        n7974), .Y(n5520) );
  MX4X1 U3305 ( .A(n5582), .B(n5572), .C(n5577), .D(n5567), .S0(n7980), .S1(
        n7974), .Y(n5583) );
  MX4X1 U3306 ( .A(n5923), .B(n5881), .C(n5902), .D(n5860), .S0(n7993), .S1(
        n7990), .Y(n5924) );
  MX4X1 U3307 ( .A(n5880), .B(n5870), .C(n5875), .D(n5865), .S0(n7984), .S1(
        n7975), .Y(n5881) );
  MX4X1 U3308 ( .A(n5859), .B(n5849), .C(n5854), .D(n5844), .S0(n7984), .S1(
        n7975), .Y(n5860) );
  MX4X1 U3309 ( .A(n5922), .B(n5912), .C(n5917), .D(n5907), .S0(n7984), .S1(
        n7975), .Y(n5923) );
  MX4X1 U3310 ( .A(n6263), .B(n6221), .C(n6242), .D(n6200), .S0(n7993), .S1(
        n7990), .Y(n6264) );
  MX4X1 U3311 ( .A(n6220), .B(n6210), .C(n6215), .D(n6205), .S0(n7985), .S1(
        n7976), .Y(n6221) );
  MX4X1 U3312 ( .A(n6199), .B(n6189), .C(n6194), .D(n6184), .S0(n7985), .S1(
        n7976), .Y(n6200) );
  MX4X1 U3313 ( .A(n6262), .B(n6252), .C(n6257), .D(n6247), .S0(n7985), .S1(
        n7976), .Y(n6263) );
  MX4X1 U3314 ( .A(n6603), .B(n6561), .C(n6582), .D(n6540), .S0(n7992), .S1(
        n7991), .Y(n6604) );
  MX4X1 U3315 ( .A(n6560), .B(n6550), .C(n6555), .D(n6545), .S0(n7986), .S1(
        n7974), .Y(n6561) );
  MX4X1 U3316 ( .A(n6539), .B(n6529), .C(n6534), .D(n6524), .S0(n7986), .S1(
        n7977), .Y(n6540) );
  MX4X1 U3317 ( .A(n6602), .B(n6592), .C(n6597), .D(n6587), .S0(n7986), .S1(
        n7973), .Y(n6603) );
  MX4X1 U3318 ( .A(n6943), .B(n6901), .C(n6922), .D(n6880), .S0(n7993), .S1(
        n7991), .Y(n6944) );
  MX4X1 U3319 ( .A(n6900), .B(n6890), .C(n6895), .D(n6885), .S0(n7988), .S1(
        n7972), .Y(n6901) );
  MX4X1 U3320 ( .A(n6879), .B(n6869), .C(n6874), .D(n6864), .S0(n7988), .S1(
        N82), .Y(n6880) );
  MX4X1 U3321 ( .A(n6942), .B(n6932), .C(n6937), .D(n6927), .S0(n7988), .S1(
        n7976), .Y(n6943) );
  MX4X1 U3322 ( .A(n7283), .B(n7241), .C(n7262), .D(n7220), .S0(n7992), .S1(
        n7991), .Y(n7284) );
  MX4X1 U3323 ( .A(n7282), .B(n7272), .C(n7277), .D(n7267), .S0(n7983), .S1(
        n7978), .Y(n7283) );
  MX4X1 U3324 ( .A(n7240), .B(n7230), .C(n7235), .D(n7225), .S0(N83), .S1(
        n8644), .Y(n7241) );
  MX4X1 U3325 ( .A(n7219), .B(n7209), .C(n7214), .D(n7204), .S0(n7987), .S1(
        n7977), .Y(n7220) );
  MX4X1 U3326 ( .A(n5243), .B(n5201), .C(n5222), .D(n5180), .S0(n7992), .S1(
        n7990), .Y(n5244) );
  MX4X1 U3327 ( .A(n5200), .B(n5190), .C(n5195), .D(n5185), .S0(n7982), .S1(
        n7973), .Y(n5201) );
  MX4X1 U3328 ( .A(n5179), .B(n5169), .C(n5174), .D(n5164), .S0(n7982), .S1(
        n7973), .Y(n5180) );
  MX4X1 U3329 ( .A(n5242), .B(n5232), .C(n5237), .D(n5227), .S0(n7982), .S1(
        n7973), .Y(n5243) );
  MX4X1 U3330 ( .A(n4903), .B(n4861), .C(n4882), .D(n4840), .S0(n7992), .S1(
        n7991), .Y(n4904) );
  MX4X1 U3331 ( .A(n4860), .B(n4850), .C(n4855), .D(n4845), .S0(n7981), .S1(
        n7971), .Y(n4861) );
  MX4X1 U3332 ( .A(n4839), .B(n4829), .C(n4834), .D(n4824), .S0(n7981), .S1(
        n7971), .Y(n4840) );
  MX4X1 U3333 ( .A(n4902), .B(n4892), .C(n4897), .D(n4887), .S0(n7981), .S1(
        n7972), .Y(n4903) );
  MX4X1 U3334 ( .A(n1432), .B(n1422), .C(n1427), .D(n1417), .S0(n4637), .S1(
        n4634), .Y(n1433) );
  MX4X1 U3335 ( .A(n1421), .B(n1419), .C(n1420), .D(n1418), .S0(n4616), .S1(
        n4528), .Y(n1422) );
  MX4X1 U3336 ( .A(n1416), .B(n1414), .C(n1415), .D(n1413), .S0(n4610), .S1(
        n4528), .Y(n1417) );
  MX4X1 U3337 ( .A(n1431), .B(n1429), .C(n1430), .D(n1428), .S0(n4618), .S1(
        n4528), .Y(n1432) );
  MX4X1 U3338 ( .A(n1523), .B(n1513), .C(n1518), .D(n1508), .S0(n4637), .S1(
        n4631), .Y(n1524) );
  MX4X1 U3339 ( .A(n1512), .B(n1510), .C(n1511), .D(n1509), .S0(n4588), .S1(
        n4530), .Y(n1513) );
  MX4X1 U3340 ( .A(n1507), .B(n1504), .C(n1506), .D(n1502), .S0(n4588), .S1(
        n4529), .Y(n1508) );
  MX4X1 U3341 ( .A(n1522), .B(n1520), .C(n1521), .D(n1519), .S0(n4588), .S1(
        n4530), .Y(n1523) );
  MX4X1 U3342 ( .A(n1790), .B(n1780), .C(n1785), .D(n1775), .S0(n4638), .S1(
        n4628), .Y(n1791) );
  MX4X1 U3343 ( .A(n1779), .B(n1777), .C(n1778), .D(n1776), .S0(n4592), .S1(
        n4533), .Y(n1780) );
  MX4X1 U3344 ( .A(n1774), .B(n1771), .C(n1772), .D(n1770), .S0(n4592), .S1(
        n4533), .Y(n1775) );
  MX4X1 U3345 ( .A(n1789), .B(n1787), .C(n1788), .D(n1786), .S0(n4592), .S1(
        n4533), .Y(n1790) );
  MX4X1 U3346 ( .A(n1879), .B(n1867), .C(n1874), .D(n1862), .S0(n4638), .S1(
        n4628), .Y(n1880) );
  MX4X1 U3347 ( .A(n1866), .B(n1864), .C(n1865), .D(n1863), .S0(n4593), .S1(
        n4534), .Y(n1867) );
  MX4X1 U3348 ( .A(n1861), .B(n1859), .C(n1860), .D(n1858), .S0(n4593), .S1(
        n4534), .Y(n1862) );
  MX4X1 U3349 ( .A(n1878), .B(n1876), .C(n1877), .D(n1875), .S0(n4593), .S1(
        n4535), .Y(n1879) );
  MX4X1 U3350 ( .A(n1615), .B(n1602), .C(n1610), .D(n1597), .S0(n4637), .S1(
        n4628), .Y(n1616) );
  MX4X1 U3351 ( .A(n1601), .B(n1599), .C(n1600), .D(n1598), .S0(n4589), .S1(
        n4531), .Y(n1602) );
  MX4X1 U3352 ( .A(n1596), .B(n1594), .C(n1595), .D(n1593), .S0(n4589), .S1(
        n4531), .Y(n1597) );
  MX4X1 U3353 ( .A(n1614), .B(n1612), .C(n1613), .D(n1611), .S0(n4589), .S1(
        n4531), .Y(n1615) );
  MX4X1 U3354 ( .A(n1702), .B(n1692), .C(n1697), .D(n1687), .S0(n4638), .S1(
        n4631), .Y(n1703) );
  MX4X1 U3355 ( .A(n1691), .B(n1689), .C(n1690), .D(n1688), .S0(n4590), .S1(
        n4532), .Y(n1692) );
  MX4X1 U3356 ( .A(n1686), .B(n1684), .C(n1685), .D(n1683), .S0(n4590), .S1(
        n4532), .Y(n1687) );
  MX4X1 U3357 ( .A(n1701), .B(n1699), .C(n1700), .D(n1698), .S0(n4590), .S1(
        n4532), .Y(n1702) );
  MX4X1 U3358 ( .A(n2143), .B(n2131), .C(n2137), .D(n2126), .S0(n4639), .S1(
        n4629), .Y(n2144) );
  MX4X1 U3359 ( .A(n2130), .B(n2128), .C(n2129), .D(n2127), .S0(n4597), .S1(
        n4538), .Y(n2131) );
  MX4X1 U3360 ( .A(n2125), .B(n2123), .C(n2124), .D(n2122), .S0(n4597), .S1(
        n4538), .Y(n2126) );
  MX4X1 U3361 ( .A(n2142), .B(n2140), .C(n2141), .D(n2139), .S0(n4597), .S1(
        n4538), .Y(n2143) );
  MX4X1 U3362 ( .A(n2230), .B(n2220), .C(n2225), .D(n2215), .S0(n4640), .S1(
        n4629), .Y(n2231) );
  MX4X1 U3363 ( .A(n2219), .B(n2217), .C(n2218), .D(n2216), .S0(n4598), .S1(
        n4539), .Y(n2220) );
  MX4X1 U3364 ( .A(n2214), .B(n2212), .C(n2213), .D(n2211), .S0(n4598), .S1(
        n4539), .Y(n2215) );
  MX4X1 U3365 ( .A(n2229), .B(n2227), .C(n2228), .D(n2226), .S0(n4598), .S1(
        n4540), .Y(n2230) );
  MX4X1 U3366 ( .A(n1966), .B(n1956), .C(n1961), .D(n1951), .S0(n4639), .S1(
        n4628), .Y(n1967) );
  MX4X1 U3367 ( .A(n1955), .B(n1953), .C(n1954), .D(n1952), .S0(n4594), .S1(
        n4536), .Y(n1956) );
  MX4X1 U3368 ( .A(n1950), .B(n1948), .C(n1949), .D(n1947), .S0(n4594), .S1(
        n4536), .Y(n1951) );
  MX4X1 U3369 ( .A(n1965), .B(n1963), .C(n1964), .D(n1962), .S0(n4594), .S1(
        n4536), .Y(n1966) );
  MX4X1 U3370 ( .A(n2054), .B(n2044), .C(n2049), .D(n2039), .S0(n4639), .S1(
        n4629), .Y(n2055) );
  MX4X1 U3371 ( .A(n2043), .B(n2041), .C(n2042), .D(n2040), .S0(n4596), .S1(
        n4537), .Y(n2044) );
  MX4X1 U3372 ( .A(n2037), .B(n2035), .C(n2036), .D(n2034), .S0(n4596), .S1(
        n4537), .Y(n2039) );
  MX4X1 U3373 ( .A(n2053), .B(n2051), .C(n2052), .D(n2050), .S0(n4596), .S1(
        n4537), .Y(n2054) );
  MX4X1 U3374 ( .A(n2556), .B(n2546), .C(n2551), .D(n2541), .S0(n4641), .S1(
        n4630), .Y(n2557) );
  MX4X1 U3375 ( .A(n2545), .B(n2543), .C(n2544), .D(n2542), .S0(n4602), .S1(
        n4543), .Y(n2546) );
  MX4X1 U3376 ( .A(n2540), .B(n2538), .C(n2539), .D(n2537), .S0(n4602), .S1(
        n4543), .Y(n2541) );
  MX4X1 U3377 ( .A(n2555), .B(n2553), .C(n2554), .D(n2552), .S0(n4602), .S1(
        n4543), .Y(n2556) );
  MX4X1 U3378 ( .A(n2641), .B(n2631), .C(n2636), .D(n2626), .S0(n4641), .S1(
        n4630), .Y(n2642) );
  MX4X1 U3379 ( .A(n2630), .B(n2628), .C(n2629), .D(n2627), .S0(n4604), .S1(
        n4545), .Y(n2631) );
  MX4X1 U3380 ( .A(n2625), .B(n2623), .C(n2624), .D(n2622), .S0(n4604), .S1(
        n4540), .Y(n2626) );
  MX4X1 U3381 ( .A(n2640), .B(n2638), .C(n2639), .D(n2637), .S0(n4604), .S1(
        n4536), .Y(n2641) );
  MX4X1 U3382 ( .A(n2318), .B(n2308), .C(n2313), .D(n2302), .S0(n4640), .S1(
        n4630), .Y(n2319) );
  MX4X1 U3383 ( .A(n2307), .B(n2305), .C(n2306), .D(n2304), .S0(n4600), .S1(
        n4541), .Y(n2308) );
  MX4X1 U3384 ( .A(n2301), .B(n2299), .C(n2300), .D(n2298), .S0(n4600), .S1(
        n4541), .Y(n2302) );
  MX4X1 U3385 ( .A(n2317), .B(n2315), .C(n2316), .D(n2314), .S0(n4600), .S1(
        n4541), .Y(n2318) );
  MX4X1 U3386 ( .A(n2471), .B(n2461), .C(n2466), .D(n2456), .S0(n4640), .S1(
        n4630), .Y(n2472) );
  MX4X1 U3387 ( .A(n2460), .B(n2458), .C(n2459), .D(n2457), .S0(n4601), .S1(
        n4542), .Y(n2461) );
  MX4X1 U3388 ( .A(n2455), .B(n2453), .C(n2454), .D(n2452), .S0(n4601), .S1(
        n4542), .Y(n2456) );
  MX4X1 U3389 ( .A(n2470), .B(n2468), .C(n2469), .D(n2467), .S0(n4601), .S1(
        n4542), .Y(n2471) );
  MX4X1 U3390 ( .A(n2896), .B(n2886), .C(n2891), .D(n2881), .S0(n4642), .S1(
        n4631), .Y(n2897) );
  MX4X1 U3391 ( .A(n2885), .B(n2883), .C(n2884), .D(n2882), .S0(n4608), .S1(
        n4547), .Y(n2886) );
  MX4X1 U3392 ( .A(n2880), .B(n2878), .C(n2879), .D(n2877), .S0(n4608), .S1(
        n4547), .Y(n2881) );
  MX4X1 U3393 ( .A(n2895), .B(n2893), .C(n2894), .D(n2892), .S0(n4608), .S1(
        n4547), .Y(n2896) );
  MX4X1 U3394 ( .A(n2981), .B(n2971), .C(n2976), .D(n2966), .S0(n4642), .S1(
        n4632), .Y(n2982) );
  MX4X1 U3395 ( .A(n2970), .B(n2968), .C(n2969), .D(n2967), .S0(n4609), .S1(
        n4548), .Y(n2971) );
  MX4X1 U3396 ( .A(n2965), .B(n2963), .C(n2964), .D(n2962), .S0(n4609), .S1(
        n4548), .Y(n2966) );
  MX4X1 U3397 ( .A(n2980), .B(n2978), .C(n2979), .D(n2977), .S0(n4609), .S1(
        n4548), .Y(n2981) );
  MX4X1 U3398 ( .A(n2726), .B(n2716), .C(n2721), .D(n2711), .S0(n4641), .S1(
        n4631), .Y(n2727) );
  MX4X1 U3399 ( .A(n2715), .B(n2713), .C(n2714), .D(n2712), .S0(n4605), .S1(
        n4545), .Y(n2716) );
  MX4X1 U3400 ( .A(n2710), .B(n2708), .C(n2709), .D(n2707), .S0(n4605), .S1(
        n4544), .Y(n2711) );
  MX4X1 U3401 ( .A(n2725), .B(n2723), .C(n2724), .D(n2722), .S0(n4605), .S1(
        n4545), .Y(n2726) );
  MX4X1 U3402 ( .A(n2811), .B(n2801), .C(n2806), .D(n2796), .S0(n4642), .S1(
        n4631), .Y(n2812) );
  MX4X1 U3403 ( .A(n2800), .B(n2798), .C(n2799), .D(n2797), .S0(n4606), .S1(
        n4546), .Y(n2801) );
  MX4X1 U3404 ( .A(n2795), .B(n2793), .C(n2794), .D(n2792), .S0(n4606), .S1(
        n4546), .Y(n2796) );
  MX4X1 U3405 ( .A(n2810), .B(n2808), .C(n2809), .D(n2807), .S0(n4606), .S1(
        n4546), .Y(n2811) );
  MX4X1 U3406 ( .A(n3236), .B(n3226), .C(n3231), .D(n3221), .S0(n4643), .S1(
        n4633), .Y(n3237) );
  MX4X1 U3407 ( .A(n3225), .B(n3223), .C(n3224), .D(n3222), .S0(n4613), .S1(
        n4552), .Y(n3226) );
  MX4X1 U3408 ( .A(n3220), .B(n3218), .C(n3219), .D(n3217), .S0(n4613), .S1(
        n4552), .Y(n3221) );
  MX4X1 U3409 ( .A(n3235), .B(n3233), .C(n3234), .D(n3232), .S0(n4613), .S1(
        n4552), .Y(n3236) );
  MX4X1 U3410 ( .A(n3321), .B(n3311), .C(n3316), .D(n3306), .S0(n4644), .S1(
        n4633), .Y(n3322) );
  MX4X1 U3411 ( .A(n3310), .B(n3308), .C(n3309), .D(n3307), .S0(n4614), .S1(
        n4553), .Y(n3311) );
  MX4X1 U3412 ( .A(n3305), .B(n3303), .C(n3304), .D(n3302), .S0(n4614), .S1(
        n4553), .Y(n3306) );
  MX4X1 U3413 ( .A(n3320), .B(n3318), .C(n3319), .D(n3317), .S0(n4614), .S1(
        n4553), .Y(n3321) );
  MX4X1 U3414 ( .A(n3066), .B(n3056), .C(n3061), .D(n3051), .S0(n4643), .S1(
        n4632), .Y(n3067) );
  MX4X1 U3415 ( .A(n3055), .B(n3053), .C(n3054), .D(n3052), .S0(n4610), .S1(
        n4549), .Y(n3056) );
  MX4X1 U3416 ( .A(n3050), .B(n3048), .C(n3049), .D(n3047), .S0(n4610), .S1(
        n4549), .Y(n3051) );
  MX4X1 U3417 ( .A(n3065), .B(n3063), .C(n3064), .D(n3062), .S0(n4610), .S1(
        n4550), .Y(n3066) );
  MX4X1 U3418 ( .A(n3151), .B(n3141), .C(n3146), .D(n3136), .S0(n4643), .S1(
        n4632), .Y(n3152) );
  MX4X1 U3419 ( .A(n3140), .B(n3138), .C(n3139), .D(n3137), .S0(n4612), .S1(
        n4551), .Y(n3141) );
  MX4X1 U3420 ( .A(n3135), .B(n3133), .C(n3134), .D(n3132), .S0(n4612), .S1(
        n4551), .Y(n3136) );
  MX4X1 U3421 ( .A(n3150), .B(n3148), .C(n3149), .D(n3147), .S0(n4612), .S1(
        n4551), .Y(n3151) );
  MX4X1 U3422 ( .A(n3576), .B(n3566), .C(n3571), .D(n3561), .S0(n4640), .S1(
        n4634), .Y(n3577) );
  MX4X1 U3423 ( .A(n3565), .B(n3563), .C(n3564), .D(n3562), .S0(n4618), .S1(
        n4557), .Y(n3566) );
  MX4X1 U3424 ( .A(n3560), .B(n3558), .C(n3559), .D(n3557), .S0(n4618), .S1(
        n4557), .Y(n3561) );
  MX4X1 U3425 ( .A(n3575), .B(n3573), .C(n3574), .D(n3572), .S0(n4618), .S1(
        n4557), .Y(n3576) );
  MX4X1 U3426 ( .A(n3661), .B(n3651), .C(n3656), .D(n3646), .S0(n4639), .S1(
        n4634), .Y(n3662) );
  MX4X1 U3427 ( .A(n3650), .B(n3648), .C(n3649), .D(n3647), .S0(n4620), .S1(
        n4560), .Y(n3651) );
  MX4X1 U3428 ( .A(n3645), .B(n3643), .C(n3644), .D(n3642), .S0(n4620), .S1(
        N70), .Y(n3646) );
  MX4X1 U3429 ( .A(n3660), .B(n3658), .C(n3659), .D(n3657), .S0(n4620), .S1(
        N70), .Y(n3661) );
  MX4X1 U3430 ( .A(n3406), .B(n3396), .C(n3401), .D(n3391), .S0(n4644), .S1(
        n4633), .Y(n3407) );
  MX4X1 U3431 ( .A(n3395), .B(n3393), .C(n3394), .D(n3392), .S0(n4616), .S1(
        n4554), .Y(n3396) );
  MX4X1 U3432 ( .A(n3390), .B(n3388), .C(n3389), .D(n3387), .S0(n4616), .S1(
        n4554), .Y(n3391) );
  MX4X1 U3433 ( .A(n3405), .B(n3403), .C(n3404), .D(n3402), .S0(n4616), .S1(
        n4555), .Y(n3406) );
  MX4X1 U3434 ( .A(n3491), .B(n3481), .C(n3486), .D(n3476), .S0(n4644), .S1(
        n4634), .Y(n3492) );
  MX4X1 U3435 ( .A(n3480), .B(n3478), .C(n3479), .D(n3477), .S0(n4617), .S1(
        n4556), .Y(n3481) );
  MX4X1 U3436 ( .A(n3475), .B(n3473), .C(n3474), .D(n3472), .S0(n4617), .S1(
        n4556), .Y(n3476) );
  MX4X1 U3437 ( .A(n3490), .B(n3488), .C(n3489), .D(n3487), .S0(n4617), .S1(
        n4556), .Y(n3491) );
  MX4X1 U3438 ( .A(n3916), .B(n3906), .C(n3911), .D(n3901), .S0(n4645), .S1(
        n4635), .Y(n3917) );
  MX4X1 U3439 ( .A(n3905), .B(n3903), .C(n3904), .D(n3902), .S0(n4624), .S1(
        n4558), .Y(n3906) );
  MX4X1 U3440 ( .A(n3900), .B(n3898), .C(n3899), .D(n3897), .S0(n4624), .S1(
        n4558), .Y(n3901) );
  MX4X1 U3441 ( .A(n3915), .B(n3913), .C(n3914), .D(n3912), .S0(n4624), .S1(
        n4558), .Y(n3916) );
  MX4X1 U3442 ( .A(n4001), .B(n3991), .C(n3996), .D(n3986), .S0(n4645), .S1(
        n4635), .Y(n4002) );
  MX4X1 U3443 ( .A(n3990), .B(n3988), .C(n3989), .D(n3987), .S0(n4568), .S1(
        n4559), .Y(n3991) );
  MX4X1 U3444 ( .A(n3985), .B(n3983), .C(n3984), .D(n3982), .S0(n4569), .S1(
        n4559), .Y(n3986) );
  MX4X1 U3445 ( .A(n4000), .B(n3998), .C(n3999), .D(n3997), .S0(N71), .S1(
        n4559), .Y(n4001) );
  MX4X1 U3446 ( .A(n3746), .B(n3736), .C(n3741), .D(n3731), .S0(n4644), .S1(
        n4634), .Y(n3747) );
  MX4X1 U3447 ( .A(n3735), .B(n3733), .C(n3734), .D(n3732), .S0(n4621), .S1(
        n4528), .Y(n3736) );
  MX4X1 U3448 ( .A(n3730), .B(n3728), .C(n3729), .D(n3727), .S0(n4621), .S1(
        n4533), .Y(n3731) );
  MX4X1 U3449 ( .A(n3745), .B(n3743), .C(n3744), .D(n3742), .S0(n4621), .S1(
        n4559), .Y(n3746) );
  MX4X1 U3450 ( .A(n3831), .B(n3821), .C(n3826), .D(n3816), .S0(n4645), .S1(
        n4635), .Y(n3832) );
  MX4X1 U3451 ( .A(n3820), .B(n3818), .C(n3819), .D(n3817), .S0(n4622), .S1(
        n4535), .Y(n3821) );
  MX4X1 U3452 ( .A(n3815), .B(n3813), .C(n3814), .D(n3812), .S0(n4622), .S1(
        n4541), .Y(n3816) );
  MX4X1 U3453 ( .A(n3830), .B(n3828), .C(n3829), .D(n3827), .S0(n4622), .S1(
        n4545), .Y(n3831) );
  MX4X1 U3454 ( .A(n4881), .B(n4871), .C(n4876), .D(n4866), .S0(n7981), .S1(
        n7971), .Y(n4882) );
  MX4X1 U3455 ( .A(n4870), .B(n4868), .C(n4869), .D(n4867), .S0(n7959), .S1(
        n7869), .Y(n4871) );
  MX4X1 U3456 ( .A(n4865), .B(n4863), .C(n4864), .D(n4862), .S0(n7953), .S1(
        n7869), .Y(n4866) );
  MX4X1 U3457 ( .A(n4880), .B(n4878), .C(n4879), .D(n4877), .S0(n7961), .S1(
        n7869), .Y(n4881) );
  MX4X1 U3458 ( .A(n4966), .B(n4956), .C(n4961), .D(n4951), .S0(n7981), .S1(
        n7972), .Y(n4967) );
  MX4X1 U3459 ( .A(n4955), .B(n4953), .C(n4954), .D(n4952), .S0(n7931), .S1(
        n7871), .Y(n4956) );
  MX4X1 U3460 ( .A(n4950), .B(n4948), .C(n4949), .D(n4947), .S0(n7931), .S1(
        n7870), .Y(n4951) );
  MX4X1 U3461 ( .A(n4965), .B(n4963), .C(n4964), .D(n4962), .S0(n7931), .S1(
        n7871), .Y(n4966) );
  MX4X1 U3462 ( .A(n5221), .B(n5211), .C(n5216), .D(n5206), .S0(n7982), .S1(
        n7973), .Y(n5222) );
  MX4X1 U3463 ( .A(n5210), .B(n5208), .C(n5209), .D(n5207), .S0(n7935), .S1(
        n7874), .Y(n5211) );
  MX4X1 U3464 ( .A(n5205), .B(n5203), .C(n5204), .D(n5202), .S0(n7935), .S1(
        n7874), .Y(n5206) );
  MX4X1 U3465 ( .A(n5220), .B(n5218), .C(n5219), .D(n5217), .S0(n7935), .S1(
        n7874), .Y(n5221) );
  MX4X1 U3466 ( .A(n5306), .B(n5296), .C(n5301), .D(n5291), .S0(n7982), .S1(
        n7973), .Y(n5307) );
  MX4X1 U3467 ( .A(n5295), .B(n5293), .C(n5294), .D(n5292), .S0(n7936), .S1(
        n7875), .Y(n5296) );
  MX4X1 U3468 ( .A(n5290), .B(n5288), .C(n5289), .D(n5287), .S0(n7936), .S1(
        n7875), .Y(n5291) );
  MX4X1 U3469 ( .A(n5305), .B(n5303), .C(n5304), .D(n5302), .S0(n7936), .S1(
        n7876), .Y(n5306) );
  MX4X1 U3470 ( .A(n5051), .B(n5041), .C(n5046), .D(n5036), .S0(n7981), .S1(
        n7972), .Y(n5052) );
  MX4X1 U3471 ( .A(n5040), .B(n5038), .C(n5039), .D(n5037), .S0(n7932), .S1(
        n7872), .Y(n5041) );
  MX4X1 U3472 ( .A(n5035), .B(n5033), .C(n5034), .D(n5032), .S0(n7932), .S1(
        n7872), .Y(n5036) );
  MX4X1 U3473 ( .A(n5050), .B(n5048), .C(n5049), .D(n5047), .S0(n7932), .S1(
        n7872), .Y(n5051) );
  MX4X1 U3474 ( .A(n5136), .B(n5126), .C(n5131), .D(n5121), .S0(n7982), .S1(
        n7972), .Y(n5137) );
  MX4X1 U3475 ( .A(n5125), .B(n5123), .C(n5124), .D(n5122), .S0(n7933), .S1(
        n7873), .Y(n5126) );
  MX4X1 U3476 ( .A(n5120), .B(n5118), .C(n5119), .D(n5117), .S0(n7933), .S1(
        n7873), .Y(n5121) );
  MX4X1 U3477 ( .A(n5135), .B(n5133), .C(n5134), .D(n5132), .S0(n7933), .S1(
        n7873), .Y(n5136) );
  MX4X1 U3478 ( .A(n5561), .B(n5551), .C(n5556), .D(n5546), .S0(n7986), .S1(
        n7974), .Y(n5562) );
  MX4X1 U3479 ( .A(n5550), .B(n5548), .C(n5549), .D(n5547), .S0(n7940), .S1(
        n7879), .Y(n5551) );
  MX4X1 U3480 ( .A(n5545), .B(n5543), .C(n5544), .D(n5542), .S0(n7940), .S1(
        n7879), .Y(n5546) );
  MX4X1 U3481 ( .A(n5560), .B(n5558), .C(n5559), .D(n5557), .S0(n7940), .S1(
        n7879), .Y(n5561) );
  MX4X1 U3482 ( .A(n5646), .B(n5636), .C(n5641), .D(n5631), .S0(n7983), .S1(
        n7974), .Y(n5647) );
  MX4X1 U3483 ( .A(n5635), .B(n5633), .C(n5634), .D(n5632), .S0(n7941), .S1(
        n7880), .Y(n5636) );
  MX4X1 U3484 ( .A(n5630), .B(n5628), .C(n5629), .D(n5627), .S0(n7941), .S1(
        n7880), .Y(n5631) );
  MX4X1 U3485 ( .A(n5645), .B(n5643), .C(n5644), .D(n5642), .S0(n7941), .S1(
        n7881), .Y(n5646) );
  MX4X1 U3486 ( .A(n5391), .B(n5381), .C(n5386), .D(n5376), .S0(n7984), .S1(
        n7973), .Y(n5392) );
  MX4X1 U3487 ( .A(n5380), .B(n5378), .C(n5379), .D(n5377), .S0(n7937), .S1(
        n7877), .Y(n5381) );
  MX4X1 U3488 ( .A(n5375), .B(n5373), .C(n5374), .D(n5372), .S0(n7937), .S1(
        n7877), .Y(n5376) );
  MX4X1 U3489 ( .A(n5390), .B(n5388), .C(n5389), .D(n5387), .S0(n7937), .S1(
        n7877), .Y(n5391) );
  MX4X1 U3490 ( .A(n5476), .B(n5466), .C(n5471), .D(n5461), .S0(n8642), .S1(
        n7974), .Y(n5477) );
  MX4X1 U3491 ( .A(n5465), .B(n5463), .C(n5464), .D(n5462), .S0(n7939), .S1(
        n7878), .Y(n5466) );
  MX4X1 U3492 ( .A(n5460), .B(n5458), .C(n5459), .D(n5457), .S0(n7939), .S1(
        n7878), .Y(n5461) );
  MX4X1 U3493 ( .A(n5475), .B(n5473), .C(n5474), .D(n5472), .S0(n7939), .S1(
        n7878), .Y(n5476) );
  MX4X1 U3494 ( .A(n5901), .B(n5891), .C(n5896), .D(n5886), .S0(n7984), .S1(
        n7975), .Y(n5902) );
  MX4X1 U3495 ( .A(n5890), .B(n5888), .C(n5889), .D(n5887), .S0(n7945), .S1(
        n7884), .Y(n5891) );
  MX4X1 U3496 ( .A(n5885), .B(n5883), .C(n5884), .D(n5882), .S0(n7945), .S1(
        n7884), .Y(n5886) );
  MX4X1 U3497 ( .A(n5900), .B(n5898), .C(n5899), .D(n5897), .S0(n7945), .S1(
        n7884), .Y(n5901) );
  MX4X1 U3498 ( .A(n5986), .B(n5976), .C(n5981), .D(n5971), .S0(n7984), .S1(
        n7975), .Y(n5987) );
  MX4X1 U3499 ( .A(n5975), .B(n5973), .C(n5974), .D(n5972), .S0(n7947), .S1(
        n7885), .Y(n5976) );
  MX4X1 U3500 ( .A(n5970), .B(n5968), .C(n5969), .D(n5967), .S0(n7947), .S1(
        n7885), .Y(n5971) );
  MX4X1 U3501 ( .A(n5985), .B(n5983), .C(n5984), .D(n5982), .S0(n7947), .S1(
        n7885), .Y(n5986) );
  MX4X1 U3502 ( .A(n5731), .B(n5721), .C(n5726), .D(n5716), .S0(n7983), .S1(
        n7975), .Y(n5732) );
  MX4X1 U3503 ( .A(n5720), .B(n5718), .C(n5719), .D(n5717), .S0(n7943), .S1(
        n7882), .Y(n5721) );
  MX4X1 U3504 ( .A(n5715), .B(n5713), .C(n5714), .D(n5712), .S0(n7943), .S1(
        n7882), .Y(n5716) );
  MX4X1 U3505 ( .A(n5730), .B(n5728), .C(n5729), .D(n5727), .S0(n7943), .S1(
        n7882), .Y(n5731) );
  MX4X1 U3506 ( .A(n5816), .B(n5806), .C(n5811), .D(n5801), .S0(n7983), .S1(
        n7975), .Y(n5817) );
  MX4X1 U3507 ( .A(n5805), .B(n5803), .C(n5804), .D(n5802), .S0(n7944), .S1(
        n7883), .Y(n5806) );
  MX4X1 U3508 ( .A(n5800), .B(n5798), .C(n5799), .D(n5797), .S0(n7944), .S1(
        n7883), .Y(n5801) );
  MX4X1 U3509 ( .A(n5815), .B(n5813), .C(n5814), .D(n5812), .S0(n7944), .S1(
        n7883), .Y(n5816) );
  MX4X1 U3510 ( .A(n6241), .B(n6231), .C(n6236), .D(n6226), .S0(n7985), .S1(
        n7976), .Y(n6242) );
  MX4X1 U3511 ( .A(n6230), .B(n6228), .C(n6229), .D(n6227), .S0(n7951), .S1(
        n7889), .Y(n6231) );
  MX4X1 U3512 ( .A(n6225), .B(n6223), .C(n6224), .D(n6222), .S0(n7951), .S1(
        n7889), .Y(n6226) );
  MX4X1 U3513 ( .A(n6240), .B(n6238), .C(n6239), .D(n6237), .S0(n7951), .S1(
        n7889), .Y(n6241) );
  MX4X1 U3514 ( .A(n6326), .B(n6316), .C(n6321), .D(n6311), .S0(n7985), .S1(
        n7977), .Y(n6327) );
  MX4X1 U3515 ( .A(n6315), .B(n6313), .C(n6314), .D(n6312), .S0(n7952), .S1(
        n7890), .Y(n6316) );
  MX4X1 U3516 ( .A(n6310), .B(n6308), .C(n6309), .D(n6307), .S0(n7952), .S1(
        n7890), .Y(n6311) );
  MX4X1 U3517 ( .A(n6325), .B(n6323), .C(n6324), .D(n6322), .S0(n7952), .S1(
        n7890), .Y(n6326) );
  MX4X1 U3518 ( .A(n6071), .B(n6061), .C(n6066), .D(n6056), .S0(n7984), .S1(
        n7976), .Y(n6072) );
  MX4X1 U3519 ( .A(n6060), .B(n6058), .C(n6059), .D(n6057), .S0(n7948), .S1(
        n7887), .Y(n6061) );
  MX4X1 U3520 ( .A(n6055), .B(n6053), .C(n6054), .D(n6052), .S0(n7948), .S1(
        n7886), .Y(n6056) );
  MX4X1 U3521 ( .A(n6070), .B(n6068), .C(n6069), .D(n6067), .S0(n7948), .S1(
        n7887), .Y(n6071) );
  MX4X1 U3522 ( .A(n6156), .B(n6146), .C(n6151), .D(n6141), .S0(n7985), .S1(
        n7976), .Y(n6157) );
  MX4X1 U3523 ( .A(n6145), .B(n6143), .C(n6144), .D(n6142), .S0(n7949), .S1(
        n7888), .Y(n6146) );
  MX4X1 U3524 ( .A(n6140), .B(n6138), .C(n6139), .D(n6137), .S0(n7949), .S1(
        n7888), .Y(n6141) );
  MX4X1 U3525 ( .A(n6155), .B(n6153), .C(n6154), .D(n6152), .S0(n7949), .S1(
        n7888), .Y(n6156) );
  MX4X1 U3526 ( .A(n6581), .B(n6571), .C(n6576), .D(n6566), .S0(n7986), .S1(
        n7973), .Y(n6582) );
  MX4X1 U3527 ( .A(n6570), .B(n6568), .C(n6569), .D(n6567), .S0(n7956), .S1(
        n7894), .Y(n6571) );
  MX4X1 U3528 ( .A(n6565), .B(n6563), .C(n6564), .D(n6562), .S0(n7956), .S1(
        n7894), .Y(n6566) );
  MX4X1 U3529 ( .A(n6580), .B(n6578), .C(n6579), .D(n6577), .S0(n7956), .S1(
        n7894), .Y(n6581) );
  MX4X1 U3530 ( .A(n6666), .B(n6656), .C(n6661), .D(n6651), .S0(n7987), .S1(
        n7975), .Y(n6667) );
  MX4X1 U3531 ( .A(n6655), .B(n6653), .C(n6654), .D(n6652), .S0(n7957), .S1(
        n7895), .Y(n6656) );
  MX4X1 U3532 ( .A(n6650), .B(n6648), .C(n6649), .D(n6647), .S0(n7957), .S1(
        n7895), .Y(n6651) );
  MX4X1 U3533 ( .A(n6665), .B(n6663), .C(n6664), .D(n6662), .S0(n7957), .S1(
        n7895), .Y(n6666) );
  MX4X1 U3534 ( .A(n6411), .B(n6401), .C(n6406), .D(n6396), .S0(n7986), .S1(
        n7977), .Y(n6412) );
  MX4X1 U3535 ( .A(n6400), .B(n6398), .C(n6399), .D(n6397), .S0(n7953), .S1(
        n7891), .Y(n6401) );
  MX4X1 U3536 ( .A(n6395), .B(n6393), .C(n6394), .D(n6392), .S0(n7953), .S1(
        n7891), .Y(n6396) );
  MX4X1 U3537 ( .A(n6410), .B(n6408), .C(n6409), .D(n6407), .S0(n7953), .S1(
        n7892), .Y(n6411) );
  MX4X1 U3538 ( .A(n6496), .B(n6486), .C(n6491), .D(n6481), .S0(n7986), .S1(
        n7977), .Y(n6497) );
  MX4X1 U3539 ( .A(n6485), .B(n6483), .C(n6484), .D(n6482), .S0(n7955), .S1(
        n7893), .Y(n6486) );
  MX4X1 U3540 ( .A(n6480), .B(n6478), .C(n6479), .D(n6477), .S0(n7955), .S1(
        n7893), .Y(n6481) );
  MX4X1 U3541 ( .A(n6495), .B(n6493), .C(n6494), .D(n6492), .S0(n7955), .S1(
        n7893), .Y(n6496) );
  MX4X1 U3542 ( .A(n6921), .B(n6911), .C(n6916), .D(n6906), .S0(n7988), .S1(
        N82), .Y(n6922) );
  MX4X1 U3543 ( .A(n6910), .B(n6908), .C(n6909), .D(n6907), .S0(n7961), .S1(
        n7897), .Y(n6911) );
  MX4X1 U3544 ( .A(n6905), .B(n6903), .C(n6904), .D(n6902), .S0(n7961), .S1(
        n7897), .Y(n6906) );
  MX4X1 U3545 ( .A(n6920), .B(n6918), .C(n6919), .D(n6917), .S0(n7961), .S1(
        n7897), .Y(n6921) );
  MX4X1 U3546 ( .A(n7006), .B(n6996), .C(n7001), .D(n6991), .S0(n7988), .S1(
        N82), .Y(n7007) );
  MX4X1 U3547 ( .A(n6995), .B(n6993), .C(n6994), .D(n6992), .S0(n7963), .S1(
        n7898), .Y(n6996) );
  MX4X1 U3548 ( .A(n6990), .B(n6988), .C(n6989), .D(n6987), .S0(n7963), .S1(
        n7898), .Y(n6991) );
  MX4X1 U3549 ( .A(n7005), .B(n7003), .C(n7004), .D(n7002), .S0(n7963), .S1(
        n7898), .Y(n7006) );
  MX4X1 U3550 ( .A(n6751), .B(n6741), .C(n6746), .D(n6736), .S0(n7987), .S1(
        n7974), .Y(n6752) );
  MX4X1 U3551 ( .A(n6740), .B(n6738), .C(n6739), .D(n6737), .S0(n7959), .S1(
        n7896), .Y(n6741) );
  MX4X1 U3552 ( .A(n6735), .B(n6733), .C(n6734), .D(n6732), .S0(n7959), .S1(
        n7896), .Y(n6736) );
  MX4X1 U3553 ( .A(n6750), .B(n6748), .C(n6749), .D(n6747), .S0(n7959), .S1(
        n7888), .Y(n6751) );
  MX4X1 U3554 ( .A(n6836), .B(n6826), .C(n6831), .D(n6821), .S0(n7987), .S1(
        n7975), .Y(n6837) );
  MX4X1 U3555 ( .A(n6825), .B(n6823), .C(n6824), .D(n6822), .S0(n7960), .S1(
        n7899), .Y(n6826) );
  MX4X1 U3556 ( .A(n6820), .B(n6818), .C(n6819), .D(n6817), .S0(n7960), .S1(
        n7900), .Y(n6821) );
  MX4X1 U3557 ( .A(n6835), .B(n6833), .C(n6834), .D(n6832), .S0(n7960), .S1(
        n7867), .Y(n6836) );
  MX4X1 U3558 ( .A(n7261), .B(n7251), .C(n7256), .D(n7246), .S0(n7988), .S1(
        N82), .Y(n7262) );
  MX4X1 U3559 ( .A(n7250), .B(n7248), .C(n7249), .D(n7247), .S0(n7967), .S1(
        n7889), .Y(n7251) );
  MX4X1 U3560 ( .A(n7245), .B(n7243), .C(n7244), .D(n7242), .S0(n7967), .S1(
        n7897), .Y(n7246) );
  MX4X1 U3561 ( .A(n7260), .B(n7258), .C(n7259), .D(n7257), .S0(n7967), .S1(
        n7896), .Y(n7261) );
  MX4X1 U3562 ( .A(n7346), .B(n7336), .C(n7341), .D(n7331), .S0(n7984), .S1(
        n7972), .Y(n7347) );
  MX4X1 U3563 ( .A(n7335), .B(n7333), .C(n7334), .D(n7332), .S0(n7910), .S1(
        n7902), .Y(n7336) );
  MX4X1 U3564 ( .A(n7330), .B(n7328), .C(n7329), .D(n7327), .S0(n7911), .S1(
        n7902), .Y(n7331) );
  MX4X1 U3565 ( .A(n7345), .B(n7343), .C(n7344), .D(n7342), .S0(N81), .S1(
        n7902), .Y(n7346) );
  MX4X1 U3566 ( .A(n7091), .B(n7081), .C(n7086), .D(n7076), .S0(n7988), .S1(
        N82), .Y(n7092) );
  MX4X1 U3567 ( .A(n7080), .B(n7078), .C(n7079), .D(n7077), .S0(n7964), .S1(
        n7899), .Y(n7081) );
  MX4X1 U3568 ( .A(n7075), .B(n7073), .C(n7074), .D(n7072), .S0(n7964), .S1(
        n7899), .Y(n7076) );
  MX4X1 U3569 ( .A(n7090), .B(n7088), .C(n7089), .D(n7087), .S0(n7964), .S1(
        n7899), .Y(n7091) );
  MX4X1 U3570 ( .A(n7176), .B(n7166), .C(n7171), .D(n7161), .S0(N83), .S1(
        n7974), .Y(n7177) );
  MX4X1 U3571 ( .A(n7165), .B(n7163), .C(n7164), .D(n7162), .S0(n7965), .S1(
        n7901), .Y(n7166) );
  MX4X1 U3572 ( .A(n7160), .B(n7158), .C(n7159), .D(n7157), .S0(n7965), .S1(
        n7900), .Y(n7161) );
  MX4X1 U3573 ( .A(n7175), .B(n7173), .C(n7174), .D(n7172), .S0(n7965), .S1(
        n7901), .Y(n7176) );
  MX4X1 U3574 ( .A(n2165), .B(n2121), .C(n2144), .D(n2099), .S0(n4649), .S1(
        N74), .Y(n2166) );
  MX4X1 U3575 ( .A(n2120), .B(n2110), .C(n2115), .D(n2105), .S0(n4639), .S1(
        n4629), .Y(n2121) );
  MX4X1 U3576 ( .A(n2098), .B(n2088), .C(n2093), .D(n2083), .S0(n4639), .S1(
        n4629), .Y(n2099) );
  MX4X1 U3577 ( .A(n2164), .B(n2154), .C(n2159), .D(n2149), .S0(n4639), .S1(
        n4629), .Y(n2165) );
  MX4X1 U3578 ( .A(n2578), .B(n2536), .C(n2557), .D(n2515), .S0(n4649), .S1(
        N74), .Y(n2579) );
  MX4X1 U3579 ( .A(n2535), .B(n2525), .C(n2530), .D(n2520), .S0(n4641), .S1(
        n4630), .Y(n2536) );
  MX4X1 U3580 ( .A(n2514), .B(n2504), .C(n2509), .D(n2499), .S0(n4641), .S1(
        n4630), .Y(n2515) );
  MX4X1 U3581 ( .A(n2577), .B(n2567), .C(n2572), .D(n2562), .S0(n4641), .S1(
        n4630), .Y(n2578) );
  MX4X1 U3582 ( .A(n2918), .B(n2876), .C(n2897), .D(n2855), .S0(n4649), .S1(
        N74), .Y(n2919) );
  MX4X1 U3583 ( .A(n2875), .B(n2865), .C(n2870), .D(n2860), .S0(n4642), .S1(
        n4631), .Y(n2876) );
  MX4X1 U3584 ( .A(n2854), .B(n2844), .C(n2849), .D(n2839), .S0(n4642), .S1(
        n4631), .Y(n2855) );
  MX4X1 U3585 ( .A(n2917), .B(n2907), .C(n2912), .D(n2902), .S0(n4642), .S1(
        n4631), .Y(n2918) );
  MX4X1 U3586 ( .A(n3258), .B(n3216), .C(n3237), .D(n3195), .S0(n4648), .S1(
        n4646), .Y(n3259) );
  MX4X1 U3587 ( .A(n3215), .B(n3205), .C(n3210), .D(n3200), .S0(n4643), .S1(
        n4633), .Y(n3216) );
  MX4X1 U3588 ( .A(n3194), .B(n3184), .C(n3189), .D(n3179), .S0(n4643), .S1(
        n4632), .Y(n3195) );
  MX4X1 U3589 ( .A(n3257), .B(n3247), .C(n3252), .D(n3242), .S0(n4643), .S1(
        n4633), .Y(n3258) );
  MX4X1 U3590 ( .A(n3598), .B(n3556), .C(n3577), .D(n3535), .S0(n4649), .S1(
        n4646), .Y(n3599) );
  MX4X1 U3591 ( .A(n3555), .B(n3545), .C(n3550), .D(n3540), .S0(n4643), .S1(
        n4634), .Y(n3556) );
  MX4X1 U3592 ( .A(n3534), .B(n3524), .C(n3529), .D(n3519), .S0(n4639), .S1(
        n4634), .Y(n3535) );
  MX4X1 U3593 ( .A(n3597), .B(n3587), .C(n3592), .D(n3582), .S0(n4643), .S1(
        n4634), .Y(n3598) );
  MX4X1 U3594 ( .A(n3938), .B(n3896), .C(n3917), .D(n3875), .S0(n4648), .S1(
        n4646), .Y(n3939) );
  MX4X1 U3595 ( .A(n3895), .B(n3885), .C(n3890), .D(n3880), .S0(n4645), .S1(
        n4635), .Y(n3896) );
  MX4X1 U3596 ( .A(n3874), .B(n3864), .C(n3869), .D(n3859), .S0(n4645), .S1(
        n4635), .Y(n3875) );
  MX4X1 U3597 ( .A(n3937), .B(n3927), .C(n3932), .D(n3922), .S0(n4645), .S1(
        n4635), .Y(n3938) );
  MX4X1 U3598 ( .A(n1546), .B(n1534), .C(n1541), .D(n1529), .S0(n4637), .S1(
        n4632), .Y(n1547) );
  MX4X1 U3599 ( .A(n1533), .B(n1531), .C(n1532), .D(n1530), .S0(n4588), .S1(
        n4530), .Y(n1534) );
  MX4X1 U3600 ( .A(n1528), .B(n1526), .C(n1527), .D(n1525), .S0(n4588), .S1(
        n4530), .Y(n1529) );
  MX4X1 U3601 ( .A(n1545), .B(n1543), .C(n1544), .D(n1542), .S0(n4588), .S1(
        n4530), .Y(n1546) );
  MX4X1 U3602 ( .A(n1900), .B(n1890), .C(n1895), .D(n1885), .S0(n4638), .S1(
        n4628), .Y(n1901) );
  MX4X1 U3603 ( .A(n1889), .B(n1887), .C(n1888), .D(n1886), .S0(n4593), .S1(
        n4535), .Y(n1890) );
  MX4X1 U3604 ( .A(n1884), .B(n1882), .C(n1883), .D(n1881), .S0(n4593), .S1(
        n4535), .Y(n1885) );
  MX4X1 U3605 ( .A(n1899), .B(n1897), .C(n1898), .D(n1896), .S0(n4593), .S1(
        n4535), .Y(n1900) );
  MX4X1 U3606 ( .A(n1636), .B(n1626), .C(n1631), .D(n1621), .S0(n4637), .S1(
        n4630), .Y(n1637) );
  MX4X1 U3607 ( .A(n1625), .B(n1623), .C(n1624), .D(n1622), .S0(n4589), .S1(
        n4531), .Y(n1626) );
  MX4X1 U3608 ( .A(n1620), .B(n1618), .C(n1619), .D(n1617), .S0(n4589), .S1(
        n4531), .Y(n1621) );
  MX4X1 U3609 ( .A(n1635), .B(n1633), .C(n1634), .D(n1632), .S0(n4589), .S1(
        n4531), .Y(n1636) );
  MX4X1 U3610 ( .A(n1724), .B(n1714), .C(n1719), .D(n1709), .S0(n4638), .S1(
        n4633), .Y(n1725) );
  MX4X1 U3611 ( .A(n1713), .B(n1711), .C(n1712), .D(n1710), .S0(n4591), .S1(
        n4532), .Y(n1714) );
  MX4X1 U3612 ( .A(n1708), .B(n1705), .C(n1706), .D(n1704), .S0(n4591), .S1(
        n4532), .Y(n1709) );
  MX4X1 U3613 ( .A(n1723), .B(n1721), .C(n1722), .D(n1720), .S0(n4591), .S1(
        n4532), .Y(n1724) );
  MX4X1 U3614 ( .A(n2252), .B(n2242), .C(n2247), .D(n2236), .S0(n4640), .S1(
        n4629), .Y(n2253) );
  MX4X1 U3615 ( .A(n2241), .B(n2239), .C(n2240), .D(n2238), .S0(n4599), .S1(
        n4540), .Y(n2242) );
  MX4X1 U3616 ( .A(n2235), .B(n2233), .C(n2234), .D(n2232), .S0(n4599), .S1(
        n4540), .Y(n2236) );
  MX4X1 U3617 ( .A(n2251), .B(n2249), .C(n2250), .D(n2248), .S0(n4599), .S1(
        n4540), .Y(n2252) );
  MX4X1 U3618 ( .A(n1988), .B(n1978), .C(n1983), .D(n1973), .S0(n4639), .S1(
        n4628), .Y(n1989) );
  MX4X1 U3619 ( .A(n1977), .B(n1975), .C(n1976), .D(n1974), .S0(n4595), .S1(
        n4536), .Y(n1978) );
  MX4X1 U3620 ( .A(n1971), .B(n1969), .C(n1970), .D(n1968), .S0(n4595), .S1(
        n4536), .Y(n1973) );
  MX4X1 U3621 ( .A(n1987), .B(n1985), .C(n1986), .D(n1984), .S0(n4595), .S1(
        n4536), .Y(n1988) );
  MX4X1 U3622 ( .A(n2076), .B(n2065), .C(n2070), .D(n2060), .S0(n4639), .S1(
        n4629), .Y(n2077) );
  MX4X1 U3623 ( .A(n2064), .B(n2062), .C(n2063), .D(n2061), .S0(n4596), .S1(
        n4537), .Y(n2065) );
  MX4X1 U3624 ( .A(n2059), .B(n2057), .C(n2058), .D(n2056), .S0(n4596), .S1(
        n4537), .Y(n2060) );
  MX4X1 U3625 ( .A(n2075), .B(n2073), .C(n2074), .D(n2072), .S0(n4596), .S1(
        n4537), .Y(n2076) );
  MX4X1 U3626 ( .A(n2662), .B(n2652), .C(n2657), .D(n2647), .S0(n4641), .S1(
        n4631), .Y(n2663) );
  MX4X1 U3627 ( .A(n2651), .B(n2649), .C(n2650), .D(n2648), .S0(n4604), .S1(
        n4544), .Y(n2652) );
  MX4X1 U3628 ( .A(n2646), .B(n2644), .C(n2645), .D(n2643), .S0(n4604), .S1(
        n4544), .Y(n2647) );
  MX4X1 U3629 ( .A(n2661), .B(n2659), .C(n2660), .D(n2658), .S0(n4604), .S1(
        n4544), .Y(n2662) );
  MX4X1 U3630 ( .A(n2345), .B(n2329), .C(n2334), .D(n2324), .S0(n4640), .S1(
        n4630), .Y(n2347) );
  MX4X1 U3631 ( .A(n2328), .B(n2326), .C(n2327), .D(n2325), .S0(n4600), .S1(
        n4541), .Y(n2329) );
  MX4X1 U3632 ( .A(n2323), .B(n2321), .C(n2322), .D(n2320), .S0(n4600), .S1(
        n4541), .Y(n2324) );
  MX4X1 U3633 ( .A(n2343), .B(n2339), .C(n2341), .D(n2335), .S0(n4600), .S1(
        n4541), .Y(n2345) );
  MX4X1 U3634 ( .A(n2492), .B(n2482), .C(n2487), .D(n2477), .S0(n4640), .S1(
        n4630), .Y(n2493) );
  MX4X1 U3635 ( .A(n2481), .B(n2479), .C(n2480), .D(n2478), .S0(n4601), .S1(
        n4542), .Y(n2482) );
  MX4X1 U3636 ( .A(n2476), .B(n2474), .C(n2475), .D(n2473), .S0(n4601), .S1(
        n4542), .Y(n2477) );
  MX4X1 U3637 ( .A(n2491), .B(n2489), .C(n2490), .D(n2488), .S0(n4601), .S1(
        n4542), .Y(n2492) );
  MX4X1 U3638 ( .A(n3002), .B(n2992), .C(n2997), .D(n2987), .S0(n4642), .S1(
        n4632), .Y(n3003) );
  MX4X1 U3639 ( .A(n2991), .B(n2989), .C(n2990), .D(n2988), .S0(n4609), .S1(
        n4549), .Y(n2992) );
  MX4X1 U3640 ( .A(n2986), .B(n2984), .C(n2985), .D(n2983), .S0(n4609), .S1(
        n4548), .Y(n2987) );
  MX4X1 U3641 ( .A(n3001), .B(n2999), .C(n3000), .D(n2998), .S0(n4609), .S1(
        n4549), .Y(n3002) );
  MX4X1 U3642 ( .A(n2747), .B(n2737), .C(n2742), .D(n2732), .S0(n4641), .S1(
        n4631), .Y(n2748) );
  MX4X1 U3643 ( .A(n2736), .B(n2734), .C(n2735), .D(n2733), .S0(n4605), .S1(
        n4545), .Y(n2737) );
  MX4X1 U3644 ( .A(n2731), .B(n2729), .C(n2730), .D(n2728), .S0(n4605), .S1(
        n4545), .Y(n2732) );
  MX4X1 U3645 ( .A(n2746), .B(n2744), .C(n2745), .D(n2743), .S0(n4605), .S1(
        n4545), .Y(n2747) );
  MX4X1 U3646 ( .A(n2832), .B(n2822), .C(n2827), .D(n2817), .S0(n4642), .S1(
        n4631), .Y(n2833) );
  MX4X1 U3647 ( .A(n2821), .B(n2819), .C(n2820), .D(n2818), .S0(n4607), .S1(
        n4546), .Y(n2822) );
  MX4X1 U3648 ( .A(n2816), .B(n2814), .C(n2815), .D(n2813), .S0(n4607), .S1(
        n4546), .Y(n2817) );
  MX4X1 U3649 ( .A(n2831), .B(n2829), .C(n2830), .D(n2828), .S0(n4607), .S1(
        n4546), .Y(n2832) );
  MX4X1 U3650 ( .A(n3342), .B(n3332), .C(n3337), .D(n3327), .S0(n4644), .S1(
        n4633), .Y(n3343) );
  MX4X1 U3651 ( .A(n3331), .B(n3329), .C(n3330), .D(n3328), .S0(n4615), .S1(
        n4553), .Y(n3332) );
  MX4X1 U3652 ( .A(n3326), .B(n3324), .C(n3325), .D(n3323), .S0(n4615), .S1(
        n4553), .Y(n3327) );
  MX4X1 U3653 ( .A(n3341), .B(n3339), .C(n3340), .D(n3338), .S0(n4615), .S1(
        n4554), .Y(n3342) );
  MX4X1 U3654 ( .A(n3087), .B(n3077), .C(n3082), .D(n3072), .S0(n4643), .S1(
        n4632), .Y(n3088) );
  MX4X1 U3655 ( .A(n3076), .B(n3074), .C(n3075), .D(n3073), .S0(n4611), .S1(
        n4550), .Y(n3077) );
  MX4X1 U3656 ( .A(n3071), .B(n3069), .C(n3070), .D(n3068), .S0(n4611), .S1(
        n4550), .Y(n3072) );
  MX4X1 U3657 ( .A(n3086), .B(n3084), .C(n3085), .D(n3083), .S0(n4611), .S1(
        n4550), .Y(n3087) );
  MX4X1 U3658 ( .A(n3172), .B(n3162), .C(n3167), .D(n3157), .S0(n4643), .S1(
        n4632), .Y(n3173) );
  MX4X1 U3659 ( .A(n3161), .B(n3159), .C(n3160), .D(n3158), .S0(n4612), .S1(
        n4551), .Y(n3162) );
  MX4X1 U3660 ( .A(n3156), .B(n3154), .C(n3155), .D(n3153), .S0(n4612), .S1(
        n4551), .Y(n3157) );
  MX4X1 U3661 ( .A(n3171), .B(n3169), .C(n3170), .D(n3168), .S0(n4612), .S1(
        n4551), .Y(n3172) );
  MX4X1 U3662 ( .A(n3682), .B(n3672), .C(n3677), .D(n3667), .S0(n4641), .S1(
        n4634), .Y(n3683) );
  MX4X1 U3663 ( .A(n3671), .B(n3669), .C(n3670), .D(n3668), .S0(n4620), .S1(
        N70), .Y(n3672) );
  MX4X1 U3664 ( .A(n3666), .B(n3664), .C(n3665), .D(n3663), .S0(n4620), .S1(
        n4508), .Y(n3667) );
  MX4X1 U3665 ( .A(n3681), .B(n3679), .C(n3680), .D(n3678), .S0(n4620), .S1(
        n4531), .Y(n3682) );
  MX4X1 U3666 ( .A(n3427), .B(n3417), .C(n3422), .D(n3412), .S0(n4644), .S1(
        n4633), .Y(n3428) );
  MX4X1 U3667 ( .A(n3416), .B(n3414), .C(n3415), .D(n3413), .S0(n4616), .S1(
        n4555), .Y(n3417) );
  MX4X1 U3668 ( .A(n3411), .B(n3409), .C(n3410), .D(n3408), .S0(n4616), .S1(
        n4555), .Y(n3412) );
  MX4X1 U3669 ( .A(n3426), .B(n3424), .C(n3425), .D(n3423), .S0(n4616), .S1(
        n4555), .Y(n3427) );
  MX4X1 U3670 ( .A(n3512), .B(n3502), .C(n3507), .D(n3497), .S0(n4644), .S1(
        n4634), .Y(n3513) );
  MX4X1 U3671 ( .A(n3501), .B(n3499), .C(n3500), .D(n3498), .S0(n4617), .S1(
        n4556), .Y(n3502) );
  MX4X1 U3672 ( .A(n3496), .B(n3494), .C(n3495), .D(n3493), .S0(n4617), .S1(
        n4556), .Y(n3497) );
  MX4X1 U3673 ( .A(n3511), .B(n3509), .C(n3510), .D(n3508), .S0(n4617), .S1(
        n4556), .Y(n3512) );
  MX4X1 U3674 ( .A(n3767), .B(n3757), .C(n3762), .D(n3752), .S0(n4642), .S1(
        n4635), .Y(n3768) );
  MX4X1 U3675 ( .A(n3756), .B(n3754), .C(n3755), .D(n3753), .S0(n4621), .S1(
        n4545), .Y(n3757) );
  MX4X1 U3676 ( .A(n3751), .B(n3749), .C(n3750), .D(n3748), .S0(n4621), .S1(
        n4558), .Y(n3752) );
  MX4X1 U3677 ( .A(n3766), .B(n3764), .C(n3765), .D(n3763), .S0(n4621), .S1(
        n4542), .Y(n3767) );
  MX4X1 U3678 ( .A(n3852), .B(n3842), .C(n3847), .D(n3837), .S0(n4645), .S1(
        n4635), .Y(n3853) );
  MX4X1 U3679 ( .A(n3841), .B(n3839), .C(n3840), .D(n3838), .S0(n4623), .S1(
        n4533), .Y(n3842) );
  MX4X1 U3680 ( .A(n3836), .B(n3834), .C(n3835), .D(n3833), .S0(n4623), .S1(
        n4537), .Y(n3837) );
  MX4X1 U3681 ( .A(n3851), .B(n3849), .C(n3850), .D(n3848), .S0(n4623), .S1(
        n4544), .Y(n3852) );
  MX4X1 U3682 ( .A(n4987), .B(n4977), .C(n4982), .D(n4972), .S0(n7981), .S1(
        n7972), .Y(n4988) );
  MX4X1 U3683 ( .A(n4976), .B(n4974), .C(n4975), .D(n4973), .S0(n7931), .S1(
        n7871), .Y(n4977) );
  MX4X1 U3684 ( .A(n4971), .B(n4969), .C(n4970), .D(n4968), .S0(n7931), .S1(
        n7871), .Y(n4972) );
  MX4X1 U3685 ( .A(n4986), .B(n4984), .C(n4985), .D(n4983), .S0(n7931), .S1(
        n7871), .Y(n4987) );
  MX4X1 U3686 ( .A(n5327), .B(n5317), .C(n5322), .D(n5312), .S0(n7982), .S1(
        n7973), .Y(n5328) );
  MX4X1 U3687 ( .A(n5316), .B(n5314), .C(n5315), .D(n5313), .S0(n7936), .S1(
        n7876), .Y(n5317) );
  MX4X1 U3688 ( .A(n5311), .B(n5309), .C(n5310), .D(n5308), .S0(n7936), .S1(
        n7876), .Y(n5312) );
  MX4X1 U3689 ( .A(n5326), .B(n5324), .C(n5325), .D(n5323), .S0(n7936), .S1(
        n7876), .Y(n5327) );
  MX4X1 U3690 ( .A(n5072), .B(n5062), .C(n5067), .D(n5057), .S0(n7981), .S1(
        n7972), .Y(n5073) );
  MX4X1 U3691 ( .A(n5061), .B(n5059), .C(n5060), .D(n5058), .S0(n7932), .S1(
        n7872), .Y(n5062) );
  MX4X1 U3692 ( .A(n5056), .B(n5054), .C(n5055), .D(n5053), .S0(n7932), .S1(
        n7872), .Y(n5057) );
  MX4X1 U3693 ( .A(n5071), .B(n5069), .C(n5070), .D(n5068), .S0(n7932), .S1(
        n7872), .Y(n5072) );
  MX4X1 U3694 ( .A(n5157), .B(n5147), .C(n5152), .D(n5142), .S0(n7982), .S1(
        n7972), .Y(n5158) );
  MX4X1 U3695 ( .A(n5146), .B(n5144), .C(n5145), .D(n5143), .S0(n7934), .S1(
        n7873), .Y(n5147) );
  MX4X1 U3696 ( .A(n5141), .B(n5139), .C(n5140), .D(n5138), .S0(n7934), .S1(
        n7873), .Y(n5142) );
  MX4X1 U3697 ( .A(n5156), .B(n5154), .C(n5155), .D(n5153), .S0(n7934), .S1(
        n7873), .Y(n5157) );
  MX4X1 U3698 ( .A(n5667), .B(n5657), .C(n5662), .D(n5652), .S0(n7983), .S1(
        n7974), .Y(n5668) );
  MX4X1 U3699 ( .A(n5656), .B(n5654), .C(n5655), .D(n5653), .S0(n7942), .S1(
        n7881), .Y(n5657) );
  MX4X1 U3700 ( .A(n5651), .B(n5649), .C(n5650), .D(n5648), .S0(n7942), .S1(
        n7881), .Y(n5652) );
  MX4X1 U3701 ( .A(n5666), .B(n5664), .C(n5665), .D(n5663), .S0(n7942), .S1(
        n7881), .Y(n5667) );
  MX4X1 U3702 ( .A(n5412), .B(n5402), .C(n5407), .D(n5397), .S0(n8642), .S1(
        n7973), .Y(n5413) );
  MX4X1 U3703 ( .A(n5401), .B(n5399), .C(n5400), .D(n5398), .S0(n7938), .S1(
        n7877), .Y(n5402) );
  MX4X1 U3704 ( .A(n5396), .B(n5394), .C(n5395), .D(n5393), .S0(n7938), .S1(
        n7877), .Y(n5397) );
  MX4X1 U3705 ( .A(n5411), .B(n5409), .C(n5410), .D(n5408), .S0(n7938), .S1(
        n7877), .Y(n5412) );
  MX4X1 U3706 ( .A(n5497), .B(n5487), .C(n5492), .D(n5482), .S0(n7980), .S1(
        n7974), .Y(n5498) );
  MX4X1 U3707 ( .A(n5486), .B(n5484), .C(n5485), .D(n5483), .S0(n7939), .S1(
        n7878), .Y(n5487) );
  MX4X1 U3708 ( .A(n5481), .B(n5479), .C(n5480), .D(n5478), .S0(n7939), .S1(
        n7878), .Y(n5482) );
  MX4X1 U3709 ( .A(n5496), .B(n5494), .C(n5495), .D(n5493), .S0(n7939), .S1(
        n7878), .Y(n5497) );
  MX4X1 U3710 ( .A(n6007), .B(n5997), .C(n6002), .D(n5992), .S0(n7984), .S1(
        n7976), .Y(n6008) );
  MX4X1 U3711 ( .A(n5996), .B(n5994), .C(n5995), .D(n5993), .S0(n7947), .S1(
        n7886), .Y(n5997) );
  MX4X1 U3712 ( .A(n5991), .B(n5989), .C(n5990), .D(n5988), .S0(n7947), .S1(
        n7886), .Y(n5992) );
  MX4X1 U3713 ( .A(n6006), .B(n6004), .C(n6005), .D(n6003), .S0(n7947), .S1(
        n7886), .Y(n6007) );
  MX4X1 U3714 ( .A(n5752), .B(n5742), .C(n5747), .D(n5737), .S0(n7983), .S1(
        n7975), .Y(n5753) );
  MX4X1 U3715 ( .A(n5741), .B(n5739), .C(n5740), .D(n5738), .S0(n7943), .S1(
        n7882), .Y(n5742) );
  MX4X1 U3716 ( .A(n5736), .B(n5734), .C(n5735), .D(n5733), .S0(n7943), .S1(
        n7882), .Y(n5737) );
  MX4X1 U3717 ( .A(n5751), .B(n5749), .C(n5750), .D(n5748), .S0(n7943), .S1(
        n7882), .Y(n5752) );
  MX4X1 U3718 ( .A(n5837), .B(n5827), .C(n5832), .D(n5822), .S0(n7983), .S1(
        n7975), .Y(n5838) );
  MX4X1 U3719 ( .A(n5826), .B(n5824), .C(n5825), .D(n5823), .S0(n7944), .S1(
        n7883), .Y(n5827) );
  MX4X1 U3720 ( .A(n5821), .B(n5819), .C(n5820), .D(n5818), .S0(n7944), .S1(
        n7883), .Y(n5822) );
  MX4X1 U3721 ( .A(n5836), .B(n5834), .C(n5835), .D(n5833), .S0(n7944), .S1(
        n7883), .Y(n5837) );
  MX4X1 U3722 ( .A(n6347), .B(n6337), .C(n6342), .D(n6332), .S0(n7985), .S1(
        n7977), .Y(n6348) );
  MX4X1 U3723 ( .A(n6336), .B(n6334), .C(n6335), .D(n6333), .S0(n7952), .S1(
        n7891), .Y(n6337) );
  MX4X1 U3724 ( .A(n6331), .B(n6329), .C(n6330), .D(n6328), .S0(n7952), .S1(
        n7890), .Y(n6332) );
  MX4X1 U3725 ( .A(n6346), .B(n6344), .C(n6345), .D(n6343), .S0(n7952), .S1(
        n7891), .Y(n6347) );
  MX4X1 U3726 ( .A(n6092), .B(n6082), .C(n6087), .D(n6077), .S0(n7984), .S1(
        n7976), .Y(n6093) );
  MX4X1 U3727 ( .A(n6081), .B(n6079), .C(n6080), .D(n6078), .S0(n7948), .S1(
        n7887), .Y(n6082) );
  MX4X1 U3728 ( .A(n6076), .B(n6074), .C(n6075), .D(n6073), .S0(n7948), .S1(
        n7887), .Y(n6077) );
  MX4X1 U3729 ( .A(n6091), .B(n6089), .C(n6090), .D(n6088), .S0(n7948), .S1(
        n7887), .Y(n6092) );
  MX4X1 U3730 ( .A(n6177), .B(n6167), .C(n6172), .D(n6162), .S0(n7985), .S1(
        n7976), .Y(n6178) );
  MX4X1 U3731 ( .A(n6166), .B(n6164), .C(n6165), .D(n6163), .S0(n7950), .S1(
        n7888), .Y(n6167) );
  MX4X1 U3732 ( .A(n6161), .B(n6159), .C(n6160), .D(n6158), .S0(n7950), .S1(
        n7888), .Y(n6162) );
  MX4X1 U3733 ( .A(n6176), .B(n6174), .C(n6175), .D(n6173), .S0(n7950), .S1(
        n7888), .Y(n6177) );
  MX4X1 U3734 ( .A(n6687), .B(n6677), .C(n6682), .D(n6672), .S0(n7987), .S1(
        n7972), .Y(n6688) );
  MX4X1 U3735 ( .A(n6676), .B(n6674), .C(n6675), .D(n6673), .S0(n7958), .S1(
        n7895), .Y(n6677) );
  MX4X1 U3736 ( .A(n6671), .B(n6669), .C(n6670), .D(n6668), .S0(n7958), .S1(
        n7895), .Y(n6672) );
  MX4X1 U3737 ( .A(n6686), .B(n6684), .C(n6685), .D(n6683), .S0(n7958), .S1(
        n7896), .Y(n6687) );
  MX4X1 U3738 ( .A(n6432), .B(n6422), .C(n6427), .D(n6417), .S0(n7986), .S1(
        n7977), .Y(n6433) );
  MX4X1 U3739 ( .A(n6421), .B(n6419), .C(n6420), .D(n6418), .S0(n7954), .S1(
        n7892), .Y(n6422) );
  MX4X1 U3740 ( .A(n6416), .B(n6414), .C(n6415), .D(n6413), .S0(n7954), .S1(
        n7892), .Y(n6417) );
  MX4X1 U3741 ( .A(n6431), .B(n6429), .C(n6430), .D(n6428), .S0(n7954), .S1(
        n7892), .Y(n6432) );
  MX4X1 U3742 ( .A(n6517), .B(n6507), .C(n6512), .D(n6502), .S0(n7986), .S1(
        n7977), .Y(n6518) );
  MX4X1 U3743 ( .A(n6506), .B(n6504), .C(n6505), .D(n6503), .S0(n7955), .S1(
        n7893), .Y(n6507) );
  MX4X1 U3744 ( .A(n6501), .B(n6499), .C(n6500), .D(n6498), .S0(n7955), .S1(
        n7893), .Y(n6502) );
  MX4X1 U3745 ( .A(n6516), .B(n6514), .C(n6515), .D(n6513), .S0(n7955), .S1(
        n7893), .Y(n6517) );
  MX4X1 U3746 ( .A(n7027), .B(n7017), .C(n7022), .D(n7012), .S0(n7988), .S1(
        n7971), .Y(n7028) );
  MX4X1 U3747 ( .A(n7016), .B(n7014), .C(n7015), .D(n7013), .S0(n7963), .S1(
        n7898), .Y(n7017) );
  MX4X1 U3748 ( .A(n7011), .B(n7009), .C(n7010), .D(n7008), .S0(n7963), .S1(
        n7898), .Y(n7012) );
  MX4X1 U3749 ( .A(n7026), .B(n7024), .C(n7025), .D(n7023), .S0(n7963), .S1(
        n7899), .Y(n7027) );
  MX4X1 U3750 ( .A(n6772), .B(n6762), .C(n6767), .D(n6757), .S0(n7987), .S1(
        n7971), .Y(n6773) );
  MX4X1 U3751 ( .A(n6761), .B(n6759), .C(n6760), .D(n6758), .S0(n7959), .S1(
        n7890), .Y(n6762) );
  MX4X1 U3752 ( .A(n6756), .B(n6754), .C(n6755), .D(n6753), .S0(n7959), .S1(
        n7868), .Y(n6757) );
  MX4X1 U3753 ( .A(n6771), .B(n6769), .C(n6770), .D(n6768), .S0(n7959), .S1(
        n7900), .Y(n6772) );
  MX4X1 U3754 ( .A(n6857), .B(n6847), .C(n6852), .D(n6842), .S0(n7987), .S1(
        n8644), .Y(n6858) );
  MX4X1 U3755 ( .A(n6846), .B(n6844), .C(n6845), .D(n6843), .S0(n7960), .S1(
        n7894), .Y(n6847) );
  MX4X1 U3756 ( .A(n6841), .B(n6839), .C(n6840), .D(n6838), .S0(n7960), .S1(
        n7895), .Y(n6842) );
  MX4X1 U3757 ( .A(n6856), .B(n6854), .C(n6855), .D(n6853), .S0(n7960), .S1(
        n7891), .Y(n6857) );
  MX4X1 U3758 ( .A(n7367), .B(n7357), .C(n7362), .D(n7352), .S0(n7985), .S1(
        n7971), .Y(n7368) );
  MX4X1 U3759 ( .A(n7356), .B(n7354), .C(n7355), .D(n7353), .S0(N81), .S1(
        n7902), .Y(n7357) );
  MX4X1 U3760 ( .A(n7351), .B(n7349), .C(n7350), .D(n7348), .S0(n7911), .S1(
        n7902), .Y(n7352) );
  MX4X1 U3761 ( .A(n7366), .B(n7364), .C(n7365), .D(n7363), .S0(N81), .S1(
        n7902), .Y(n7367) );
  MX4X1 U3762 ( .A(n7112), .B(n7102), .C(n7107), .D(n7097), .S0(n7988), .S1(
        N82), .Y(n7113) );
  MX4X1 U3763 ( .A(n7101), .B(n7099), .C(n7100), .D(n7098), .S0(n7964), .S1(
        n7900), .Y(n7102) );
  MX4X1 U3764 ( .A(n7096), .B(n7094), .C(n7095), .D(n7093), .S0(n7964), .S1(
        n7900), .Y(n7097) );
  MX4X1 U3765 ( .A(n7111), .B(n7109), .C(n7110), .D(n7108), .S0(n7964), .S1(
        n7900), .Y(n7112) );
  MX4X1 U3766 ( .A(n7197), .B(n7187), .C(n7192), .D(n7182), .S0(n7982), .S1(
        n7971), .Y(n7198) );
  MX4X1 U3767 ( .A(n7186), .B(n7184), .C(n7185), .D(n7183), .S0(n7966), .S1(
        n7901), .Y(n7187) );
  MX4X1 U3768 ( .A(n7181), .B(n7179), .C(n7180), .D(n7178), .S0(n7966), .S1(
        n7901), .Y(n7182) );
  MX4X1 U3769 ( .A(n7196), .B(n7194), .C(n7195), .D(n7193), .S0(n7966), .S1(
        n7901), .Y(n7197) );
  MX4X1 U3770 ( .A(n1479), .B(n1467), .C(n1474), .D(n1462), .S0(n4637), .S1(
        n4628), .Y(n1480) );
  MX4X1 U3771 ( .A(n1466), .B(n1464), .C(n1465), .D(n1463), .S0(n4587), .S1(
        n4529), .Y(n1467) );
  MX4X1 U3772 ( .A(n1461), .B(n1459), .C(n1460), .D(n1458), .S0(n4587), .S1(
        n4529), .Y(n1462) );
  MX4X1 U3773 ( .A(n1478), .B(n1476), .C(n1477), .D(n1475), .S0(n4587), .S1(
        n4529), .Y(n1479) );
  MX4X1 U3774 ( .A(n1834), .B(n1824), .C(n1829), .D(n1819), .S0(n4638), .S1(
        n4628), .Y(n1835) );
  MX4X1 U3775 ( .A(n1823), .B(n1821), .C(n1822), .D(n1820), .S0(n4592), .S1(
        n4534), .Y(n1824) );
  MX4X1 U3776 ( .A(n1818), .B(n1816), .C(n1817), .D(n1815), .S0(n4592), .S1(
        n4534), .Y(n1819) );
  MX4X1 U3777 ( .A(n1833), .B(n1831), .C(n1832), .D(n1830), .S0(n4592), .S1(
        n4534), .Y(n1834) );
  MX4X1 U3778 ( .A(n1568), .B(n1558), .C(n1563), .D(n1553), .S0(n4637), .S1(
        n4629), .Y(n1569) );
  MX4X1 U3779 ( .A(n1557), .B(n1555), .C(n1556), .D(n1554), .S0(n4588), .S1(
        n4530), .Y(n1558) );
  MX4X1 U3780 ( .A(n1552), .B(n1550), .C(n1551), .D(n1549), .S0(n4588), .S1(
        n4530), .Y(n1553) );
  MX4X1 U3781 ( .A(n1567), .B(n1565), .C(n1566), .D(n1564), .S0(n4588), .S1(
        n4530), .Y(n1568) );
  MX4X1 U3782 ( .A(n1659), .B(n1649), .C(n1654), .D(n1644), .S0(n4638), .S1(
        n4630), .Y(n1660) );
  MX4X1 U3783 ( .A(n1648), .B(n1646), .C(n1647), .D(n1645), .S0(n4590), .S1(
        n4531), .Y(n1649) );
  MX4X1 U3784 ( .A(n1643), .B(n1640), .C(n1642), .D(n1639), .S0(n4590), .S1(
        n4531), .Y(n1644) );
  MX4X1 U3785 ( .A(n1658), .B(n1656), .C(n1657), .D(n1655), .S0(n4590), .S1(
        n4532), .Y(n1659) );
  MX4X1 U3786 ( .A(n2187), .B(n2177), .C(n2182), .D(n2172), .S0(n4640), .S1(
        n4629), .Y(n2188) );
  MX4X1 U3787 ( .A(n2176), .B(n2174), .C(n2175), .D(n2173), .S0(n4598), .S1(
        n4539), .Y(n2177) );
  MX4X1 U3788 ( .A(n2170), .B(n2168), .C(n2169), .D(n2167), .S0(n4598), .S1(
        n4539), .Y(n2172) );
  MX4X1 U3789 ( .A(n2186), .B(n2184), .C(n2185), .D(n2183), .S0(n4598), .S1(
        n4539), .Y(n2187) );
  MX4X1 U3790 ( .A(n1923), .B(n1913), .C(n1918), .D(n1908), .S0(n4639), .S1(
        n4628), .Y(n1924) );
  MX4X1 U3791 ( .A(n1912), .B(n1910), .C(n1911), .D(n1909), .S0(n4594), .S1(
        n4535), .Y(n1913) );
  MX4X1 U3792 ( .A(n1907), .B(n1904), .C(n1905), .D(n1903), .S0(n4594), .S1(
        n4535), .Y(n1908) );
  MX4X1 U3793 ( .A(n1922), .B(n1920), .C(n1921), .D(n1919), .S0(n4594), .S1(
        n4535), .Y(n1923) );
  MX4X1 U3794 ( .A(n2011), .B(n2000), .C(n2006), .D(n1995), .S0(n4639), .S1(
        n4628), .Y(n2012) );
  MX4X1 U3795 ( .A(n1999), .B(n1997), .C(n1998), .D(n1996), .S0(n4595), .S1(
        n4536), .Y(n2000) );
  MX4X1 U3796 ( .A(n1994), .B(n1992), .C(n1993), .D(n1991), .S0(n4595), .S1(
        n4536), .Y(n1995) );
  MX4X1 U3797 ( .A(n2010), .B(n2008), .C(n2009), .D(n2007), .S0(n4595), .S1(
        n4536), .Y(n2011) );
  MX4X1 U3798 ( .A(n2599), .B(n2589), .C(n2594), .D(n2584), .S0(n4641), .S1(
        n4630), .Y(n2600) );
  MX4X1 U3799 ( .A(n2588), .B(n2586), .C(n2587), .D(n2585), .S0(n4603), .S1(
        n4538), .Y(n2589) );
  MX4X1 U3800 ( .A(n2583), .B(n2581), .C(n2582), .D(n2580), .S0(n4603), .S1(
        n4543), .Y(n2584) );
  MX4X1 U3801 ( .A(n2598), .B(n2596), .C(n2597), .D(n2595), .S0(n4603), .S1(
        n4544), .Y(n2599) );
  MX4X1 U3802 ( .A(n2275), .B(n2264), .C(n2269), .D(n2259), .S0(n4640), .S1(
        n4629), .Y(n2276) );
  MX4X1 U3803 ( .A(n2263), .B(n2261), .C(n2262), .D(n2260), .S0(n4599), .S1(
        n4540), .Y(n2264) );
  MX4X1 U3804 ( .A(n2258), .B(n2256), .C(n2257), .D(n2255), .S0(n4599), .S1(
        n4540), .Y(n2259) );
  MX4X1 U3805 ( .A(n2274), .B(n2272), .C(n2273), .D(n2271), .S0(n4599), .S1(
        n4540), .Y(n2275) );
  MX4X1 U3806 ( .A(n2374), .B(n2362), .C(n2368), .D(n2357), .S0(n4640), .S1(
        n4630), .Y(n2375) );
  MX4X1 U3807 ( .A(n2361), .B(n2359), .C(n2360), .D(n2358), .S0(n4600), .S1(
        n4541), .Y(n2362) );
  MX4X1 U3808 ( .A(n2356), .B(n2353), .C(n2355), .D(n2351), .S0(n4600), .S1(
        n4541), .Y(n2357) );
  MX4X1 U3809 ( .A(n2373), .B(n2370), .C(n2371), .D(n2369), .S0(n4600), .S1(
        n4541), .Y(n2374) );
  MX4X1 U3810 ( .A(n2939), .B(n2929), .C(n2934), .D(n2924), .S0(n4642), .S1(
        n4632), .Y(n2940) );
  MX4X1 U3811 ( .A(n2928), .B(n2926), .C(n2927), .D(n2925), .S0(n4608), .S1(
        n4548), .Y(n2929) );
  MX4X1 U3812 ( .A(n2923), .B(n2921), .C(n2922), .D(n2920), .S0(n4608), .S1(
        n4548), .Y(n2924) );
  MX4X1 U3813 ( .A(n2938), .B(n2936), .C(n2937), .D(n2935), .S0(n4608), .S1(
        n4548), .Y(n2939) );
  MX4X1 U3814 ( .A(n2684), .B(n2674), .C(n2679), .D(n2669), .S0(n4641), .S1(
        n4631), .Y(n2685) );
  MX4X1 U3815 ( .A(n2673), .B(n2671), .C(n2672), .D(n2670), .S0(n4604), .S1(
        n4544), .Y(n2674) );
  MX4X1 U3816 ( .A(n2668), .B(n2666), .C(n2667), .D(n2665), .S0(n4604), .S1(
        n4544), .Y(n2669) );
  MX4X1 U3817 ( .A(n2683), .B(n2681), .C(n2682), .D(n2680), .S0(n4604), .S1(
        n4544), .Y(n2684) );
  MX4X1 U3818 ( .A(n2769), .B(n2759), .C(n2764), .D(n2754), .S0(n4642), .S1(
        n4631), .Y(n2770) );
  MX4X1 U3819 ( .A(n2758), .B(n2756), .C(n2757), .D(n2755), .S0(n4606), .S1(
        n4545), .Y(n2759) );
  MX4X1 U3820 ( .A(n2753), .B(n2751), .C(n2752), .D(n2750), .S0(n4606), .S1(
        n4545), .Y(n2754) );
  MX4X1 U3821 ( .A(n2768), .B(n2766), .C(n2767), .D(n2765), .S0(n4606), .S1(
        n4545), .Y(n2769) );
  MX4X1 U3822 ( .A(n3279), .B(n3269), .C(n3274), .D(n3264), .S0(n4644), .S1(
        n4633), .Y(n3280) );
  MX4X1 U3823 ( .A(n3268), .B(n3266), .C(n3267), .D(n3265), .S0(n4614), .S1(
        n4553), .Y(n3269) );
  MX4X1 U3824 ( .A(n3263), .B(n3261), .C(n3262), .D(n3260), .S0(n4614), .S1(
        n4552), .Y(n3264) );
  MX4X1 U3825 ( .A(n3278), .B(n3276), .C(n3277), .D(n3275), .S0(n4614), .S1(
        n4553), .Y(n3279) );
  MX4X1 U3826 ( .A(n3024), .B(n3014), .C(n3019), .D(n3009), .S0(n4643), .S1(
        n4632), .Y(n3025) );
  MX4X1 U3827 ( .A(n3013), .B(n3011), .C(n3012), .D(n3010), .S0(n4610), .S1(
        n4549), .Y(n3014) );
  MX4X1 U3828 ( .A(n3008), .B(n3006), .C(n3007), .D(n3005), .S0(n4610), .S1(
        n4549), .Y(n3009) );
  MX4X1 U3829 ( .A(n3023), .B(n3021), .C(n3022), .D(n3020), .S0(n4610), .S1(
        n4549), .Y(n3024) );
  MX4X1 U3830 ( .A(n3109), .B(n3099), .C(n3104), .D(n3094), .S0(n4643), .S1(
        n4632), .Y(n3110) );
  MX4X1 U3831 ( .A(n3098), .B(n3096), .C(n3097), .D(n3095), .S0(n4611), .S1(
        n4550), .Y(n3099) );
  MX4X1 U3832 ( .A(n3093), .B(n3091), .C(n3092), .D(n3090), .S0(n4611), .S1(
        n4550), .Y(n3094) );
  MX4X1 U3833 ( .A(n3108), .B(n3106), .C(n3107), .D(n3105), .S0(n4611), .S1(
        n4550), .Y(n3109) );
  MX4X1 U3834 ( .A(n3619), .B(n3609), .C(n3614), .D(n3604), .S0(n4638), .S1(
        n4634), .Y(n3620) );
  MX4X1 U3835 ( .A(n3608), .B(n3606), .C(n3607), .D(n3605), .S0(n4619), .S1(
        n4557), .Y(n3609) );
  MX4X1 U3836 ( .A(n3603), .B(n3601), .C(n3602), .D(n3600), .S0(n4619), .S1(
        n4557), .Y(n3604) );
  MX4X1 U3837 ( .A(n3618), .B(n3616), .C(n3617), .D(n3615), .S0(n4619), .S1(
        n4509), .Y(n3619) );
  MX4X1 U3838 ( .A(n3364), .B(n3354), .C(n3359), .D(n3349), .S0(n4644), .S1(
        n4633), .Y(n3365) );
  MX4X1 U3839 ( .A(n3353), .B(n3351), .C(n3352), .D(n3350), .S0(n4615), .S1(
        n4554), .Y(n3354) );
  MX4X1 U3840 ( .A(n3348), .B(n3346), .C(n3347), .D(n3345), .S0(n4615), .S1(
        n4554), .Y(n3349) );
  MX4X1 U3841 ( .A(n3363), .B(n3361), .C(n3362), .D(n3360), .S0(n4615), .S1(
        n4554), .Y(n3364) );
  MX4X1 U3842 ( .A(n3449), .B(n3439), .C(n3444), .D(n3434), .S0(n4644), .S1(
        n4633), .Y(n3450) );
  MX4X1 U3843 ( .A(n3438), .B(n3436), .C(n3437), .D(n3435), .S0(n4616), .S1(
        n4555), .Y(n3439) );
  MX4X1 U3844 ( .A(n3433), .B(n3431), .C(n3432), .D(n3430), .S0(n4616), .S1(
        n4555), .Y(n3434) );
  MX4X1 U3845 ( .A(n3448), .B(n3446), .C(n3447), .D(n3445), .S0(n4616), .S1(
        n4555), .Y(n3449) );
  MX4X1 U3846 ( .A(n4022), .B(n4012), .C(n4017), .D(n4007), .S0(n4645), .S1(
        n4635), .Y(n4023) );
  MX4X1 U3847 ( .A(n4011), .B(n4009), .C(n4010), .D(n4008), .S0(N71), .S1(
        n4559), .Y(n4012) );
  MX4X1 U3848 ( .A(n4006), .B(n4004), .C(n4005), .D(n4003), .S0(n4569), .S1(
        n4559), .Y(n4007) );
  MX4X1 U3849 ( .A(n4021), .B(n4019), .C(n4020), .D(n4018), .S0(N71), .S1(
        n4559), .Y(n4022) );
  MX4X1 U3850 ( .A(n3959), .B(n3949), .C(n3954), .D(n3944), .S0(n4645), .S1(
        n4635), .Y(n3960) );
  MX4X1 U3851 ( .A(n3948), .B(n3946), .C(n3947), .D(n3945), .S0(n4624), .S1(
        n4558), .Y(n3949) );
  MX4X1 U3852 ( .A(n3943), .B(n3941), .C(n3942), .D(n3940), .S0(n4624), .S1(
        n4558), .Y(n3944) );
  MX4X1 U3853 ( .A(n3958), .B(n3956), .C(n3957), .D(n3955), .S0(n4624), .S1(
        n4559), .Y(n3959) );
  MX4X1 U3854 ( .A(n3704), .B(n3694), .C(n3699), .D(n3689), .S0(n4644), .S1(
        n4634), .Y(n3705) );
  MX4X1 U3855 ( .A(n3693), .B(n3691), .C(n3692), .D(n3690), .S0(n4620), .S1(
        n4558), .Y(n3694) );
  MX4X1 U3856 ( .A(n3688), .B(n3686), .C(n3687), .D(n3685), .S0(n4620), .S1(
        n4535), .Y(n3689) );
  MX4X1 U3857 ( .A(n3703), .B(n3701), .C(n3702), .D(n3700), .S0(n4620), .S1(
        n4530), .Y(n3704) );
  MX4X1 U3858 ( .A(n3789), .B(n3779), .C(n3784), .D(n3774), .S0(n4645), .S1(
        n4635), .Y(n3790) );
  MX4X1 U3859 ( .A(n3778), .B(n3776), .C(n3777), .D(n3775), .S0(n4622), .S1(
        n4526), .Y(n3779) );
  MX4X1 U3860 ( .A(n3773), .B(n3771), .C(n3772), .D(n3770), .S0(n4622), .S1(
        n4538), .Y(n3774) );
  MX4X1 U3861 ( .A(n3788), .B(n3786), .C(n3787), .D(n3785), .S0(n4622), .S1(
        n4531), .Y(n3789) );
  MX4X1 U3862 ( .A(n4924), .B(n4914), .C(n4919), .D(n4909), .S0(n7981), .S1(
        n7972), .Y(n4925) );
  MX4X1 U3863 ( .A(n4913), .B(n4911), .C(n4912), .D(n4910), .S0(n7930), .S1(
        n7870), .Y(n4914) );
  MX4X1 U3864 ( .A(n4908), .B(n4906), .C(n4907), .D(n4905), .S0(n7930), .S1(
        n7870), .Y(n4909) );
  MX4X1 U3865 ( .A(n4923), .B(n4921), .C(n4922), .D(n4920), .S0(n7930), .S1(
        n7870), .Y(n4924) );
  MX4X1 U3866 ( .A(n4754), .B(n4744), .C(n4749), .D(n4739), .S0(n8642), .S1(
        n7971), .Y(n4755) );
  MX4X1 U3867 ( .A(n4743), .B(n4741), .C(n4742), .D(n4740), .S0(n7933), .S1(
        n7867), .Y(n4744) );
  MX4X1 U3868 ( .A(n4738), .B(n4736), .C(n4737), .D(n4735), .S0(n7930), .S1(
        n7867), .Y(n4739) );
  MX4X1 U3869 ( .A(n4753), .B(n4751), .C(n4752), .D(n4750), .S0(n7951), .S1(
        n7868), .Y(n4754) );
  MX4X1 U3870 ( .A(n5264), .B(n5254), .C(n5259), .D(n5249), .S0(n7982), .S1(
        n7973), .Y(n5265) );
  MX4X1 U3871 ( .A(n5253), .B(n5251), .C(n5252), .D(n5250), .S0(n7935), .S1(
        n7875), .Y(n5254) );
  MX4X1 U3872 ( .A(n5248), .B(n5246), .C(n5247), .D(n5245), .S0(n7935), .S1(
        n7875), .Y(n5249) );
  MX4X1 U3873 ( .A(n5263), .B(n5261), .C(n5262), .D(n5260), .S0(n7935), .S1(
        n7875), .Y(n5264) );
  MX4X1 U3874 ( .A(n5009), .B(n4999), .C(n5004), .D(n4994), .S0(n7981), .S1(
        n7972), .Y(n5010) );
  MX4X1 U3875 ( .A(n4998), .B(n4996), .C(n4997), .D(n4995), .S0(n7931), .S1(
        n7871), .Y(n4999) );
  MX4X1 U3876 ( .A(n4993), .B(n4991), .C(n4992), .D(n4990), .S0(n7931), .S1(
        n7871), .Y(n4994) );
  MX4X1 U3877 ( .A(n5008), .B(n5006), .C(n5007), .D(n5005), .S0(n7931), .S1(
        n7871), .Y(n5009) );
  MX4X1 U3878 ( .A(n5094), .B(n5084), .C(n5089), .D(n5079), .S0(n7982), .S1(
        n7972), .Y(n5095) );
  MX4X1 U3879 ( .A(n5083), .B(n5081), .C(n5082), .D(n5080), .S0(n7933), .S1(
        n7872), .Y(n5084) );
  MX4X1 U3880 ( .A(n5078), .B(n5076), .C(n5077), .D(n5075), .S0(n7933), .S1(
        n7872), .Y(n5079) );
  MX4X1 U3881 ( .A(n5093), .B(n5091), .C(n5092), .D(n5090), .S0(n7933), .S1(
        n7873), .Y(n5094) );
  MX4X1 U3882 ( .A(n5604), .B(n5594), .C(n5599), .D(n5589), .S0(n7983), .S1(
        n7974), .Y(n5605) );
  MX4X1 U3883 ( .A(n5593), .B(n5591), .C(n5592), .D(n5590), .S0(n7941), .S1(
        n7880), .Y(n5594) );
  MX4X1 U3884 ( .A(n5588), .B(n5586), .C(n5587), .D(n5585), .S0(n7941), .S1(
        n7880), .Y(n5589) );
  MX4X1 U3885 ( .A(n5603), .B(n5601), .C(n5602), .D(n5600), .S0(n7941), .S1(
        n7880), .Y(n5604) );
  MX4X1 U3886 ( .A(n5349), .B(n5339), .C(n5344), .D(n5334), .S0(n7982), .S1(
        n7973), .Y(n5350) );
  MX4X1 U3887 ( .A(n5338), .B(n5336), .C(n5337), .D(n5335), .S0(n7937), .S1(
        n7876), .Y(n5339) );
  MX4X1 U3888 ( .A(n5333), .B(n5331), .C(n5332), .D(n5330), .S0(n7937), .S1(
        n7876), .Y(n5334) );
  MX4X1 U3889 ( .A(n5348), .B(n5346), .C(n5347), .D(n5345), .S0(n7937), .S1(
        n7876), .Y(n5349) );
  MX4X1 U3890 ( .A(n5434), .B(n5424), .C(n5429), .D(n5419), .S0(n7988), .S1(
        n7973), .Y(n5435) );
  MX4X1 U3891 ( .A(n5423), .B(n5421), .C(n5422), .D(n5420), .S0(n7938), .S1(
        n7877), .Y(n5424) );
  MX4X1 U3892 ( .A(n5418), .B(n5416), .C(n5417), .D(n5415), .S0(n7938), .S1(
        n7877), .Y(n5419) );
  MX4X1 U3893 ( .A(n5433), .B(n5431), .C(n5432), .D(n5430), .S0(n7938), .S1(
        n7877), .Y(n5434) );
  MX4X1 U3894 ( .A(n5944), .B(n5934), .C(n5939), .D(n5929), .S0(n7984), .S1(
        n7975), .Y(n5945) );
  MX4X1 U3895 ( .A(n5933), .B(n5931), .C(n5932), .D(n5930), .S0(n7946), .S1(
        n7885), .Y(n5934) );
  MX4X1 U3896 ( .A(n5928), .B(n5926), .C(n5927), .D(n5925), .S0(n7946), .S1(
        n7885), .Y(n5929) );
  MX4X1 U3897 ( .A(n5943), .B(n5941), .C(n5942), .D(n5940), .S0(n7946), .S1(
        n7885), .Y(n5944) );
  MX4X1 U3898 ( .A(n5689), .B(n5679), .C(n5684), .D(n5674), .S0(n7983), .S1(
        n7974), .Y(n5690) );
  MX4X1 U3899 ( .A(n5678), .B(n5676), .C(n5677), .D(n5675), .S0(n7942), .S1(
        n7881), .Y(n5679) );
  MX4X1 U3900 ( .A(n5673), .B(n5671), .C(n5672), .D(n5670), .S0(n7942), .S1(
        n7881), .Y(n5674) );
  MX4X1 U3901 ( .A(n5688), .B(n5686), .C(n5687), .D(n5685), .S0(n7942), .S1(
        n7881), .Y(n5689) );
  MX4X1 U3902 ( .A(n5774), .B(n5764), .C(n5769), .D(n5759), .S0(n7983), .S1(
        n7975), .Y(n5775) );
  MX4X1 U3903 ( .A(n5763), .B(n5761), .C(n5762), .D(n5760), .S0(n7943), .S1(
        n7882), .Y(n5764) );
  MX4X1 U3904 ( .A(n5758), .B(n5756), .C(n5757), .D(n5755), .S0(n7943), .S1(
        n7882), .Y(n5759) );
  MX4X1 U3905 ( .A(n5773), .B(n5771), .C(n5772), .D(n5770), .S0(n7943), .S1(
        n7882), .Y(n5774) );
  MX4X1 U3906 ( .A(n6284), .B(n6274), .C(n6279), .D(n6269), .S0(n7985), .S1(
        n7977), .Y(n6285) );
  MX4X1 U3907 ( .A(n6273), .B(n6271), .C(n6272), .D(n6270), .S0(n7951), .S1(
        n7890), .Y(n6274) );
  MX4X1 U3908 ( .A(n6268), .B(n6266), .C(n6267), .D(n6265), .S0(n7951), .S1(
        n7890), .Y(n6269) );
  MX4X1 U3909 ( .A(n6283), .B(n6281), .C(n6282), .D(n6280), .S0(n7951), .S1(
        n7890), .Y(n6284) );
  MX4X1 U3910 ( .A(n6029), .B(n6019), .C(n6024), .D(n6014), .S0(n7984), .S1(
        n7976), .Y(n6030) );
  MX4X1 U3911 ( .A(n6018), .B(n6016), .C(n6017), .D(n6015), .S0(n7947), .S1(
        n7886), .Y(n6019) );
  MX4X1 U3912 ( .A(n6013), .B(n6011), .C(n6012), .D(n6010), .S0(n7947), .S1(
        n7886), .Y(n6014) );
  MX4X1 U3913 ( .A(n6028), .B(n6026), .C(n6027), .D(n6025), .S0(n7947), .S1(
        n7886), .Y(n6029) );
  MX4X1 U3914 ( .A(n6114), .B(n6104), .C(n6109), .D(n6099), .S0(n7985), .S1(
        n7976), .Y(n6115) );
  MX4X1 U3915 ( .A(n6103), .B(n6101), .C(n6102), .D(n6100), .S0(n7949), .S1(
        n7887), .Y(n6104) );
  MX4X1 U3916 ( .A(n6098), .B(n6096), .C(n6097), .D(n6095), .S0(n7949), .S1(
        n7887), .Y(n6099) );
  MX4X1 U3917 ( .A(n6113), .B(n6111), .C(n6112), .D(n6110), .S0(n7949), .S1(
        n7887), .Y(n6114) );
  MX4X1 U3918 ( .A(n6624), .B(n6614), .C(n6619), .D(n6609), .S0(n7987), .S1(
        n7978), .Y(n6625) );
  MX4X1 U3919 ( .A(n6613), .B(n6611), .C(n6612), .D(n6610), .S0(n7957), .S1(
        n7895), .Y(n6614) );
  MX4X1 U3920 ( .A(n6608), .B(n6606), .C(n6607), .D(n6605), .S0(n7957), .S1(
        n7894), .Y(n6609) );
  MX4X1 U3921 ( .A(n6623), .B(n6621), .C(n6622), .D(n6620), .S0(n7957), .S1(
        n7895), .Y(n6624) );
  MX4X1 U3922 ( .A(n6369), .B(n6359), .C(n6364), .D(n6354), .S0(n7986), .S1(
        n7977), .Y(n6370) );
  MX4X1 U3923 ( .A(n6358), .B(n6356), .C(n6357), .D(n6355), .S0(n7953), .S1(
        n7891), .Y(n6359) );
  MX4X1 U3924 ( .A(n6353), .B(n6351), .C(n6352), .D(n6350), .S0(n7953), .S1(
        n7891), .Y(n6354) );
  MX4X1 U3925 ( .A(n6368), .B(n6366), .C(n6367), .D(n6365), .S0(n7953), .S1(
        n7891), .Y(n6369) );
  MX4X1 U3926 ( .A(n6454), .B(n6444), .C(n6449), .D(n6439), .S0(n7986), .S1(
        n7977), .Y(n6455) );
  MX4X1 U3927 ( .A(n6443), .B(n6441), .C(n6442), .D(n6440), .S0(n7954), .S1(
        n7892), .Y(n6444) );
  MX4X1 U3928 ( .A(n6438), .B(n6436), .C(n6437), .D(n6435), .S0(n7954), .S1(
        n7892), .Y(n6439) );
  MX4X1 U3929 ( .A(n6453), .B(n6451), .C(n6452), .D(n6450), .S0(n7954), .S1(
        n7892), .Y(n6454) );
  MX4X1 U3930 ( .A(n6964), .B(n6954), .C(n6959), .D(n6949), .S0(n7988), .S1(
        N82), .Y(n6965) );
  MX4X1 U3931 ( .A(n6953), .B(n6951), .C(n6952), .D(n6950), .S0(n7962), .S1(
        n7897), .Y(n6954) );
  MX4X1 U3932 ( .A(n6948), .B(n6946), .C(n6947), .D(n6945), .S0(n7962), .S1(
        n7897), .Y(n6949) );
  MX4X1 U3933 ( .A(n6963), .B(n6961), .C(n6962), .D(n6960), .S0(n7962), .S1(
        n7898), .Y(n6964) );
  MX4X1 U3934 ( .A(n6709), .B(n6699), .C(n6704), .D(n6694), .S0(n7987), .S1(
        n7976), .Y(n6710) );
  MX4X1 U3935 ( .A(n6698), .B(n6696), .C(n6697), .D(n6695), .S0(n7958), .S1(
        n7896), .Y(n6699) );
  MX4X1 U3936 ( .A(n6693), .B(n6691), .C(n6692), .D(n6690), .S0(n7958), .S1(
        n7896), .Y(n6694) );
  MX4X1 U3937 ( .A(n6708), .B(n6706), .C(n6707), .D(n6705), .S0(n7958), .S1(
        n7896), .Y(n6709) );
  MX4X1 U3938 ( .A(n6794), .B(n6784), .C(n6789), .D(n6779), .S0(n7987), .S1(
        n7976), .Y(n6795) );
  MX4X1 U3939 ( .A(n6783), .B(n6781), .C(n6782), .D(n6780), .S0(n7959), .S1(
        n7895), .Y(n6784) );
  MX4X1 U3940 ( .A(n6778), .B(n6776), .C(n6777), .D(n6775), .S0(n7959), .S1(
        n7893), .Y(n6779) );
  MX4X1 U3941 ( .A(n6793), .B(n6791), .C(n6792), .D(n6790), .S0(n7959), .S1(
        n7898), .Y(n6794) );
  MX4X1 U3942 ( .A(n7304), .B(n7294), .C(n7299), .D(n7289), .S0(N83), .S1(
        n7977), .Y(n7305) );
  MX4X1 U3943 ( .A(n7293), .B(n7291), .C(n7292), .D(n7290), .S0(n7967), .S1(
        n7897), .Y(n7294) );
  MX4X1 U3944 ( .A(n7288), .B(n7286), .C(n7287), .D(n7285), .S0(n7967), .S1(
        n7894), .Y(n7289) );
  MX4X1 U3945 ( .A(n7303), .B(n7301), .C(n7302), .D(n7300), .S0(n7967), .S1(
        n7902), .Y(n7304) );
  MX4X1 U3946 ( .A(n7049), .B(n7039), .C(n7044), .D(n7034), .S0(n7988), .S1(
        N82), .Y(n7050) );
  MX4X1 U3947 ( .A(n7038), .B(n7036), .C(n7037), .D(n7035), .S0(n7963), .S1(
        n7899), .Y(n7039) );
  MX4X1 U3948 ( .A(n7033), .B(n7031), .C(n7032), .D(n7030), .S0(n7963), .S1(
        n7899), .Y(n7034) );
  MX4X1 U3949 ( .A(n7048), .B(n7046), .C(n7047), .D(n7045), .S0(n7963), .S1(
        n7899), .Y(n7049) );
  MX4X1 U3950 ( .A(n7134), .B(n7124), .C(n7129), .D(n7119), .S0(N83), .S1(
        n7977), .Y(n7135) );
  MX4X1 U3951 ( .A(n7123), .B(n7121), .C(n7122), .D(n7120), .S0(n7965), .S1(
        n7900), .Y(n7124) );
  MX4X1 U3952 ( .A(n7118), .B(n7116), .C(n7117), .D(n7115), .S0(n7965), .S1(
        n7900), .Y(n7119) );
  MX4X1 U3953 ( .A(n7133), .B(n7131), .C(n7132), .D(n7130), .S0(n7965), .S1(
        n7900), .Y(n7134) );
  MX4X1 U3954 ( .A(n1813), .B(n1769), .C(n1791), .D(n1748), .S0(n4648), .S1(
        N74), .Y(n1814) );
  MX4X1 U3955 ( .A(n1768), .B(n1758), .C(n1763), .D(n1753), .S0(n4638), .S1(
        n4628), .Y(n1769) );
  MX4X1 U3956 ( .A(n1747), .B(n1736), .C(n1742), .D(n1731), .S0(n4638), .S1(
        n4628), .Y(n1748) );
  MX4X1 U3957 ( .A(n1812), .B(n1801), .C(n1807), .D(n1796), .S0(n4638), .S1(
        n4628), .Y(n1813) );
  MX4X1 U3958 ( .A(n1106), .B(n1096), .C(n1101), .D(n1091), .S0(n4645), .S1(
        n4632), .Y(n1107) );
  MX4X1 U3959 ( .A(n1095), .B(n1093), .C(n1094), .D(n1092), .S0(n4593), .S1(
        n4526), .Y(n1096) );
  MX4X1 U3960 ( .A(n1090), .B(n1088), .C(n1089), .D(n1087), .S0(n4592), .S1(
        n4526), .Y(n1091) );
  MX4X1 U3961 ( .A(n1105), .B(n1103), .C(n1104), .D(n1102), .S0(n4589), .S1(
        n4526), .Y(n1106) );
  MX4X1 U3962 ( .A(n1342), .B(n1329), .C(n1337), .D(n1319), .S0(N73), .S1(
        n4634), .Y(n1343) );
  MX4X1 U3963 ( .A(n1327), .B(n1323), .C(n1325), .D(n1321), .S0(n4602), .S1(
        n4527), .Y(n1329) );
  MX4X1 U3964 ( .A(n1317), .B(n1313), .C(n1315), .D(n1311), .S0(n4600), .S1(
        n4527), .Y(n1319) );
  MX4X1 U3965 ( .A(n1341), .B(n1339), .C(n1340), .D(n1338), .S0(n4595), .S1(
        n4527), .Y(n1342) );
  MX4X1 U3966 ( .A(n4711), .B(n4701), .C(n4706), .D(n4696), .S0(n7980), .S1(
        n7971), .Y(n4712) );
  MX4X1 U3967 ( .A(n4700), .B(n4698), .C(n4699), .D(n4697), .S0(n7936), .S1(
        n7867), .Y(n4701) );
  MX4X1 U3968 ( .A(n4695), .B(n4693), .C(n4694), .D(n4692), .S0(n7935), .S1(
        n7867), .Y(n4696) );
  MX4X1 U3969 ( .A(n4710), .B(n4708), .C(n4709), .D(n4707), .S0(n7932), .S1(
        n7867), .Y(n4711) );
  MX4X1 U3970 ( .A(n4796), .B(n4786), .C(n4791), .D(n4781), .S0(N83), .S1(
        n7971), .Y(n4797) );
  MX4X1 U3971 ( .A(n4785), .B(n4783), .C(n4784), .D(n4782), .S0(n7945), .S1(
        n7868), .Y(n4786) );
  MX4X1 U3972 ( .A(n4780), .B(n4778), .C(n4779), .D(n4777), .S0(n7943), .S1(
        n7868), .Y(n4781) );
  MX4X1 U3973 ( .A(n4795), .B(n4793), .C(n4794), .D(n4792), .S0(n7938), .S1(
        n7868), .Y(n4796) );
  MX4X1 U3974 ( .A(n1456), .B(n1412), .C(n1433), .D(n1389), .S0(n4648), .S1(
        n4646), .Y(n1457) );
  MX4X1 U3975 ( .A(n1411), .B(n1399), .C(n1406), .D(n1394), .S0(n4637), .S1(
        n4632), .Y(n1412) );
  MX4X1 U3976 ( .A(n1388), .B(n1378), .C(n1383), .D(n1373), .S0(n4637), .S1(
        n4633), .Y(n1389) );
  MX4X1 U3977 ( .A(n1455), .B(n1445), .C(n1450), .D(n1440), .S0(n4637), .S1(
        n4629), .Y(n1456) );
  MX4X1 U3978 ( .A(n1169), .B(n1159), .C(n1164), .D(n1154), .S0(N73), .S1(
        n4633), .Y(n1170) );
  MX4X1 U3979 ( .A(n1158), .B(n1156), .C(n1157), .D(n1155), .S0(n4593), .S1(
        n4526), .Y(n1159) );
  MX4X1 U3980 ( .A(n1153), .B(n1151), .C(n1152), .D(n1150), .S0(n4594), .S1(
        n4526), .Y(n1154) );
  MX4X1 U3981 ( .A(n1168), .B(n1166), .C(n1167), .D(n1165), .S0(n4613), .S1(
        n4526), .Y(n1169) );
  MX4X1 U3982 ( .A(n1363), .B(n1353), .C(n1358), .D(n1348), .S0(N73), .S1(
        n4635), .Y(n1364) );
  MX4X1 U3983 ( .A(n1352), .B(n1350), .C(n1351), .D(n1349), .S0(n4598), .S1(
        n4527), .Y(n1353) );
  MX4X1 U3984 ( .A(n1347), .B(n1345), .C(n1346), .D(n1344), .S0(n4597), .S1(
        n4527), .Y(n1348) );
  MX4X1 U3985 ( .A(n1362), .B(n1360), .C(n1361), .D(n1359), .S0(n4617), .S1(
        n4528), .Y(n1363) );
  MX4X1 U3986 ( .A(n4732), .B(n4722), .C(n4727), .D(n4717), .S0(N83), .S1(
        n7971), .Y(n4733) );
  MX4X1 U3987 ( .A(n4721), .B(n4719), .C(n4720), .D(n4718), .S0(n7936), .S1(
        n7867), .Y(n4722) );
  MX4X1 U3988 ( .A(n4716), .B(n4714), .C(n4715), .D(n4713), .S0(n7937), .S1(
        n7867), .Y(n4717) );
  MX4X1 U3989 ( .A(n4731), .B(n4729), .C(n4730), .D(n4728), .S0(n7956), .S1(
        n7867), .Y(n4732) );
  MX4X1 U3990 ( .A(n4817), .B(n4807), .C(n4812), .D(n4802), .S0(N83), .S1(
        n7971), .Y(n4818) );
  MX4X1 U3991 ( .A(n4806), .B(n4804), .C(n4805), .D(n4803), .S0(n7941), .S1(
        n7868), .Y(n4807) );
  MX4X1 U3992 ( .A(n4801), .B(n4799), .C(n4800), .D(n4798), .S0(n7940), .S1(
        n7868), .Y(n4802) );
  MX4X1 U3993 ( .A(n4816), .B(n4814), .C(n4815), .D(n4813), .S0(n7960), .S1(
        n7869), .Y(n4817) );
  MX4X1 U3994 ( .A(n1500), .B(n1490), .C(n1495), .D(n1485), .S0(n4637), .S1(
        N72), .Y(n1501) );
  MX4X1 U3995 ( .A(n1489), .B(n1487), .C(n1488), .D(n1486), .S0(n4587), .S1(
        n4529), .Y(n1490) );
  MX4X1 U3996 ( .A(n1484), .B(n1482), .C(n1483), .D(n1481), .S0(n4587), .S1(
        n4529), .Y(n1485) );
  MX4X1 U3997 ( .A(n1499), .B(n1497), .C(n1498), .D(n1496), .S0(n4587), .S1(
        n4529), .Y(n1500) );
  MX4X1 U3998 ( .A(n1856), .B(n1846), .C(n1851), .D(n1841), .S0(n4638), .S1(
        n4628), .Y(n1857) );
  MX4X1 U3999 ( .A(n1845), .B(n1843), .C(n1844), .D(n1842), .S0(n4593), .S1(
        n4534), .Y(n1846) );
  MX4X1 U4000 ( .A(n1840), .B(n1837), .C(n1838), .D(n1836), .S0(n4593), .S1(
        n4534), .Y(n1841) );
  MX4X1 U4001 ( .A(n1855), .B(n1853), .C(n1854), .D(n1852), .S0(n4593), .S1(
        n4534), .Y(n1856) );
  MX4X1 U4002 ( .A(n1591), .B(n1581), .C(n1586), .D(n1576), .S0(n4637), .S1(
        N72), .Y(n1592) );
  MX4X1 U4003 ( .A(n1580), .B(n1578), .C(n1579), .D(n1577), .S0(n4589), .S1(
        n4530), .Y(n1581) );
  MX4X1 U4004 ( .A(n1575), .B(n1572), .C(n1574), .D(n1570), .S0(n4589), .S1(
        n4530), .Y(n1576) );
  MX4X1 U4005 ( .A(n1590), .B(n1588), .C(n1589), .D(n1587), .S0(n4589), .S1(
        n4531), .Y(n1591) );
  MX4X1 U4006 ( .A(n1681), .B(n1670), .C(n1676), .D(n1665), .S0(n4638), .S1(
        N72), .Y(n1682) );
  MX4X1 U4007 ( .A(n1669), .B(n1667), .C(n1668), .D(n1666), .S0(n4590), .S1(
        n4532), .Y(n1670) );
  MX4X1 U4008 ( .A(n1664), .B(n1662), .C(n1663), .D(n1661), .S0(n4590), .S1(
        n4532), .Y(n1665) );
  MX4X1 U4009 ( .A(n1680), .B(n1678), .C(n1679), .D(n1677), .S0(n4590), .S1(
        n4532), .Y(n1681) );
  MX4X1 U4010 ( .A(n2209), .B(n2198), .C(n2203), .D(n2193), .S0(n4640), .S1(
        n4629), .Y(n2210) );
  MX4X1 U4011 ( .A(n2197), .B(n2195), .C(n2196), .D(n2194), .S0(n4598), .S1(
        n4539), .Y(n2198) );
  MX4X1 U4012 ( .A(n2192), .B(n2190), .C(n2191), .D(n2189), .S0(n4598), .S1(
        n4539), .Y(n2193) );
  MX4X1 U4013 ( .A(n2208), .B(n2206), .C(n2207), .D(n2205), .S0(n4598), .S1(
        n4539), .Y(n2209) );
  MX4X1 U4014 ( .A(n1945), .B(n1934), .C(n1940), .D(n1929), .S0(n4639), .S1(
        n4628), .Y(n1946) );
  MX4X1 U4015 ( .A(n1933), .B(n1931), .C(n1932), .D(n1930), .S0(n4594), .S1(
        n4535), .Y(n1934) );
  MX4X1 U4016 ( .A(n1928), .B(n1926), .C(n1927), .D(n1925), .S0(n4594), .S1(
        n4535), .Y(n1929) );
  MX4X1 U4017 ( .A(n1944), .B(n1942), .C(n1943), .D(n1941), .S0(n4594), .S1(
        n4536), .Y(n1945) );
  MX4X1 U4018 ( .A(n2032), .B(n2022), .C(n2027), .D(n2017), .S0(n4639), .S1(
        n4629), .Y(n2033) );
  MX4X1 U4019 ( .A(n2021), .B(n2019), .C(n2020), .D(n2018), .S0(n4595), .S1(
        n4537), .Y(n2022) );
  MX4X1 U4020 ( .A(n2016), .B(n2014), .C(n2015), .D(n2013), .S0(n4595), .S1(
        n4537), .Y(n2017) );
  MX4X1 U4021 ( .A(n2031), .B(n2029), .C(n2030), .D(n2028), .S0(n4595), .S1(
        n4537), .Y(n2032) );
  MX4X1 U4022 ( .A(n2620), .B(n2610), .C(n2615), .D(n2605), .S0(n4641), .S1(
        n4630), .Y(n2621) );
  MX4X1 U4023 ( .A(n2609), .B(n2607), .C(n2608), .D(n2606), .S0(n4603), .S1(
        n4532), .Y(n2610) );
  MX4X1 U4024 ( .A(n2604), .B(n2602), .C(n2603), .D(n2601), .S0(n4603), .S1(
        n4537), .Y(n2605) );
  MX4X1 U4025 ( .A(n2619), .B(n2617), .C(n2618), .D(n2616), .S0(n4603), .S1(
        n4539), .Y(n2620) );
  MX4X1 U4026 ( .A(n2296), .B(n2286), .C(n2291), .D(n2281), .S0(n4640), .S1(
        n4629), .Y(n2297) );
  MX4X1 U4027 ( .A(n2285), .B(n2283), .C(n2284), .D(n2282), .S0(n4599), .S1(
        n4540), .Y(n2286) );
  MX4X1 U4028 ( .A(n2280), .B(n2278), .C(n2279), .D(n2277), .S0(n4599), .S1(
        n4540), .Y(n2281) );
  MX4X1 U4029 ( .A(n2295), .B(n2293), .C(n2294), .D(n2292), .S0(n4599), .S1(
        n4540), .Y(n2296) );
  MX4X1 U4030 ( .A(n2450), .B(n2440), .C(n2445), .D(n2380), .S0(n4640), .S1(
        n4630), .Y(n2451) );
  MX4X1 U4031 ( .A(n2439), .B(n2437), .C(n2438), .D(n2382), .S0(n4601), .S1(
        n4542), .Y(n2440) );
  MX4X1 U4032 ( .A(n2379), .B(n2377), .C(n2378), .D(n2376), .S0(n4601), .S1(
        n4541), .Y(n2380) );
  MX4X1 U4033 ( .A(n2449), .B(n2447), .C(n2448), .D(n2446), .S0(n4601), .S1(
        n4542), .Y(n2450) );
  MX4X1 U4034 ( .A(n2960), .B(n2950), .C(n2955), .D(n2945), .S0(n4642), .S1(
        n4632), .Y(n2961) );
  MX4X1 U4035 ( .A(n2949), .B(n2947), .C(n2948), .D(n2946), .S0(n4609), .S1(
        n4548), .Y(n2950) );
  MX4X1 U4036 ( .A(n2944), .B(n2942), .C(n2943), .D(n2941), .S0(n4609), .S1(
        n4548), .Y(n2945) );
  MX4X1 U4037 ( .A(n2959), .B(n2957), .C(n2958), .D(n2956), .S0(n4609), .S1(
        n4548), .Y(n2960) );
  MX4X1 U4038 ( .A(n2705), .B(n2695), .C(n2700), .D(n2690), .S0(n4641), .S1(
        n4631), .Y(n2706) );
  MX4X1 U4039 ( .A(n2694), .B(n2692), .C(n2693), .D(n2691), .S0(n4605), .S1(
        n4544), .Y(n2695) );
  MX4X1 U4040 ( .A(n2689), .B(n2687), .C(n2688), .D(n2686), .S0(n4605), .S1(
        n4544), .Y(n2690) );
  MX4X1 U4041 ( .A(n2704), .B(n2702), .C(n2703), .D(n2701), .S0(n4605), .S1(
        n4544), .Y(n2705) );
  MX4X1 U4042 ( .A(n2790), .B(n2780), .C(n2785), .D(n2775), .S0(n4642), .S1(
        n4631), .Y(n2791) );
  MX4X1 U4043 ( .A(n2779), .B(n2777), .C(n2778), .D(n2776), .S0(n4606), .S1(
        n4545), .Y(n2780) );
  MX4X1 U4044 ( .A(n2774), .B(n2772), .C(n2773), .D(n2771), .S0(n4606), .S1(
        n4545), .Y(n2775) );
  MX4X1 U4045 ( .A(n2789), .B(n2787), .C(n2788), .D(n2786), .S0(n4606), .S1(
        n4546), .Y(n2790) );
  MX4X1 U4046 ( .A(n3300), .B(n3290), .C(n3295), .D(n3285), .S0(n4644), .S1(
        n4633), .Y(n3301) );
  MX4X1 U4047 ( .A(n3289), .B(n3287), .C(n3288), .D(n3286), .S0(n4614), .S1(
        n4553), .Y(n3290) );
  MX4X1 U4048 ( .A(n3284), .B(n3282), .C(n3283), .D(n3281), .S0(n4614), .S1(
        n4553), .Y(n3285) );
  MX4X1 U4049 ( .A(n3299), .B(n3297), .C(n3298), .D(n3296), .S0(n4614), .S1(
        n4553), .Y(n3300) );
  MX4X1 U4050 ( .A(n3045), .B(n3035), .C(n3040), .D(n3030), .S0(n4643), .S1(
        n4632), .Y(n3046) );
  MX4X1 U4051 ( .A(n3034), .B(n3032), .C(n3033), .D(n3031), .S0(n4610), .S1(
        n4549), .Y(n3035) );
  MX4X1 U4052 ( .A(n3029), .B(n3027), .C(n3028), .D(n3026), .S0(n4610), .S1(
        n4549), .Y(n3030) );
  MX4X1 U4053 ( .A(n3044), .B(n3042), .C(n3043), .D(n3041), .S0(n4610), .S1(
        n4549), .Y(n3045) );
  MX4X1 U4054 ( .A(n3130), .B(n3120), .C(n3125), .D(n3115), .S0(n4643), .S1(
        n4632), .Y(n3131) );
  MX4X1 U4055 ( .A(n3119), .B(n3117), .C(n3118), .D(n3116), .S0(n4611), .S1(
        n4550), .Y(n3120) );
  MX4X1 U4056 ( .A(n3114), .B(n3112), .C(n3113), .D(n3111), .S0(n4611), .S1(
        n4550), .Y(n3115) );
  MX4X1 U4057 ( .A(n3129), .B(n3127), .C(n3128), .D(n3126), .S0(n4611), .S1(
        n4551), .Y(n3130) );
  MX4X1 U4058 ( .A(n3640), .B(n3630), .C(n3635), .D(n3625), .S0(n4640), .S1(
        n4634), .Y(n3641) );
  MX4X1 U4059 ( .A(n3629), .B(n3627), .C(n3628), .D(n3626), .S0(n4619), .S1(
        N70), .Y(n3630) );
  MX4X1 U4060 ( .A(n3624), .B(n3622), .C(n3623), .D(n3621), .S0(n4619), .S1(
        N70), .Y(n3625) );
  MX4X1 U4061 ( .A(n3639), .B(n3637), .C(n3638), .D(n3636), .S0(n4619), .S1(
        N70), .Y(n3640) );
  MX4X1 U4062 ( .A(n3385), .B(n3375), .C(n3380), .D(n3370), .S0(n4644), .S1(
        n4633), .Y(n3386) );
  MX4X1 U4063 ( .A(n3374), .B(n3372), .C(n3373), .D(n3371), .S0(n4615), .S1(
        n4554), .Y(n3375) );
  MX4X1 U4064 ( .A(n3369), .B(n3367), .C(n3368), .D(n3366), .S0(n4615), .S1(
        n4554), .Y(n3370) );
  MX4X1 U4065 ( .A(n3384), .B(n3382), .C(n3383), .D(n3381), .S0(n4615), .S1(
        n4554), .Y(n3385) );
  MX4X1 U4066 ( .A(n3470), .B(n3460), .C(n3465), .D(n3455), .S0(n4644), .S1(
        n4633), .Y(n3471) );
  MX4X1 U4067 ( .A(n3459), .B(n3457), .C(n3458), .D(n3456), .S0(n4617), .S1(
        n4555), .Y(n3460) );
  MX4X1 U4068 ( .A(n3454), .B(n3452), .C(n3453), .D(n3451), .S0(n4617), .S1(
        n4555), .Y(n3455) );
  MX4X1 U4069 ( .A(n3469), .B(n3467), .C(n3468), .D(n3466), .S0(n4617), .S1(
        n4555), .Y(n3470) );
  MX4X1 U4070 ( .A(n3980), .B(n3970), .C(n3975), .D(n3965), .S0(n4645), .S1(
        n4635), .Y(n3981) );
  MX4X1 U4071 ( .A(n3969), .B(n3967), .C(n3968), .D(n3966), .S0(N71), .S1(
        n4559), .Y(n3970) );
  MX4X1 U4072 ( .A(n3964), .B(n3962), .C(n3963), .D(n3961), .S0(n4592), .S1(
        n4559), .Y(n3965) );
  MX4X1 U4073 ( .A(n3979), .B(n3977), .C(n3978), .D(n3976), .S0(N71), .S1(
        n4559), .Y(n3980) );
  MX4X1 U4074 ( .A(n3725), .B(n3715), .C(n3720), .D(n3710), .S0(n4641), .S1(
        n4634), .Y(n3726) );
  MX4X1 U4075 ( .A(n3714), .B(n3712), .C(n3713), .D(n3711), .S0(n4621), .S1(
        n4542), .Y(n3715) );
  MX4X1 U4076 ( .A(n3709), .B(n3707), .C(n3708), .D(n3706), .S0(n4621), .S1(
        n4536), .Y(n3710) );
  MX4X1 U4077 ( .A(n3724), .B(n3722), .C(n3723), .D(n3721), .S0(n4621), .S1(
        n4541), .Y(n3725) );
  MX4X1 U4078 ( .A(n3810), .B(n3800), .C(n3805), .D(n3795), .S0(n4645), .S1(
        n4635), .Y(n3811) );
  MX4X1 U4079 ( .A(n3799), .B(n3797), .C(n3798), .D(n3796), .S0(n4622), .S1(
        n4529), .Y(n3800) );
  MX4X1 U4080 ( .A(n3794), .B(n3792), .C(n3793), .D(n3791), .S0(n4622), .S1(
        n4534), .Y(n3795) );
  MX4X1 U4081 ( .A(n3809), .B(n3807), .C(n3808), .D(n3806), .S0(n4622), .S1(
        n4534), .Y(n3810) );
  MX4X1 U4082 ( .A(n4945), .B(n4935), .C(n4940), .D(n4930), .S0(n7981), .S1(
        n7972), .Y(n4946) );
  MX4X1 U4083 ( .A(n4934), .B(n4932), .C(n4933), .D(n4931), .S0(n7930), .S1(
        n7870), .Y(n4935) );
  MX4X1 U4084 ( .A(n4929), .B(n4927), .C(n4928), .D(n4926), .S0(n7930), .S1(
        n7870), .Y(n4930) );
  MX4X1 U4085 ( .A(n4944), .B(n4942), .C(n4943), .D(n4941), .S0(n7930), .S1(
        n7870), .Y(n4945) );
  MX4X1 U4086 ( .A(n5285), .B(n5275), .C(n5280), .D(n5270), .S0(n7982), .S1(
        n7973), .Y(n5286) );
  MX4X1 U4087 ( .A(n5274), .B(n5272), .C(n5273), .D(n5271), .S0(n7936), .S1(
        n7875), .Y(n5275) );
  MX4X1 U4088 ( .A(n5269), .B(n5267), .C(n5268), .D(n5266), .S0(n7936), .S1(
        n7875), .Y(n5270) );
  MX4X1 U4089 ( .A(n5284), .B(n5282), .C(n5283), .D(n5281), .S0(n7936), .S1(
        n7875), .Y(n5285) );
  MX4X1 U4090 ( .A(n5030), .B(n5020), .C(n5025), .D(n5015), .S0(n7981), .S1(
        n7972), .Y(n5031) );
  MX4X1 U4091 ( .A(n5019), .B(n5017), .C(n5018), .D(n5016), .S0(n7932), .S1(
        n7871), .Y(n5020) );
  MX4X1 U4092 ( .A(n5014), .B(n5012), .C(n5013), .D(n5011), .S0(n7932), .S1(
        n7871), .Y(n5015) );
  MX4X1 U4093 ( .A(n5029), .B(n5027), .C(n5028), .D(n5026), .S0(n7932), .S1(
        n7872), .Y(n5030) );
  MX4X1 U4094 ( .A(n5115), .B(n5105), .C(n5110), .D(n5100), .S0(n7982), .S1(
        n7972), .Y(n5116) );
  MX4X1 U4095 ( .A(n5104), .B(n5102), .C(n5103), .D(n5101), .S0(n7933), .S1(
        n7873), .Y(n5105) );
  MX4X1 U4096 ( .A(n5099), .B(n5097), .C(n5098), .D(n5096), .S0(n7933), .S1(
        n7873), .Y(n5100) );
  MX4X1 U4097 ( .A(n5114), .B(n5112), .C(n5113), .D(n5111), .S0(n7933), .S1(
        n7873), .Y(n5115) );
  MX4X1 U4098 ( .A(n5625), .B(n5615), .C(n5620), .D(n5610), .S0(n7983), .S1(
        n7974), .Y(n5626) );
  MX4X1 U4099 ( .A(n5614), .B(n5612), .C(n5613), .D(n5611), .S0(n7941), .S1(
        n7880), .Y(n5615) );
  MX4X1 U4100 ( .A(n5609), .B(n5607), .C(n5608), .D(n5606), .S0(n7941), .S1(
        n7880), .Y(n5610) );
  MX4X1 U4101 ( .A(n5624), .B(n5622), .C(n5623), .D(n5621), .S0(n7941), .S1(
        n7880), .Y(n5625) );
  MX4X1 U4102 ( .A(n5370), .B(n5360), .C(n5365), .D(n5355), .S0(n7987), .S1(
        n7973), .Y(n5371) );
  MX4X1 U4103 ( .A(n5359), .B(n5357), .C(n5358), .D(n5356), .S0(n7937), .S1(
        n7876), .Y(n5360) );
  MX4X1 U4104 ( .A(n5354), .B(n5352), .C(n5353), .D(n5351), .S0(n7937), .S1(
        n7876), .Y(n5355) );
  MX4X1 U4105 ( .A(n5369), .B(n5367), .C(n5368), .D(n5366), .S0(n7937), .S1(
        n7877), .Y(n5370) );
  MX4X1 U4106 ( .A(n5455), .B(n5445), .C(n5450), .D(n5440), .S0(n7980), .S1(
        n7974), .Y(n5456) );
  MX4X1 U4107 ( .A(n5444), .B(n5442), .C(n5443), .D(n5441), .S0(n7938), .S1(
        n7878), .Y(n5445) );
  MX4X1 U4108 ( .A(n5439), .B(n5437), .C(n5438), .D(n5436), .S0(n7938), .S1(
        n7878), .Y(n5440) );
  MX4X1 U4109 ( .A(n5454), .B(n5452), .C(n5453), .D(n5451), .S0(n7938), .S1(
        n7878), .Y(n5455) );
  MX4X1 U4110 ( .A(n5965), .B(n5955), .C(n5960), .D(n5950), .S0(n7984), .S1(
        n7975), .Y(n5966) );
  MX4X1 U4111 ( .A(n5954), .B(n5952), .C(n5953), .D(n5951), .S0(n7946), .S1(
        n7885), .Y(n5955) );
  MX4X1 U4112 ( .A(n5949), .B(n5947), .C(n5948), .D(n5946), .S0(n7946), .S1(
        n7885), .Y(n5950) );
  MX4X1 U4113 ( .A(n5964), .B(n5962), .C(n5963), .D(n5961), .S0(n7946), .S1(
        n7885), .Y(n5965) );
  MX4X1 U4114 ( .A(n5710), .B(n5700), .C(n5705), .D(n5695), .S0(n7983), .S1(
        n7974), .Y(n5711) );
  MX4X1 U4115 ( .A(n5699), .B(n5697), .C(n5698), .D(n5696), .S0(n7942), .S1(
        n7881), .Y(n5700) );
  MX4X1 U4116 ( .A(n5694), .B(n5692), .C(n5693), .D(n5691), .S0(n7942), .S1(
        n7881), .Y(n5695) );
  MX4X1 U4117 ( .A(n5709), .B(n5707), .C(n5708), .D(n5706), .S0(n7942), .S1(
        n7881), .Y(n5710) );
  MX4X1 U4118 ( .A(n5795), .B(n5785), .C(n5790), .D(n5780), .S0(n7983), .S1(
        n7975), .Y(n5796) );
  MX4X1 U4119 ( .A(n5784), .B(n5782), .C(n5783), .D(n5781), .S0(n7944), .S1(
        n7883), .Y(n5785) );
  MX4X1 U4120 ( .A(n5779), .B(n5777), .C(n5778), .D(n5776), .S0(n7944), .S1(
        n7882), .Y(n5780) );
  MX4X1 U4121 ( .A(n5794), .B(n5792), .C(n5793), .D(n5791), .S0(n7944), .S1(
        n7883), .Y(n5795) );
  MX4X1 U4122 ( .A(n6305), .B(n6295), .C(n6300), .D(n6290), .S0(n7985), .S1(
        n7977), .Y(n6306) );
  MX4X1 U4123 ( .A(n6294), .B(n6292), .C(n6293), .D(n6291), .S0(n7952), .S1(
        n7890), .Y(n6295) );
  MX4X1 U4124 ( .A(n6289), .B(n6287), .C(n6288), .D(n6286), .S0(n7952), .S1(
        n7890), .Y(n6290) );
  MX4X1 U4125 ( .A(n6304), .B(n6302), .C(n6303), .D(n6301), .S0(n7952), .S1(
        n7890), .Y(n6305) );
  MX4X1 U4126 ( .A(n6050), .B(n6040), .C(n6045), .D(n6035), .S0(n7984), .S1(
        n7976), .Y(n6051) );
  MX4X1 U4127 ( .A(n6039), .B(n6037), .C(n6038), .D(n6036), .S0(n7948), .S1(
        n7886), .Y(n6040) );
  MX4X1 U4128 ( .A(n6034), .B(n6032), .C(n6033), .D(n6031), .S0(n7948), .S1(
        n7886), .Y(n6035) );
  MX4X1 U4129 ( .A(n6049), .B(n6047), .C(n6048), .D(n6046), .S0(n7948), .S1(
        n7886), .Y(n6050) );
  MX4X1 U4130 ( .A(n6135), .B(n6125), .C(n6130), .D(n6120), .S0(n7985), .S1(
        n7976), .Y(n6136) );
  MX4X1 U4131 ( .A(n6124), .B(n6122), .C(n6123), .D(n6121), .S0(n7949), .S1(
        n7887), .Y(n6125) );
  MX4X1 U4132 ( .A(n6119), .B(n6117), .C(n6118), .D(n6116), .S0(n7949), .S1(
        n7887), .Y(n6120) );
  MX4X1 U4133 ( .A(n6134), .B(n6132), .C(n6133), .D(n6131), .S0(n7949), .S1(
        n7888), .Y(n6135) );
  MX4X1 U4134 ( .A(n6645), .B(n6635), .C(n6640), .D(n6630), .S0(n7987), .S1(
        n7975), .Y(n6646) );
  MX4X1 U4135 ( .A(n6634), .B(n6632), .C(n6633), .D(n6631), .S0(n7957), .S1(
        n7895), .Y(n6635) );
  MX4X1 U4136 ( .A(n6629), .B(n6627), .C(n6628), .D(n6626), .S0(n7957), .S1(
        n7895), .Y(n6630) );
  MX4X1 U4137 ( .A(n6644), .B(n6642), .C(n6643), .D(n6641), .S0(n7957), .S1(
        n7895), .Y(n6645) );
  MX4X1 U4138 ( .A(n6390), .B(n6380), .C(n6385), .D(n6375), .S0(n7986), .S1(
        n7977), .Y(n6391) );
  MX4X1 U4139 ( .A(n6379), .B(n6377), .C(n6378), .D(n6376), .S0(n7953), .S1(
        n7891), .Y(n6380) );
  MX4X1 U4140 ( .A(n6374), .B(n6372), .C(n6373), .D(n6371), .S0(n7953), .S1(
        n7891), .Y(n6375) );
  MX4X1 U4141 ( .A(n6389), .B(n6387), .C(n6388), .D(n6386), .S0(n7953), .S1(
        n7891), .Y(n6390) );
  MX4X1 U4142 ( .A(n6475), .B(n6465), .C(n6470), .D(n6460), .S0(n7986), .S1(
        n7977), .Y(n6476) );
  MX4X1 U4143 ( .A(n6464), .B(n6462), .C(n6463), .D(n6461), .S0(n7954), .S1(
        n7892), .Y(n6465) );
  MX4X1 U4144 ( .A(n6459), .B(n6457), .C(n6458), .D(n6456), .S0(n7954), .S1(
        n7892), .Y(n6460) );
  MX4X1 U4145 ( .A(n6474), .B(n6472), .C(n6473), .D(n6471), .S0(n7954), .S1(
        n7893), .Y(n6475) );
  MX4X1 U4146 ( .A(n6985), .B(n6975), .C(n6980), .D(n6970), .S0(n7988), .S1(
        n8644), .Y(n6986) );
  MX4X1 U4147 ( .A(n6974), .B(n6972), .C(n6973), .D(n6971), .S0(n7962), .S1(
        n7898), .Y(n6975) );
  MX4X1 U4148 ( .A(n6969), .B(n6967), .C(n6968), .D(n6966), .S0(n7962), .S1(
        n7898), .Y(n6970) );
  MX4X1 U4149 ( .A(n6984), .B(n6982), .C(n6983), .D(n6981), .S0(n7962), .S1(
        n7898), .Y(n6985) );
  MX4X1 U4150 ( .A(n6730), .B(n6720), .C(n6725), .D(n6715), .S0(n7987), .S1(
        n8644), .Y(n6731) );
  MX4X1 U4151 ( .A(n6719), .B(n6717), .C(n6718), .D(n6716), .S0(n7958), .S1(
        n7896), .Y(n6720) );
  MX4X1 U4152 ( .A(n6714), .B(n6712), .C(n6713), .D(n6711), .S0(n7958), .S1(
        n7896), .Y(n6715) );
  MX4X1 U4153 ( .A(n6729), .B(n6727), .C(n6728), .D(n6726), .S0(n7958), .S1(
        n7896), .Y(n6730) );
  MX4X1 U4154 ( .A(n6815), .B(n6805), .C(n6810), .D(n6800), .S0(n7987), .S1(
        n7971), .Y(n6816) );
  MX4X1 U4155 ( .A(n6804), .B(n6802), .C(n6803), .D(n6801), .S0(n7960), .S1(
        n7899), .Y(n6805) );
  MX4X1 U4156 ( .A(n6799), .B(n6797), .C(n6798), .D(n6796), .S0(n7960), .S1(
        n7869), .Y(n6800) );
  MX4X1 U4157 ( .A(n6814), .B(n6812), .C(n6813), .D(n6811), .S0(n7960), .S1(
        n7868), .Y(n6815) );
  MX4X1 U4158 ( .A(n7325), .B(n7315), .C(n7320), .D(n7310), .S0(n7985), .S1(
        N82), .Y(n7326) );
  MX4X1 U4159 ( .A(n7314), .B(n7312), .C(n7313), .D(n7311), .S0(N81), .S1(
        n7902), .Y(n7315) );
  MX4X1 U4160 ( .A(n7309), .B(n7307), .C(n7308), .D(n7306), .S0(n7935), .S1(
        n7902), .Y(n7310) );
  MX4X1 U4161 ( .A(n7324), .B(n7322), .C(n7323), .D(n7321), .S0(N81), .S1(
        n7902), .Y(n7325) );
  MX4X1 U4162 ( .A(n7070), .B(n7060), .C(n7065), .D(n7055), .S0(n7988), .S1(
        n7973), .Y(n7071) );
  MX4X1 U4163 ( .A(n7059), .B(n7057), .C(n7058), .D(n7056), .S0(n7964), .S1(
        n7899), .Y(n7060) );
  MX4X1 U4164 ( .A(n7054), .B(n7052), .C(n7053), .D(n7051), .S0(n7964), .S1(
        n7899), .Y(n7055) );
  MX4X1 U4165 ( .A(n7069), .B(n7067), .C(n7068), .D(n7066), .S0(n7964), .S1(
        n7899), .Y(n7070) );
  MX4X1 U4166 ( .A(n7155), .B(n7145), .C(n7150), .D(n7140), .S0(n7986), .S1(
        N82), .Y(n7156) );
  MX4X1 U4167 ( .A(n7144), .B(n7142), .C(n7143), .D(n7141), .S0(n7965), .S1(
        n7900), .Y(n7145) );
  MX4X1 U4168 ( .A(n7139), .B(n7137), .C(n7138), .D(n7136), .S0(n7965), .S1(
        n7900), .Y(n7140) );
  MX4X1 U4169 ( .A(n7154), .B(n7152), .C(n7153), .D(n7151), .S0(n7965), .S1(
        n7900), .Y(n7155) );
  MX4X1 U4170 ( .A(n1064), .B(n1054), .C(n1059), .D(n1049), .S0(n4637), .S1(
        n4635), .Y(n1065) );
  MX4X1 U4171 ( .A(n1053), .B(n1051), .C(n1052), .D(n1050), .S0(n4620), .S1(
        n4525), .Y(n1054) );
  MX4X1 U4172 ( .A(n1048), .B(n1046), .C(n1047), .D(n1045), .S0(n4623), .S1(
        n4525), .Y(n1049) );
  MX4X1 U4173 ( .A(n1063), .B(n1061), .C(n1062), .D(n1060), .S0(n4623), .S1(
        n4525), .Y(n1064) );
  MX4X1 U4174 ( .A(n1207), .B(n1181), .C(n1198), .D(n1176), .S0(n4645), .S1(
        n4634), .Y(n1209) );
  MX4X1 U4175 ( .A(n1180), .B(n1178), .C(n1179), .D(n1177), .S0(n4590), .S1(
        n4526), .Y(n1181) );
  MX4X1 U4176 ( .A(n1175), .B(n1173), .C(n1174), .D(n1172), .S0(n4587), .S1(
        n4526), .Y(n1176) );
  MX4X1 U4177 ( .A(n1205), .B(n1202), .C(n1204), .D(n1201), .S0(n4608), .S1(
        n4527), .Y(n1207) );
  MX4X1 U4178 ( .A(n4669), .B(n4659), .C(n4664), .D(n4654), .S0(n7981), .S1(
        n7971), .Y(n4670) );
  MX4X1 U4179 ( .A(n4658), .B(n4656), .C(n4657), .D(n4655), .S0(n7963), .S1(
        n7866), .Y(n4659) );
  MX4X1 U4180 ( .A(n4653), .B(n4651), .C(n4652), .D(n4650), .S0(n7966), .S1(
        n7866), .Y(n4654) );
  MX4X1 U4181 ( .A(n4668), .B(n4666), .C(n4667), .D(n4665), .S0(n7966), .S1(
        n7866), .Y(n4669) );
  MX4X1 U4182 ( .A(n1085), .B(n1075), .C(n1080), .D(n1070), .S0(n4637), .S1(
        n4635), .Y(n1086) );
  MX4X1 U4183 ( .A(n1074), .B(n1072), .C(n1073), .D(n1071), .S0(n4587), .S1(
        n4526), .Y(n1075) );
  MX4X1 U4184 ( .A(n1069), .B(n1067), .C(n1068), .D(n1066), .S0(n4621), .S1(
        n4525), .Y(n1070) );
  MX4X1 U4185 ( .A(n1084), .B(n1082), .C(n1083), .D(n1081), .S0(n4622), .S1(
        n4526), .Y(n1085) );
  MX4X1 U4186 ( .A(n1307), .B(n1287), .C(n1297), .D(n1277), .S0(N73), .S1(N72), 
        .Y(n1309) );
  MX4X1 U4187 ( .A(n1285), .B(n1281), .C(n1283), .D(n1279), .S0(n4614), .S1(
        n4527), .Y(n1287) );
  MX4X1 U4188 ( .A(n1275), .B(n1270), .C(n1273), .D(n1210), .S0(n4596), .S1(
        n4527), .Y(n1277) );
  MX4X1 U4189 ( .A(n1305), .B(n1301), .C(n1303), .D(n1299), .S0(n4603), .S1(
        n4527), .Y(n1307) );
  MX4X1 U4190 ( .A(n4690), .B(n4680), .C(n4685), .D(n4675), .S0(n7981), .S1(
        n7971), .Y(n4691) );
  MX4X1 U4191 ( .A(n4679), .B(n4677), .C(n4678), .D(n4676), .S0(n7930), .S1(
        n7867), .Y(n4680) );
  MX4X1 U4192 ( .A(n4674), .B(n4672), .C(n4673), .D(n4671), .S0(n7964), .S1(
        n7866), .Y(n4675) );
  MX4X1 U4193 ( .A(n4689), .B(n4687), .C(n4688), .D(n4686), .S0(n7965), .S1(
        n7867), .Y(n4690) );
  MX4X1 U4194 ( .A(n4775), .B(n4765), .C(n4770), .D(n4760), .S0(N83), .S1(
        n7971), .Y(n4776) );
  MX4X1 U4195 ( .A(n4764), .B(n4762), .C(n4763), .D(n4761), .S0(n7957), .S1(
        n7868), .Y(n4765) );
  MX4X1 U4196 ( .A(n4759), .B(n4757), .C(n4758), .D(n4756), .S0(n7939), .S1(
        n7868), .Y(n4760) );
  MX4X1 U4197 ( .A(n4774), .B(n4772), .C(n4773), .D(n4771), .S0(n7946), .S1(
        n7868), .Y(n4775) );
  INVX1 U4198 ( .A(n4502), .Y(n4503) );
  INVX1 U4199 ( .A(n8658), .Y(n4502) );
  INVX1 U4200 ( .A(n8659), .Y(n8658) );
  INVX1 U4201 ( .A(N69), .Y(n8659) );
  AOI21X2 U4202 ( .A0(n1267), .A1(n8660), .B0(rst), .Y(n1266) );
  NOR3X2 U4203 ( .A(Address[0]), .B(Address[2]), .C(n8971), .Y(n2342) );
  NOR2X2 U4204 ( .A(n8967), .B(Address[9]), .Y(n1606) );
  NOR2BX2 U4205 ( .AN(Address[9]), .B(Address[8]), .Y(n1871) );
  NOR2BX2 U4206 ( .AN(Address[9]), .B(n8967), .Y(n2136) );
  NOR2X2 U4207 ( .A(Address[8]), .B(Address[9]), .Y(n1366) );
  NOR2X2 U4208 ( .A(n8970), .B(Address[4]), .Y(n2354) );
  NOR2BX2 U4209 ( .AN(Address[4]), .B(Address[3]), .Y(n2363) );
  NOR2BX2 U4210 ( .AN(Address[4]), .B(n8970), .Y(n2372) );
  NOR3X2 U4211 ( .A(Address[1]), .B(Address[2]), .C(Address[0]), .Y(n2337) );
  NOR3X2 U4212 ( .A(Address[1]), .B(Address[2]), .C(n8972), .Y(n2340) );
  NOR3X2 U4213 ( .A(n8972), .B(Address[2]), .C(n8971), .Y(n2344) );
  NOR3X2 U4214 ( .A(Address[6]), .B(Address[7]), .C(n8969), .Y(n1367) );
  NOR3X2 U4215 ( .A(Address[5]), .B(Address[7]), .C(n8968), .Y(n1401) );
  NOR3X2 U4216 ( .A(n8969), .B(Address[7]), .C(n8968), .Y(n1435) );
  BUFX3 U4217 ( .A(n2338), .Y(n8439) );
  NOR2X1 U4218 ( .A(Address[3]), .B(Address[4]), .Y(n2338) );
  INVX1 U4219 ( .A(Address[5]), .Y(n8969) );
  INVX1 U4220 ( .A(Address[0]), .Y(n8972) );
  INVX1 U4221 ( .A(Address[6]), .Y(n8968) );
  INVX1 U4222 ( .A(Address[1]), .Y(n8971) );
  INVX1 U4223 ( .A(Address[8]), .Y(n8967) );
  INVX1 U4224 ( .A(Address[3]), .Y(n8970) );
  NOR3X2 U4225 ( .A(Address[6]), .B(Address[7]), .C(Address[5]), .Y(n1605) );
  AND3X2 U4226 ( .A(n8972), .B(n8971), .C(Address[2]), .Y(n2346) );
  INVX1 U4227 ( .A(n1212), .Y(n8960) );
  AND3X2 U4228 ( .A(Address[0]), .B(n8971), .C(Address[2]), .Y(n2348) );
  AND3X2 U4229 ( .A(Address[1]), .B(n8972), .C(Address[2]), .Y(n2350) );
  AND3X2 U4230 ( .A(Address[1]), .B(Address[0]), .C(Address[2]), .Y(n2352) );
  AND3X2 U4231 ( .A(n8969), .B(n8968), .C(Address[7]), .Y(n1469) );
  AND3X2 U4232 ( .A(Address[5]), .B(n8968), .C(Address[7]), .Y(n1503) );
  AND3X2 U4233 ( .A(Address[6]), .B(n8969), .C(Address[7]), .Y(n1537) );
  AND3X2 U4234 ( .A(Address[6]), .B(Address[5]), .C(Address[7]), .Y(n1571) );
  CLKINVX3 U4235 ( .A(n8662), .Y(n8660) );
  INVX1 U4236 ( .A(ena_in), .Y(n8662) );
  NOR2X1 U4237 ( .A(n1200), .B(n1206), .Y(n1187) );
  AOI21X1 U4238 ( .A0(n8964), .A1(n8961), .B0(n8958), .Y(n1239) );
  NAND2X1 U4239 ( .A(n1212), .B(n1241), .Y(n1197) );
  OAI22X1 U4240 ( .A0(n1237), .A1(n8966), .B0(n8965), .B1(n1238), .Y(n2426) );
  NOR2BX1 U4241 ( .AN(n1239), .B(n8961), .Y(n1237) );
  BUFX3 U4242 ( .A(n1196), .Y(n8443) );
  NAND3X1 U4243 ( .A(n8964), .B(n8966), .C(n1189), .Y(n1196) );
  BUFX3 U4244 ( .A(n1193), .Y(n8444) );
  NAND2X1 U4245 ( .A(n1192), .B(n8964), .Y(n1193) );
  BUFX3 U4246 ( .A(n1243), .Y(n8440) );
  NOR2X1 U4247 ( .A(rst), .B(n1257), .Y(n1243) );
  INVX1 U4248 ( .A(n8765), .Y(n8768) );
  INVX1 U4249 ( .A(n8692), .Y(n8719) );
  INVX1 U4250 ( .A(n8720), .Y(n8747) );
  NOR2X1 U4251 ( .A(n8966), .B(n8965), .Y(n1186) );
  INVX1 U4252 ( .A(rst), .Y(n8973) );
  INVX1 U4253 ( .A(n1217), .Y(n8956) );
  AOI22X1 U4254 ( .A0(N1366), .A1(n8442), .B0(block_i[17]), .B1(n8436), .Y(
        n1217) );
  INVX1 U4255 ( .A(n1219), .Y(n8955) );
  AOI22X1 U4256 ( .A0(N1365), .A1(n8442), .B0(block_i[16]), .B1(n8436), .Y(
        n1219) );
  INVX1 U4257 ( .A(n1220), .Y(n8954) );
  AOI22X1 U4258 ( .A0(N1364), .A1(n8442), .B0(block_i[15]), .B1(n8436), .Y(
        n1220) );
  INVX1 U4259 ( .A(n1221), .Y(n8953) );
  AOI22X1 U4260 ( .A0(N1363), .A1(n8442), .B0(block_i[14]), .B1(n8436), .Y(
        n1221) );
  INVX1 U4261 ( .A(n1222), .Y(n8952) );
  AOI22X1 U4262 ( .A0(N1362), .A1(n8442), .B0(block_i[13]), .B1(n8436), .Y(
        n1222) );
  INVX1 U4263 ( .A(n1223), .Y(n8951) );
  AOI22X1 U4264 ( .A0(N1361), .A1(n8442), .B0(block_i[12]), .B1(n8436), .Y(
        n1223) );
  INVX1 U4265 ( .A(n1224), .Y(n8950) );
  AOI22X1 U4266 ( .A0(N1360), .A1(n8442), .B0(block_i[11]), .B1(n8436), .Y(
        n1224) );
  INVX1 U4267 ( .A(n1225), .Y(n8949) );
  AOI22X1 U4268 ( .A0(N1359), .A1(n8442), .B0(block_i[10]), .B1(n8436), .Y(
        n1225) );
  INVX1 U4269 ( .A(n1226), .Y(n8948) );
  AOI22X1 U4270 ( .A0(N1358), .A1(n8442), .B0(block_i[9]), .B1(n8435), .Y(
        n1226) );
  INVX1 U4271 ( .A(n1227), .Y(n8947) );
  AOI22X1 U4272 ( .A0(N1357), .A1(n8442), .B0(block_i[8]), .B1(n8435), .Y(
        n1227) );
  INVX1 U4273 ( .A(n1228), .Y(n8946) );
  AOI22X1 U4274 ( .A0(N1356), .A1(n8442), .B0(block_i[7]), .B1(n8435), .Y(
        n1228) );
  INVX1 U4275 ( .A(n1229), .Y(n8945) );
  AOI22X1 U4276 ( .A0(N1355), .A1(n8442), .B0(block_i[6]), .B1(n8435), .Y(
        n1229) );
  INVX1 U4277 ( .A(n1230), .Y(n8944) );
  AOI22X1 U4278 ( .A0(N1354), .A1(n8442), .B0(block_i[5]), .B1(n8435), .Y(
        n1230) );
  INVX1 U4279 ( .A(n1231), .Y(n8943) );
  AOI22X1 U4280 ( .A0(N1353), .A1(n8442), .B0(block_i[4]), .B1(n8435), .Y(
        n1231) );
  INVX1 U4281 ( .A(n1232), .Y(n8942) );
  AOI22X1 U4282 ( .A0(N1352), .A1(n8442), .B0(block_i[3]), .B1(n8435), .Y(
        n1232) );
  INVX1 U4283 ( .A(n1233), .Y(n8941) );
  AOI22X1 U4284 ( .A0(N1351), .A1(n8442), .B0(block_i[2]), .B1(n8435), .Y(
        n1233) );
  INVX1 U4285 ( .A(n1234), .Y(n8940) );
  AOI22X1 U4286 ( .A0(N1350), .A1(n8442), .B0(block_i[1]), .B1(n8435), .Y(
        n1234) );
  INVX1 U4287 ( .A(n1235), .Y(n8939) );
  INVX1 U4288 ( .A(n1236), .Y(n8938) );
  AOI22X1 U4289 ( .A0(N1367), .A1(n8442), .B0(block_i[18]), .B1(n8435), .Y(
        n1236) );
  OAI31X1 U4290 ( .A0(n8937), .A1(n8436), .A2(n8960), .B0(n1216), .Y(n2425) );
  NAND2X1 U4291 ( .A(Image_Done), .B(n8436), .Y(n1216) );
  INVX1 U4292 ( .A(N1408), .Y(n8937) );
  INVX1 U4293 ( .A(n8664), .Y(n8663) );
  INVX1 U4294 ( .A(data_in[0]), .Y(n8664) );
  INVX1 U4295 ( .A(n8693), .Y(n8692) );
  INVX1 U4296 ( .A(data_in[1]), .Y(n8693) );
  INVX1 U4297 ( .A(n8721), .Y(n8720) );
  INVX1 U4298 ( .A(data_in[2]), .Y(n8721) );
  INVX1 U4299 ( .A(n8749), .Y(n8748) );
  INVX1 U4300 ( .A(data_in[3]), .Y(n8749) );
  INVX1 U4301 ( .A(n8772), .Y(n8771) );
  INVX1 U4302 ( .A(data_in[4]), .Y(n8772) );
  INVX1 U4303 ( .A(n8801), .Y(n8800) );
  INVX1 U4304 ( .A(data_in[5]), .Y(n8801) );
  INVX1 U4305 ( .A(n8830), .Y(n8829) );
  INVX1 U4306 ( .A(data_in[6]), .Y(n8830) );
  INVX1 U4307 ( .A(n8859), .Y(n8858) );
  INVX1 U4308 ( .A(data_in[7]), .Y(n8859) );
  NOR2BX1 U4309 ( .AN(n1208), .B(pixel_i[1]), .Y(n1203) );
  AND2X2 U4310 ( .A(n1208), .B(pixel_i[1]), .Y(n1199) );
  AND3X2 U4311 ( .A(N1197), .B(n1199), .C(n1206), .Y(n1040) );
  AND3X2 U4312 ( .A(N1197), .B(n1200), .C(n1203), .Y(n1041) );
  AND3X2 U4313 ( .A(n1203), .B(N1197), .C(n1206), .Y(n1042) );
  AND3X2 U4314 ( .A(n1199), .B(n1200), .C(N1197), .Y(n1043) );
  AND4X2 U4315 ( .A(n1211), .B(n1212), .C(n1213), .D(n1214), .Y(n1208) );
  NOR3X1 U4316 ( .A(pixel_i[11]), .B(pixel_i[2]), .C(pixel_i[12]), .Y(n1213)
         );
  NOR2XL U4317 ( .A(pixel_i[10]), .B(N1195), .Y(n1211) );
  INVX1 U4318 ( .A(pixel_i[3]), .Y(n8916) );
  INVX1 U4319 ( .A(N1197), .Y(n8915) );
  INVX1 U4320 ( .A(n1255), .Y(n8925) );
  AOI22X1 U4321 ( .A0(N1197), .A1(n8440), .B0(N1235), .B1(n8441), .Y(n1255) );
  INVX1 U4322 ( .A(n1252), .Y(n8928) );
  AOI22X1 U4323 ( .A0(n8440), .A1(pixel_i[3]), .B0(N1238), .B1(n8441), .Y(
        n1252) );
  INVX1 U4324 ( .A(n1249), .Y(n8931) );
  AOI22X1 U4325 ( .A0(n8440), .A1(pixel_i[6]), .B0(N1241), .B1(n8441), .Y(
        n1249) );
  INVX1 U4326 ( .A(n1254), .Y(n8926) );
  AOI22X1 U4327 ( .A0(pixel_i[1]), .A1(n8440), .B0(N1236), .B1(n8441), .Y(
        n1254) );
  INVX1 U4328 ( .A(n1251), .Y(n8929) );
  AOI22X1 U4329 ( .A0(n8440), .A1(pixel_i[4]), .B0(N1239), .B1(n8441), .Y(
        n1251) );
  INVX1 U4330 ( .A(n1253), .Y(n8927) );
  AOI22X1 U4331 ( .A0(n8440), .A1(pixel_i[2]), .B0(N1237), .B1(n8441), .Y(
        n1253) );
  INVX1 U4332 ( .A(n1246), .Y(n8934) );
  AOI22X1 U4333 ( .A0(n8440), .A1(pixel_i[9]), .B0(N1244), .B1(n8441), .Y(
        n1246) );
  INVX1 U4334 ( .A(n1248), .Y(n8932) );
  AOI22X1 U4335 ( .A0(n8440), .A1(pixel_i[7]), .B0(N1242), .B1(n8441), .Y(
        n1248) );
  INVX1 U4336 ( .A(n1250), .Y(n8930) );
  INVX1 U4337 ( .A(n1247), .Y(n8933) );
  INVX1 U4338 ( .A(n1245), .Y(n8935) );
  AOI22X1 U4339 ( .A0(n8440), .A1(pixel_i[10]), .B0(N1245), .B1(n8441), .Y(
        n1245) );
  INVX1 U4340 ( .A(n1242), .Y(n8936) );
  AOI22X1 U4341 ( .A0(n8440), .A1(pixel_i[11]), .B0(N1246), .B1(n8441), .Y(
        n1242) );
  INVX1 U4342 ( .A(n1256), .Y(n8924) );
  AOI22X1 U4343 ( .A0(n8440), .A1(pixel_i[12]), .B0(N1247), .B1(n8441), .Y(
        n1256) );
  INVX1 U4344 ( .A(pixel_i[8]), .Y(n8917) );
  INVX1 U4345 ( .A(n1258), .Y(n8921) );
  AOI32X1 U4346 ( .A0(n1206), .A1(n8923), .A2(n1212), .B0(state[0]), .B1(n1259), .Y(n1258) );
  INVX1 U4347 ( .A(n1260), .Y(n8922) );
  AOI32X1 U4348 ( .A0(n1200), .A1(n8923), .A2(n1212), .B0(n1259), .B1(state[1]), .Y(n1260) );
  MX4X1 U4349 ( .A(\registers[1012][0] ), .B(\registers[1013][0] ), .C(
        \registers[1014][0] ), .D(\registers[1015][0] ), .S0(n4106), .S1(n4350), .Y(n1047) );
  MX4X1 U4350 ( .A(\registers[996][0] ), .B(\registers[997][0] ), .C(
        \registers[998][0] ), .D(\registers[999][0] ), .S0(n4250), .S1(n4501), 
        .Y(n1052) );
  MX4X1 U4351 ( .A(\registers[1012][0] ), .B(\registers[1013][0] ), .C(
        \registers[1014][0] ), .D(\registers[1015][0] ), .S0(n7578), .S1(n7808), .Y(n4652) );
  MX4X1 U4352 ( .A(\registers[996][0] ), .B(\registers[997][0] ), .C(
        \registers[998][0] ), .D(\registers[999][0] ), .S0(n7607), .S1(n7811), 
        .Y(n4657) );
  MX4X1 U4353 ( .A(\registers[340][0] ), .B(\registers[341][0] ), .C(
        \registers[342][0] ), .D(\registers[343][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1425) );
  MX4X1 U4354 ( .A(\registers[324][0] ), .B(\registers[325][0] ), .C(
        \registers[326][0] ), .D(\registers[327][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1430) );
  MX4X1 U4355 ( .A(\registers[372][0] ), .B(\registers[373][0] ), .C(
        \registers[374][0] ), .D(\registers[375][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1415) );
  MX4X1 U4356 ( .A(\registers[356][0] ), .B(\registers[357][0] ), .C(
        \registers[358][0] ), .D(\registers[359][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1420) );
  MX4X1 U4357 ( .A(\registers[276][0] ), .B(\registers[277][0] ), .C(
        \registers[278][0] ), .D(\registers[279][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1448) );
  MX4X1 U4358 ( .A(\registers[260][0] ), .B(\registers[261][0] ), .C(
        \registers[262][0] ), .D(\registers[263][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1453) );
  MX4X1 U4359 ( .A(\registers[308][0] ), .B(\registers[309][0] ), .C(
        \registers[310][0] ), .D(\registers[311][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1438) );
  MX4X1 U4360 ( .A(\registers[292][0] ), .B(\registers[293][0] ), .C(
        \registers[294][0] ), .D(\registers[295][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1443) );
  MX4X1 U4361 ( .A(\registers[468][0] ), .B(\registers[469][0] ), .C(
        \registers[470][0] ), .D(\registers[471][0] ), .S0(n4115), .S1(n4357), 
        .Y(n1381) );
  MX4X1 U4362 ( .A(\registers[452][0] ), .B(\registers[453][0] ), .C(
        \registers[454][0] ), .D(\registers[455][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1386) );
  MX4X1 U4363 ( .A(\registers[500][0] ), .B(\registers[501][0] ), .C(
        \registers[502][0] ), .D(\registers[503][0] ), .S0(n4115), .S1(n4356), 
        .Y(n1371) );
  MX4X1 U4364 ( .A(\registers[484][0] ), .B(\registers[485][0] ), .C(
        \registers[486][0] ), .D(\registers[487][0] ), .S0(n4115), .S1(n4356), 
        .Y(n1376) );
  MX4X1 U4365 ( .A(\registers[404][0] ), .B(\registers[405][0] ), .C(
        \registers[406][0] ), .D(\registers[407][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1404) );
  MX4X1 U4366 ( .A(\registers[388][0] ), .B(\registers[389][0] ), .C(
        \registers[390][0] ), .D(\registers[391][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1409) );
  MX4X1 U4367 ( .A(\registers[436][0] ), .B(\registers[437][0] ), .C(
        \registers[438][0] ), .D(\registers[439][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1392) );
  MX4X1 U4368 ( .A(\registers[420][0] ), .B(\registers[421][0] ), .C(
        \registers[422][0] ), .D(\registers[423][0] ), .S0(n4116), .S1(n4358), 
        .Y(n1397) );
  MX4X1 U4369 ( .A(\registers[84][0] ), .B(\registers[85][0] ), .C(
        \registers[86][0] ), .D(\registers[87][0] ), .S0(n4123), .S1(n4364), 
        .Y(n1516) );
  MX4X1 U4370 ( .A(\registers[68][0] ), .B(\registers[69][0] ), .C(
        \registers[70][0] ), .D(\registers[71][0] ), .S0(n4124), .S1(n4364), 
        .Y(n1521) );
  MX4X1 U4371 ( .A(\registers[116][0] ), .B(\registers[117][0] ), .C(
        \registers[118][0] ), .D(\registers[119][0] ), .S0(n4123), .S1(n4363), 
        .Y(n1506) );
  MX4X1 U4372 ( .A(\registers[100][0] ), .B(\registers[101][0] ), .C(
        \registers[102][0] ), .D(\registers[103][0] ), .S0(n4123), .S1(n4364), 
        .Y(n1511) );
  MX4X1 U4373 ( .A(\registers[20][0] ), .B(\registers[21][0] ), .C(
        \registers[22][0] ), .D(\registers[23][0] ), .S0(n4125), .S1(n4365), 
        .Y(n1538) );
  MX4X1 U4374 ( .A(\registers[4][0] ), .B(\registers[5][0] ), .C(
        \registers[6][0] ), .D(\registers[7][0] ), .S0(n4125), .S1(n4366), .Y(
        n1544) );
  MX4X1 U4375 ( .A(\registers[52][0] ), .B(\registers[53][0] ), .C(
        \registers[54][0] ), .D(\registers[55][0] ), .S0(n4124), .S1(n4365), 
        .Y(n1527) );
  MX4X1 U4376 ( .A(\registers[36][0] ), .B(\registers[37][0] ), .C(
        \registers[38][0] ), .D(\registers[39][0] ), .S0(n4124), .S1(n4365), 
        .Y(n1532) );
  MX4X1 U4377 ( .A(\registers[212][0] ), .B(\registers[213][0] ), .C(
        \registers[214][0] ), .D(\registers[215][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1472) );
  MX4X1 U4378 ( .A(\registers[196][0] ), .B(\registers[197][0] ), .C(
        \registers[198][0] ), .D(\registers[199][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1477) );
  MX4X1 U4379 ( .A(\registers[244][0] ), .B(\registers[245][0] ), .C(
        \registers[246][0] ), .D(\registers[247][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1460) );
  MX4X1 U4380 ( .A(\registers[228][0] ), .B(\registers[229][0] ), .C(
        \registers[230][0] ), .D(\registers[231][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1465) );
  MX4X1 U4381 ( .A(\registers[148][0] ), .B(\registers[149][0] ), .C(
        \registers[150][0] ), .D(\registers[151][0] ), .S0(n4122), .S1(n4363), 
        .Y(n1493) );
  MX4X1 U4382 ( .A(\registers[132][0] ), .B(\registers[133][0] ), .C(
        \registers[134][0] ), .D(\registers[135][0] ), .S0(n4122), .S1(n4363), 
        .Y(n1498) );
  MX4X1 U4383 ( .A(\registers[180][0] ), .B(\registers[181][0] ), .C(
        \registers[182][0] ), .D(\registers[183][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1483) );
  MX4X1 U4384 ( .A(\registers[164][0] ), .B(\registers[165][0] ), .C(
        \registers[166][0] ), .D(\registers[167][0] ), .S0(n4122), .S1(n4362), 
        .Y(n1488) );
  MX4X1 U4385 ( .A(\registers[852][0] ), .B(\registers[853][0] ), .C(
        \registers[854][0] ), .D(\registers[855][0] ), .S0(n4107), .S1(n4458), 
        .Y(n1099) );
  MX4X1 U4386 ( .A(\registers[836][0] ), .B(\registers[837][0] ), .C(
        \registers[838][0] ), .D(\registers[839][0] ), .S0(n4108), .S1(n4465), 
        .Y(n1104) );
  MX4X1 U4387 ( .A(\registers[884][0] ), .B(\registers[885][0] ), .C(
        \registers[886][0] ), .D(\registers[887][0] ), .S0(n4107), .S1(n4457), 
        .Y(n1089) );
  MX4X1 U4388 ( .A(\registers[868][0] ), .B(\registers[869][0] ), .C(
        \registers[870][0] ), .D(\registers[871][0] ), .S0(n4107), .S1(n4496), 
        .Y(n1094) );
  MX4X1 U4389 ( .A(\registers[788][0] ), .B(\registers[789][0] ), .C(
        \registers[790][0] ), .D(\registers[791][0] ), .S0(n4109), .S1(n4467), 
        .Y(n1162) );
  MX4X1 U4390 ( .A(\registers[772][0] ), .B(\registers[773][0] ), .C(
        \registers[774][0] ), .D(\registers[775][0] ), .S0(n4109), .S1(n4351), 
        .Y(n1167) );
  MX4X1 U4391 ( .A(\registers[820][0] ), .B(\registers[821][0] ), .C(
        \registers[822][0] ), .D(\registers[823][0] ), .S0(n4108), .S1(n4477), 
        .Y(n1152) );
  MX4X1 U4392 ( .A(\registers[804][0] ), .B(\registers[805][0] ), .C(
        \registers[806][0] ), .D(\registers[807][0] ), .S0(n4108), .S1(n4444), 
        .Y(n1157) );
  MX4X1 U4393 ( .A(\registers[980][0] ), .B(\registers[981][0] ), .C(
        \registers[982][0] ), .D(\registers[983][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1057) );
  MX4X1 U4394 ( .A(\registers[964][0] ), .B(\registers[965][0] ), .C(
        \registers[966][0] ), .D(\registers[967][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1062) );
  MX4X1 U4395 ( .A(\registers[916][0] ), .B(\registers[917][0] ), .C(
        \registers[918][0] ), .D(\registers[919][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1078) );
  MX4X1 U4396 ( .A(\registers[900][0] ), .B(\registers[901][0] ), .C(
        \registers[902][0] ), .D(\registers[903][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1083) );
  MX4X1 U4397 ( .A(\registers[948][0] ), .B(\registers[949][0] ), .C(
        \registers[950][0] ), .D(\registers[951][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1068) );
  MX4X1 U4398 ( .A(\registers[932][0] ), .B(\registers[933][0] ), .C(
        \registers[934][0] ), .D(\registers[935][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1073) );
  MX4X1 U4399 ( .A(\registers[596][0] ), .B(\registers[597][0] ), .C(
        \registers[598][0] ), .D(\registers[599][0] ), .S0(n4113), .S1(n4354), 
        .Y(n1335) );
  MX4X1 U4400 ( .A(\registers[580][0] ), .B(\registers[581][0] ), .C(
        \registers[582][0] ), .D(\registers[583][0] ), .S0(n4113), .S1(n4354), 
        .Y(n1340) );
  MX4X1 U4401 ( .A(\registers[628][0] ), .B(\registers[629][0] ), .C(
        \registers[630][0] ), .D(\registers[631][0] ), .S0(n4112), .S1(n4354), 
        .Y(n1315) );
  MX4X1 U4402 ( .A(\registers[612][0] ), .B(\registers[613][0] ), .C(
        \registers[614][0] ), .D(\registers[615][0] ), .S0(n4112), .S1(n4354), 
        .Y(n1325) );
  MX4X1 U4403 ( .A(\registers[532][0] ), .B(\registers[533][0] ), .C(
        \registers[534][0] ), .D(\registers[535][0] ), .S0(n4114), .S1(n4355), 
        .Y(n1356) );
  MX4X1 U4404 ( .A(\registers[516][0] ), .B(\registers[517][0] ), .C(
        \registers[518][0] ), .D(\registers[519][0] ), .S0(n4114), .S1(n4356), 
        .Y(n1361) );
  MX4X1 U4405 ( .A(\registers[564][0] ), .B(\registers[565][0] ), .C(
        \registers[566][0] ), .D(\registers[567][0] ), .S0(n4113), .S1(n4355), 
        .Y(n1346) );
  MX4X1 U4406 ( .A(\registers[548][0] ), .B(\registers[549][0] ), .C(
        \registers[550][0] ), .D(\registers[551][0] ), .S0(n4114), .S1(n4355), 
        .Y(n1351) );
  MX4X1 U4407 ( .A(\registers[724][0] ), .B(\registers[725][0] ), .C(
        \registers[726][0] ), .D(\registers[727][0] ), .S0(n4110), .S1(n4352), 
        .Y(n1184) );
  MX4X1 U4408 ( .A(\registers[708][0] ), .B(\registers[709][0] ), .C(
        \registers[710][0] ), .D(\registers[711][0] ), .S0(n4110), .S1(n4352), 
        .Y(n1204) );
  MX4X1 U4409 ( .A(\registers[756][0] ), .B(\registers[757][0] ), .C(
        \registers[758][0] ), .D(\registers[759][0] ), .S0(n4109), .S1(n4351), 
        .Y(n1174) );
  MX4X1 U4410 ( .A(\registers[740][0] ), .B(\registers[741][0] ), .C(
        \registers[742][0] ), .D(\registers[743][0] ), .S0(n4110), .S1(n4351), 
        .Y(n1179) );
  MX4X1 U4411 ( .A(\registers[660][0] ), .B(\registers[661][0] ), .C(
        \registers[662][0] ), .D(\registers[663][0] ), .S0(n4111), .S1(n4353), 
        .Y(n1293) );
  MX4X1 U4412 ( .A(\registers[644][0] ), .B(\registers[645][0] ), .C(
        \registers[646][0] ), .D(\registers[647][0] ), .S0(n4112), .S1(n4353), 
        .Y(n1303) );
  MX4X1 U4413 ( .A(\registers[692][0] ), .B(\registers[693][0] ), .C(
        \registers[694][0] ), .D(\registers[695][0] ), .S0(n4111), .S1(n4352), 
        .Y(n1273) );
  MX4X1 U4414 ( .A(\registers[676][0] ), .B(\registers[677][0] ), .C(
        \registers[678][0] ), .D(\registers[679][0] ), .S0(n4111), .S1(n4353), 
        .Y(n1283) );
  MX4X1 U4415 ( .A(\registers[340][1] ), .B(\registers[341][1] ), .C(
        \registers[342][1] ), .D(\registers[343][1] ), .S0(n4139), .S1(n4379), 
        .Y(n1783) );
  MX4X1 U4416 ( .A(\registers[324][1] ), .B(\registers[325][1] ), .C(
        \registers[326][1] ), .D(\registers[327][1] ), .S0(n4140), .S1(n4379), 
        .Y(n1788) );
  MX4X1 U4417 ( .A(\registers[372][1] ), .B(\registers[373][1] ), .C(
        \registers[374][1] ), .D(\registers[375][1] ), .S0(n4139), .S1(n4378), 
        .Y(n1772) );
  MX4X1 U4418 ( .A(\registers[356][1] ), .B(\registers[357][1] ), .C(
        \registers[358][1] ), .D(\registers[359][1] ), .S0(n4139), .S1(n4378), 
        .Y(n1778) );
  MX4X1 U4419 ( .A(\registers[276][1] ), .B(\registers[277][1] ), .C(
        \registers[278][1] ), .D(\registers[279][1] ), .S0(n4141), .S1(n4380), 
        .Y(n1804) );
  MX4X1 U4420 ( .A(\registers[260][1] ), .B(\registers[261][1] ), .C(
        \registers[262][1] ), .D(\registers[263][1] ), .S0(n4141), .S1(n4380), 
        .Y(n1810) );
  MX4X1 U4421 ( .A(\registers[308][1] ), .B(\registers[309][1] ), .C(
        \registers[310][1] ), .D(\registers[311][1] ), .S0(n4140), .S1(n4379), 
        .Y(n1794) );
  MX4X1 U4422 ( .A(\registers[292][1] ), .B(\registers[293][1] ), .C(
        \registers[294][1] ), .D(\registers[295][1] ), .S0(n4140), .S1(n4380), 
        .Y(n1799) );
  MX4X1 U4423 ( .A(\registers[468][1] ), .B(\registers[469][1] ), .C(
        \registers[470][1] ), .D(\registers[471][1] ), .S0(n4137), .S1(n4376), 
        .Y(n1739) );
  MX4X1 U4424 ( .A(\registers[452][1] ), .B(\registers[453][1] ), .C(
        \registers[454][1] ), .D(\registers[455][1] ), .S0(n4137), .S1(n4377), 
        .Y(n1745) );
  MX4X1 U4425 ( .A(\registers[500][1] ), .B(\registers[501][1] ), .C(
        \registers[502][1] ), .D(\registers[503][1] ), .S0(n4136), .S1(n4376), 
        .Y(n1729) );
  MX4X1 U4426 ( .A(\registers[484][1] ), .B(\registers[485][1] ), .C(
        \registers[486][1] ), .D(\registers[487][1] ), .S0(n4136), .S1(n4376), 
        .Y(n1734) );
  MX4X1 U4427 ( .A(\registers[404][1] ), .B(\registers[405][1] ), .C(
        \registers[406][1] ), .D(\registers[407][1] ), .S0(n4138), .S1(n4378), 
        .Y(n1761) );
  MX4X1 U4428 ( .A(\registers[388][1] ), .B(\registers[389][1] ), .C(
        \registers[390][1] ), .D(\registers[391][1] ), .S0(n4138), .S1(n4378), 
        .Y(n1766) );
  MX4X1 U4429 ( .A(\registers[436][1] ), .B(\registers[437][1] ), .C(
        \registers[438][1] ), .D(\registers[439][1] ), .S0(n4137), .S1(n4377), 
        .Y(n1751) );
  MX4X1 U4430 ( .A(\registers[420][1] ), .B(\registers[421][1] ), .C(
        \registers[422][1] ), .D(\registers[423][1] ), .S0(n4138), .S1(n4377), 
        .Y(n1756) );
  MX4X1 U4431 ( .A(\registers[84][1] ), .B(\registers[85][1] ), .C(
        \registers[86][1] ), .D(\registers[87][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1870) );
  MX4X1 U4432 ( .A(\registers[68][1] ), .B(\registers[69][1] ), .C(
        \registers[70][1] ), .D(\registers[71][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1877) );
  MX4X1 U4433 ( .A(\registers[116][1] ), .B(\registers[117][1] ), .C(
        \registers[118][1] ), .D(\registers[119][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1860) );
  MX4X1 U4434 ( .A(\registers[100][1] ), .B(\registers[101][1] ), .C(
        \registers[102][1] ), .D(\registers[103][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1865) );
  MX4X1 U4435 ( .A(\registers[20][1] ), .B(\registers[21][1] ), .C(
        \registers[22][1] ), .D(\registers[23][1] ), .S0(n4146), .S1(n4385), 
        .Y(n1893) );
  MX4X1 U4436 ( .A(\registers[4][1] ), .B(\registers[5][1] ), .C(
        \registers[6][1] ), .D(\registers[7][1] ), .S0(n4146), .S1(n4385), .Y(
        n1898) );
  MX4X1 U4437 ( .A(\registers[52][1] ), .B(\registers[53][1] ), .C(
        \registers[54][1] ), .D(\registers[55][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1883) );
  MX4X1 U4438 ( .A(\registers[36][1] ), .B(\registers[37][1] ), .C(
        \registers[38][1] ), .D(\registers[39][1] ), .S0(n4146), .S1(n4385), 
        .Y(n1888) );
  MX4X1 U4439 ( .A(\registers[212][1] ), .B(\registers[213][1] ), .C(
        \registers[214][1] ), .D(\registers[215][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1827) );
  MX4X1 U4440 ( .A(\registers[196][1] ), .B(\registers[197][1] ), .C(
        \registers[198][1] ), .D(\registers[199][1] ), .S0(n4142), .S1(n4382), 
        .Y(n1832) );
  MX4X1 U4441 ( .A(\registers[244][1] ), .B(\registers[245][1] ), .C(
        \registers[246][1] ), .D(\registers[247][1] ), .S0(n4141), .S1(n4381), 
        .Y(n1817) );
  MX4X1 U4442 ( .A(\registers[228][1] ), .B(\registers[229][1] ), .C(
        \registers[230][1] ), .D(\registers[231][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1822) );
  MX4X1 U4443 ( .A(\registers[148][1] ), .B(\registers[149][1] ), .C(
        \registers[150][1] ), .D(\registers[151][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1849) );
  MX4X1 U4444 ( .A(\registers[132][1] ), .B(\registers[133][1] ), .C(
        \registers[134][1] ), .D(\registers[135][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1854) );
  MX4X1 U4445 ( .A(\registers[180][1] ), .B(\registers[181][1] ), .C(
        \registers[182][1] ), .D(\registers[183][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1838) );
  MX4X1 U4446 ( .A(\registers[164][1] ), .B(\registers[165][1] ), .C(
        \registers[166][1] ), .D(\registers[167][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1844) );
  MX4X1 U4447 ( .A(\registers[852][1] ), .B(\registers[853][1] ), .C(
        \registers[854][1] ), .D(\registers[855][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1607) );
  MX4X1 U4448 ( .A(\registers[836][1] ), .B(\registers[837][1] ), .C(
        \registers[838][1] ), .D(\registers[839][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1613) );
  MX4X1 U4449 ( .A(\registers[884][1] ), .B(\registers[885][1] ), .C(
        \registers[886][1] ), .D(\registers[887][1] ), .S0(n4128), .S1(n4368), 
        .Y(n1595) );
  MX4X1 U4450 ( .A(\registers[868][1] ), .B(\registers[869][1] ), .C(
        \registers[870][1] ), .D(\registers[871][1] ), .S0(n4128), .S1(n4369), 
        .Y(n1600) );
  MX4X1 U4451 ( .A(\registers[788][1] ), .B(\registers[789][1] ), .C(
        \registers[790][1] ), .D(\registers[791][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1629) );
  MX4X1 U4452 ( .A(\registers[772][1] ), .B(\registers[773][1] ), .C(
        \registers[774][1] ), .D(\registers[775][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1634) );
  MX4X1 U4453 ( .A(\registers[820][1] ), .B(\registers[821][1] ), .C(
        \registers[822][1] ), .D(\registers[823][1] ), .S0(n4129), .S1(n4370), 
        .Y(n1619) );
  MX4X1 U4454 ( .A(\registers[804][1] ), .B(\registers[805][1] ), .C(
        \registers[806][1] ), .D(\registers[807][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1624) );
  MX4X1 U4455 ( .A(\registers[980][1] ), .B(\registers[981][1] ), .C(
        \registers[982][1] ), .D(\registers[983][1] ), .S0(n4126), .S1(n4366), 
        .Y(n1561) );
  MX4X1 U4456 ( .A(\registers[964][1] ), .B(\registers[965][1] ), .C(
        \registers[966][1] ), .D(\registers[967][1] ), .S0(n4126), .S1(n4367), 
        .Y(n1566) );
  MX4X1 U4457 ( .A(\registers[1012][1] ), .B(\registers[1013][1] ), .C(
        \registers[1014][1] ), .D(\registers[1015][1] ), .S0(n4125), .S1(n4366), .Y(n1551) );
  MX4X1 U4458 ( .A(\registers[996][1] ), .B(\registers[997][1] ), .C(
        \registers[998][1] ), .D(\registers[999][1] ), .S0(n4126), .S1(n4366), 
        .Y(n1556) );
  MX4X1 U4459 ( .A(\registers[916][1] ), .B(\registers[917][1] ), .C(
        \registers[918][1] ), .D(\registers[919][1] ), .S0(n4127), .S1(n4368), 
        .Y(n1584) );
  MX4X1 U4460 ( .A(\registers[900][1] ), .B(\registers[901][1] ), .C(
        \registers[902][1] ), .D(\registers[903][1] ), .S0(n4128), .S1(n4368), 
        .Y(n1589) );
  MX4X1 U4461 ( .A(\registers[948][1] ), .B(\registers[949][1] ), .C(
        \registers[950][1] ), .D(\registers[951][1] ), .S0(n4127), .S1(n4367), 
        .Y(n1574) );
  MX4X1 U4462 ( .A(\registers[932][1] ), .B(\registers[933][1] ), .C(
        \registers[934][1] ), .D(\registers[935][1] ), .S0(n4127), .S1(n4367), 
        .Y(n1579) );
  MX4X1 U4463 ( .A(\registers[596][1] ), .B(\registers[597][1] ), .C(
        \registers[598][1] ), .D(\registers[599][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1695) );
  MX4X1 U4464 ( .A(\registers[580][1] ), .B(\registers[581][1] ), .C(
        \registers[582][1] ), .D(\registers[583][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1700) );
  MX4X1 U4465 ( .A(\registers[628][1] ), .B(\registers[629][1] ), .C(
        \registers[630][1] ), .D(\registers[631][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1685) );
  MX4X1 U4466 ( .A(\registers[612][1] ), .B(\registers[613][1] ), .C(
        \registers[614][1] ), .D(\registers[615][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1690) );
  MX4X1 U4467 ( .A(\registers[532][1] ), .B(\registers[533][1] ), .C(
        \registers[534][1] ), .D(\registers[535][1] ), .S0(n4135), .S1(n4375), 
        .Y(n1717) );
  MX4X1 U4468 ( .A(\registers[516][1] ), .B(\registers[517][1] ), .C(
        \registers[518][1] ), .D(\registers[519][1] ), .S0(n4136), .S1(n4375), 
        .Y(n1722) );
  MX4X1 U4469 ( .A(\registers[564][1] ), .B(\registers[565][1] ), .C(
        \registers[566][1] ), .D(\registers[567][1] ), .S0(n4135), .S1(n4374), 
        .Y(n1706) );
  MX4X1 U4470 ( .A(\registers[548][1] ), .B(\registers[549][1] ), .C(
        \registers[550][1] ), .D(\registers[551][1] ), .S0(n4135), .S1(n4375), 
        .Y(n1712) );
  MX4X1 U4471 ( .A(\registers[724][1] ), .B(\registers[725][1] ), .C(
        \registers[726][1] ), .D(\registers[727][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1652) );
  MX4X1 U4472 ( .A(\registers[708][1] ), .B(\registers[709][1] ), .C(
        \registers[710][1] ), .D(\registers[711][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1657) );
  MX4X1 U4473 ( .A(\registers[756][1] ), .B(\registers[757][1] ), .C(
        \registers[758][1] ), .D(\registers[759][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1642) );
  MX4X1 U4474 ( .A(\registers[740][1] ), .B(\registers[741][1] ), .C(
        \registers[742][1] ), .D(\registers[743][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1647) );
  MX4X1 U4475 ( .A(\registers[660][1] ), .B(\registers[661][1] ), .C(
        \registers[662][1] ), .D(\registers[663][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1673) );
  MX4X1 U4476 ( .A(\registers[644][1] ), .B(\registers[645][1] ), .C(
        \registers[646][1] ), .D(\registers[647][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1679) );
  MX4X1 U4477 ( .A(\registers[692][1] ), .B(\registers[693][1] ), .C(
        \registers[694][1] ), .D(\registers[695][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1663) );
  MX4X1 U4478 ( .A(\registers[676][1] ), .B(\registers[677][1] ), .C(
        \registers[678][1] ), .D(\registers[679][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1668) );
  MX4X1 U4479 ( .A(\registers[340][2] ), .B(\registers[341][2] ), .C(
        \registers[342][2] ), .D(\registers[343][2] ), .S0(n4161), .S1(n4398), 
        .Y(n2134) );
  MX4X1 U4480 ( .A(\registers[324][2] ), .B(\registers[325][2] ), .C(
        \registers[326][2] ), .D(\registers[327][2] ), .S0(n4161), .S1(n4399), 
        .Y(n2141) );
  MX4X1 U4481 ( .A(\registers[372][2] ), .B(\registers[373][2] ), .C(
        \registers[374][2] ), .D(\registers[375][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2124) );
  MX4X1 U4482 ( .A(\registers[356][2] ), .B(\registers[357][2] ), .C(
        \registers[358][2] ), .D(\registers[359][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2129) );
  MX4X1 U4483 ( .A(\registers[276][2] ), .B(\registers[277][2] ), .C(
        \registers[278][2] ), .D(\registers[279][2] ), .S0(n4162), .S1(n4400), 
        .Y(n2157) );
  MX4X1 U4484 ( .A(\registers[260][2] ), .B(\registers[261][2] ), .C(
        \registers[262][2] ), .D(\registers[263][2] ), .S0(n4162), .S1(n4400), 
        .Y(n2162) );
  MX4X1 U4485 ( .A(\registers[308][2] ), .B(\registers[309][2] ), .C(
        \registers[310][2] ), .D(\registers[311][2] ), .S0(n4161), .S1(n4399), 
        .Y(n2147) );
  MX4X1 U4486 ( .A(\registers[292][2] ), .B(\registers[293][2] ), .C(
        \registers[294][2] ), .D(\registers[295][2] ), .S0(n4162), .S1(n4399), 
        .Y(n2152) );
  MX4X1 U4487 ( .A(\registers[468][2] ), .B(\registers[469][2] ), .C(
        \registers[470][2] ), .D(\registers[471][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2091) );
  MX4X1 U4488 ( .A(\registers[452][2] ), .B(\registers[453][2] ), .C(
        \registers[454][2] ), .D(\registers[455][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2096) );
  MX4X1 U4489 ( .A(\registers[500][2] ), .B(\registers[501][2] ), .C(
        \registers[502][2] ), .D(\registers[503][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2081) );
  MX4X1 U4490 ( .A(\registers[484][2] ), .B(\registers[485][2] ), .C(
        \registers[486][2] ), .D(\registers[487][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2086) );
  MX4X1 U4491 ( .A(\registers[404][2] ), .B(\registers[405][2] ), .C(
        \registers[406][2] ), .D(\registers[407][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2113) );
  MX4X1 U4492 ( .A(\registers[388][2] ), .B(\registers[389][2] ), .C(
        \registers[390][2] ), .D(\registers[391][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2118) );
  MX4X1 U4493 ( .A(\registers[436][2] ), .B(\registers[437][2] ), .C(
        \registers[438][2] ), .D(\registers[439][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2102) );
  MX4X1 U4494 ( .A(\registers[420][2] ), .B(\registers[421][2] ), .C(
        \registers[422][2] ), .D(\registers[423][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2108) );
  MX4X1 U4495 ( .A(\registers[84][2] ), .B(\registers[85][2] ), .C(
        \registers[86][2] ), .D(\registers[87][2] ), .S0(n4166), .S1(n4403), 
        .Y(n2223) );
  MX4X1 U4496 ( .A(\registers[68][2] ), .B(\registers[69][2] ), .C(
        \registers[70][2] ), .D(\registers[71][2] ), .S0(n4166), .S1(n4404), 
        .Y(n2228) );
  MX4X1 U4497 ( .A(\registers[116][2] ), .B(\registers[117][2] ), .C(
        \registers[118][2] ), .D(\registers[119][2] ), .S0(n4165), .S1(n4403), 
        .Y(n2213) );
  MX4X1 U4498 ( .A(\registers[100][2] ), .B(\registers[101][2] ), .C(
        \registers[102][2] ), .D(\registers[103][2] ), .S0(n4166), .S1(n4403), 
        .Y(n2218) );
  MX4X1 U4499 ( .A(\registers[20][2] ), .B(\registers[21][2] ), .C(
        \registers[22][2] ), .D(\registers[23][2] ), .S0(n4167), .S1(n4405), 
        .Y(n2245) );
  MX4X1 U4500 ( .A(\registers[4][2] ), .B(\registers[5][2] ), .C(
        \registers[6][2] ), .D(\registers[7][2] ), .S0(n4168), .S1(n4405), .Y(
        n2250) );
  MX4X1 U4501 ( .A(\registers[52][2] ), .B(\registers[53][2] ), .C(
        \registers[54][2] ), .D(\registers[55][2] ), .S0(n4167), .S1(n4404), 
        .Y(n2234) );
  MX4X1 U4502 ( .A(\registers[36][2] ), .B(\registers[37][2] ), .C(
        \registers[38][2] ), .D(\registers[39][2] ), .S0(n4167), .S1(n4404), 
        .Y(n2240) );
  MX4X1 U4503 ( .A(\registers[212][2] ), .B(\registers[213][2] ), .C(
        \registers[214][2] ), .D(\registers[215][2] ), .S0(n4163), .S1(n4401), 
        .Y(n2180) );
  MX4X1 U4504 ( .A(\registers[196][2] ), .B(\registers[197][2] ), .C(
        \registers[198][2] ), .D(\registers[199][2] ), .S0(n4164), .S1(n4401), 
        .Y(n2185) );
  MX4X1 U4505 ( .A(\registers[244][2] ), .B(\registers[245][2] ), .C(
        \registers[246][2] ), .D(\registers[247][2] ), .S0(n4163), .S1(n4400), 
        .Y(n2169) );
  MX4X1 U4506 ( .A(\registers[228][2] ), .B(\registers[229][2] ), .C(
        \registers[230][2] ), .D(\registers[231][2] ), .S0(n4163), .S1(n4401), 
        .Y(n2175) );
  MX4X1 U4507 ( .A(\registers[148][2] ), .B(\registers[149][2] ), .C(
        \registers[150][2] ), .D(\registers[151][2] ), .S0(n4165), .S1(n4402), 
        .Y(n2201) );
  MX4X1 U4508 ( .A(\registers[132][2] ), .B(\registers[133][2] ), .C(
        \registers[134][2] ), .D(\registers[135][2] ), .S0(n4165), .S1(n4402), 
        .Y(n2207) );
  MX4X1 U4509 ( .A(\registers[180][2] ), .B(\registers[181][2] ), .C(
        \registers[182][2] ), .D(\registers[183][2] ), .S0(n4164), .S1(n4402), 
        .Y(n2191) );
  MX4X1 U4510 ( .A(\registers[164][2] ), .B(\registers[165][2] ), .C(
        \registers[166][2] ), .D(\registers[167][2] ), .S0(n4164), .S1(n4402), 
        .Y(n2196) );
  MX4X1 U4511 ( .A(\registers[852][2] ), .B(\registers[853][2] ), .C(
        \registers[854][2] ), .D(\registers[855][2] ), .S0(n4150), .S1(n4389), 
        .Y(n1959) );
  MX4X1 U4512 ( .A(\registers[836][2] ), .B(\registers[837][2] ), .C(
        \registers[838][2] ), .D(\registers[839][2] ), .S0(n4150), .S1(n4389), 
        .Y(n1964) );
  MX4X1 U4513 ( .A(\registers[884][2] ), .B(\registers[885][2] ), .C(
        \registers[886][2] ), .D(\registers[887][2] ), .S0(n4149), .S1(n4388), 
        .Y(n1949) );
  MX4X1 U4514 ( .A(\registers[868][2] ), .B(\registers[869][2] ), .C(
        \registers[870][2] ), .D(\registers[871][2] ), .S0(n4150), .S1(n4388), 
        .Y(n1954) );
  MX4X1 U4515 ( .A(\registers[788][2] ), .B(\registers[789][2] ), .C(
        \registers[790][2] ), .D(\registers[791][2] ), .S0(n4151), .S1(n4390), 
        .Y(n1981) );
  MX4X1 U4516 ( .A(\registers[772][2] ), .B(\registers[773][2] ), .C(
        \registers[774][2] ), .D(\registers[775][2] ), .S0(n4152), .S1(n4390), 
        .Y(n1986) );
  MX4X1 U4517 ( .A(\registers[820][2] ), .B(\registers[821][2] ), .C(
        \registers[822][2] ), .D(\registers[823][2] ), .S0(n4151), .S1(n4389), 
        .Y(n1970) );
  MX4X1 U4518 ( .A(\registers[804][2] ), .B(\registers[805][2] ), .C(
        \registers[806][2] ), .D(\registers[807][2] ), .S0(n4151), .S1(n4390), 
        .Y(n1976) );
  MX4X1 U4519 ( .A(\registers[980][2] ), .B(\registers[981][2] ), .C(
        \registers[982][2] ), .D(\registers[983][2] ), .S0(n4147), .S1(n4386), 
        .Y(n1916) );
  MX4X1 U4520 ( .A(\registers[964][2] ), .B(\registers[965][2] ), .C(
        \registers[966][2] ), .D(\registers[967][2] ), .S0(n4148), .S1(n4386), 
        .Y(n1921) );
  MX4X1 U4521 ( .A(\registers[1012][2] ), .B(\registers[1013][2] ), .C(
        \registers[1014][2] ), .D(\registers[1015][2] ), .S0(n4147), .S1(n4386), .Y(n1905) );
  MX4X1 U4522 ( .A(\registers[996][2] ), .B(\registers[997][2] ), .C(
        \registers[998][2] ), .D(\registers[999][2] ), .S0(n4147), .S1(n4386), 
        .Y(n1911) );
  MX4X1 U4523 ( .A(\registers[916][2] ), .B(\registers[917][2] ), .C(
        \registers[918][2] ), .D(\registers[919][2] ), .S0(n4149), .S1(n4387), 
        .Y(n1937) );
  MX4X1 U4524 ( .A(\registers[900][2] ), .B(\registers[901][2] ), .C(
        \registers[902][2] ), .D(\registers[903][2] ), .S0(n4149), .S1(n4388), 
        .Y(n1943) );
  MX4X1 U4525 ( .A(\registers[948][2] ), .B(\registers[949][2] ), .C(
        \registers[950][2] ), .D(\registers[951][2] ), .S0(n4148), .S1(n4387), 
        .Y(n1927) );
  MX4X1 U4526 ( .A(\registers[932][2] ), .B(\registers[933][2] ), .C(
        \registers[934][2] ), .D(\registers[935][2] ), .S0(n4148), .S1(n4387), 
        .Y(n1932) );
  MX4X1 U4527 ( .A(\registers[596][2] ), .B(\registers[597][2] ), .C(
        \registers[598][2] ), .D(\registers[599][2] ), .S0(n4155), .S1(n4394), 
        .Y(n2047) );
  MX4X1 U4528 ( .A(\registers[580][2] ), .B(\registers[581][2] ), .C(
        \registers[582][2] ), .D(\registers[583][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2052) );
  MX4X1 U4529 ( .A(\registers[628][2] ), .B(\registers[629][2] ), .C(
        \registers[630][2] ), .D(\registers[631][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2036) );
  MX4X1 U4530 ( .A(\registers[612][2] ), .B(\registers[613][2] ), .C(
        \registers[614][2] ), .D(\registers[615][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2042) );
  MX4X1 U4531 ( .A(\registers[532][2] ), .B(\registers[533][2] ), .C(
        \registers[534][2] ), .D(\registers[535][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2068) );
  MX4X1 U4532 ( .A(\registers[516][2] ), .B(\registers[517][2] ), .C(
        \registers[518][2] ), .D(\registers[519][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2074) );
  MX4X1 U4533 ( .A(\registers[564][2] ), .B(\registers[565][2] ), .C(
        \registers[566][2] ), .D(\registers[567][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2058) );
  MX4X1 U4534 ( .A(\registers[548][2] ), .B(\registers[549][2] ), .C(
        \registers[550][2] ), .D(\registers[551][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2063) );
  MX4X1 U4535 ( .A(\registers[724][2] ), .B(\registers[725][2] ), .C(
        \registers[726][2] ), .D(\registers[727][2] ), .S0(n4153), .S1(n4391), 
        .Y(n2003) );
  MX4X1 U4536 ( .A(\registers[708][2] ), .B(\registers[709][2] ), .C(
        \registers[710][2] ), .D(\registers[711][2] ), .S0(n4153), .S1(n4391), 
        .Y(n2009) );
  MX4X1 U4537 ( .A(\registers[756][2] ), .B(\registers[757][2] ), .C(
        \registers[758][2] ), .D(\registers[759][2] ), .S0(n4152), .S1(n4390), 
        .Y(n1993) );
  MX4X1 U4538 ( .A(\registers[740][2] ), .B(\registers[741][2] ), .C(
        \registers[742][2] ), .D(\registers[743][2] ), .S0(n4152), .S1(n4391), 
        .Y(n1998) );
  MX4X1 U4539 ( .A(\registers[660][2] ), .B(\registers[661][2] ), .C(
        \registers[662][2] ), .D(\registers[663][2] ), .S0(n4154), .S1(n4392), 
        .Y(n2025) );
  MX4X1 U4540 ( .A(\registers[644][2] ), .B(\registers[645][2] ), .C(
        \registers[646][2] ), .D(\registers[647][2] ), .S0(n4154), .S1(n4393), 
        .Y(n2030) );
  MX4X1 U4541 ( .A(\registers[692][2] ), .B(\registers[693][2] ), .C(
        \registers[694][2] ), .D(\registers[695][2] ), .S0(n4153), .S1(n4392), 
        .Y(n2015) );
  MX4X1 U4542 ( .A(\registers[676][2] ), .B(\registers[677][2] ), .C(
        \registers[678][2] ), .D(\registers[679][2] ), .S0(n4154), .S1(n4392), 
        .Y(n2020) );
  MX4X1 U4543 ( .A(\registers[340][3] ), .B(\registers[341][3] ), .C(
        \registers[342][3] ), .D(\registers[343][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2549) );
  MX4X1 U4544 ( .A(\registers[324][3] ), .B(\registers[325][3] ), .C(
        \registers[326][3] ), .D(\registers[327][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2554) );
  MX4X1 U4545 ( .A(\registers[372][3] ), .B(\registers[373][3] ), .C(
        \registers[374][3] ), .D(\registers[375][3] ), .S0(n4181), .S1(n4418), 
        .Y(n2539) );
  MX4X1 U4546 ( .A(\registers[356][3] ), .B(\registers[357][3] ), .C(
        \registers[358][3] ), .D(\registers[359][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2544) );
  MX4X1 U4547 ( .A(\registers[276][3] ), .B(\registers[277][3] ), .C(
        \registers[278][3] ), .D(\registers[279][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2570) );
  MX4X1 U4548 ( .A(\registers[260][3] ), .B(\registers[261][3] ), .C(
        \registers[262][3] ), .D(\registers[263][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2575) );
  MX4X1 U4549 ( .A(\registers[308][3] ), .B(\registers[309][3] ), .C(
        \registers[310][3] ), .D(\registers[311][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2560) );
  MX4X1 U4550 ( .A(\registers[292][3] ), .B(\registers[293][3] ), .C(
        \registers[294][3] ), .D(\registers[295][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2565) );
  MX4X1 U4551 ( .A(\registers[468][3] ), .B(\registers[469][3] ), .C(
        \registers[470][3] ), .D(\registers[471][3] ), .S0(n4179), .S1(n4416), 
        .Y(n2507) );
  MX4X1 U4552 ( .A(\registers[452][3] ), .B(\registers[453][3] ), .C(
        \registers[454][3] ), .D(\registers[455][3] ), .S0(n4180), .S1(n4416), 
        .Y(n2512) );
  MX4X1 U4553 ( .A(\registers[500][3] ), .B(\registers[501][3] ), .C(
        \registers[502][3] ), .D(\registers[503][3] ), .S0(n4179), .S1(n4415), 
        .Y(n2497) );
  MX4X1 U4554 ( .A(\registers[484][3] ), .B(\registers[485][3] ), .C(
        \registers[486][3] ), .D(\registers[487][3] ), .S0(n4179), .S1(n4415), 
        .Y(n2502) );
  MX4X1 U4555 ( .A(\registers[404][3] ), .B(\registers[405][3] ), .C(
        \registers[406][3] ), .D(\registers[407][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2528) );
  MX4X1 U4556 ( .A(\registers[388][3] ), .B(\registers[389][3] ), .C(
        \registers[390][3] ), .D(\registers[391][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2533) );
  MX4X1 U4557 ( .A(\registers[436][3] ), .B(\registers[437][3] ), .C(
        \registers[438][3] ), .D(\registers[439][3] ), .S0(n4180), .S1(n4416), 
        .Y(n2518) );
  MX4X1 U4558 ( .A(\registers[420][3] ), .B(\registers[421][3] ), .C(
        \registers[422][3] ), .D(\registers[423][3] ), .S0(n4180), .S1(n4417), 
        .Y(n2523) );
  MX4X1 U4559 ( .A(\registers[84][3] ), .B(\registers[85][3] ), .C(
        \registers[86][3] ), .D(\registers[87][3] ), .S0(n4187), .S1(n4423), 
        .Y(n2634) );
  MX4X1 U4560 ( .A(\registers[68][3] ), .B(\registers[69][3] ), .C(
        \registers[70][3] ), .D(\registers[71][3] ), .S0(n4188), .S1(n4423), 
        .Y(n2639) );
  MX4X1 U4561 ( .A(\registers[116][3] ), .B(\registers[117][3] ), .C(
        \registers[118][3] ), .D(\registers[119][3] ), .S0(n4187), .S1(n4422), 
        .Y(n2624) );
  MX4X1 U4562 ( .A(\registers[100][3] ), .B(\registers[101][3] ), .C(
        \registers[102][3] ), .D(\registers[103][3] ), .S0(n4187), .S1(n4423), 
        .Y(n2629) );
  MX4X1 U4563 ( .A(\registers[20][3] ), .B(\registers[21][3] ), .C(
        \registers[22][3] ), .D(\registers[23][3] ), .S0(n4189), .S1(n4424), 
        .Y(n2655) );
  MX4X1 U4564 ( .A(\registers[4][3] ), .B(\registers[5][3] ), .C(
        \registers[6][3] ), .D(\registers[7][3] ), .S0(n4189), .S1(n4425), .Y(
        n2660) );
  MX4X1 U4565 ( .A(\registers[52][3] ), .B(\registers[53][3] ), .C(
        \registers[54][3] ), .D(\registers[55][3] ), .S0(n4188), .S1(n4424), 
        .Y(n2645) );
  MX4X1 U4566 ( .A(\registers[36][3] ), .B(\registers[37][3] ), .C(
        \registers[38][3] ), .D(\registers[39][3] ), .S0(n4188), .S1(n4424), 
        .Y(n2650) );
  MX4X1 U4567 ( .A(\registers[212][3] ), .B(\registers[213][3] ), .C(
        \registers[214][3] ), .D(\registers[215][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2592) );
  MX4X1 U4568 ( .A(\registers[196][3] ), .B(\registers[197][3] ), .C(
        \registers[198][3] ), .D(\registers[199][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2597) );
  MX4X1 U4569 ( .A(\registers[244][3] ), .B(\registers[245][3] ), .C(
        \registers[246][3] ), .D(\registers[247][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2582) );
  MX4X1 U4570 ( .A(\registers[228][3] ), .B(\registers[229][3] ), .C(
        \registers[230][3] ), .D(\registers[231][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2587) );
  MX4X1 U4571 ( .A(\registers[148][3] ), .B(\registers[149][3] ), .C(
        \registers[150][3] ), .D(\registers[151][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2613) );
  MX4X1 U4572 ( .A(\registers[132][3] ), .B(\registers[133][3] ), .C(
        \registers[134][3] ), .D(\registers[135][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2618) );
  MX4X1 U4573 ( .A(\registers[180][3] ), .B(\registers[181][3] ), .C(
        \registers[182][3] ), .D(\registers[183][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2603) );
  MX4X1 U4574 ( .A(\registers[164][3] ), .B(\registers[165][3] ), .C(
        \registers[166][3] ), .D(\registers[167][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2608) );
  MX4X1 U4575 ( .A(\registers[852][3] ), .B(\registers[853][3] ), .C(
        \registers[854][3] ), .D(\registers[855][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2311) );
  MX4X1 U4576 ( .A(\registers[836][3] ), .B(\registers[837][3] ), .C(
        \registers[838][3] ), .D(\registers[839][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2316) );
  MX4X1 U4577 ( .A(\registers[884][3] ), .B(\registers[885][3] ), .C(
        \registers[886][3] ), .D(\registers[887][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2300) );
  MX4X1 U4578 ( .A(\registers[868][3] ), .B(\registers[869][3] ), .C(
        \registers[870][3] ), .D(\registers[871][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2306) );
  MX4X1 U4579 ( .A(\registers[788][3] ), .B(\registers[789][3] ), .C(
        \registers[790][3] ), .D(\registers[791][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2332) );
  MX4X1 U4580 ( .A(\registers[772][3] ), .B(\registers[773][3] ), .C(
        \registers[774][3] ), .D(\registers[775][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2341) );
  MX4X1 U4581 ( .A(\registers[820][3] ), .B(\registers[821][3] ), .C(
        \registers[822][3] ), .D(\registers[823][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2322) );
  MX4X1 U4582 ( .A(\registers[804][3] ), .B(\registers[805][3] ), .C(
        \registers[806][3] ), .D(\registers[807][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2327) );
  MX4X1 U4583 ( .A(\registers[980][3] ), .B(\registers[981][3] ), .C(
        \registers[982][3] ), .D(\registers[983][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2267) );
  MX4X1 U4584 ( .A(\registers[964][3] ), .B(\registers[965][3] ), .C(
        \registers[966][3] ), .D(\registers[967][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2273) );
  MX4X1 U4585 ( .A(\registers[1012][3] ), .B(\registers[1013][3] ), .C(
        \registers[1014][3] ), .D(\registers[1015][3] ), .S0(n4168), .S1(n4405), .Y(n2257) );
  MX4X1 U4586 ( .A(\registers[996][3] ), .B(\registers[997][3] ), .C(
        \registers[998][3] ), .D(\registers[999][3] ), .S0(n4168), .S1(n4406), 
        .Y(n2262) );
  MX4X1 U4587 ( .A(\registers[916][3] ), .B(\registers[917][3] ), .C(
        \registers[918][3] ), .D(\registers[919][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2289) );
  MX4X1 U4588 ( .A(\registers[900][3] ), .B(\registers[901][3] ), .C(
        \registers[902][3] ), .D(\registers[903][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2294) );
  MX4X1 U4589 ( .A(\registers[948][3] ), .B(\registers[949][3] ), .C(
        \registers[950][3] ), .D(\registers[951][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2279) );
  MX4X1 U4590 ( .A(\registers[932][3] ), .B(\registers[933][3] ), .C(
        \registers[934][3] ), .D(\registers[935][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2284) );
  MX4X1 U4591 ( .A(\registers[596][3] ), .B(\registers[597][3] ), .C(
        \registers[598][3] ), .D(\registers[599][3] ), .S0(n4177), .S1(n4413), 
        .Y(n2464) );
  MX4X1 U4592 ( .A(\registers[580][3] ), .B(\registers[581][3] ), .C(
        \registers[582][3] ), .D(\registers[583][3] ), .S0(n4177), .S1(n4414), 
        .Y(n2469) );
  MX4X1 U4593 ( .A(\registers[628][3] ), .B(\registers[629][3] ), .C(
        \registers[630][3] ), .D(\registers[631][3] ), .S0(n4176), .S1(n4413), 
        .Y(n2454) );
  MX4X1 U4594 ( .A(\registers[612][3] ), .B(\registers[613][3] ), .C(
        \registers[614][3] ), .D(\registers[615][3] ), .S0(n4176), .S1(n4413), 
        .Y(n2459) );
  MX4X1 U4595 ( .A(\registers[532][3] ), .B(\registers[533][3] ), .C(
        \registers[534][3] ), .D(\registers[535][3] ), .S0(n4178), .S1(n4414), 
        .Y(n2485) );
  MX4X1 U4596 ( .A(\registers[516][3] ), .B(\registers[517][3] ), .C(
        \registers[518][3] ), .D(\registers[519][3] ), .S0(n4178), .S1(n4415), 
        .Y(n2490) );
  MX4X1 U4597 ( .A(\registers[564][3] ), .B(\registers[565][3] ), .C(
        \registers[566][3] ), .D(\registers[567][3] ), .S0(n4177), .S1(n4414), 
        .Y(n2475) );
  MX4X1 U4598 ( .A(\registers[548][3] ), .B(\registers[549][3] ), .C(
        \registers[550][3] ), .D(\registers[551][3] ), .S0(n4178), .S1(n4414), 
        .Y(n2480) );
  MX4X1 U4599 ( .A(\registers[724][3] ), .B(\registers[725][3] ), .C(
        \registers[726][3] ), .D(\registers[727][3] ), .S0(n4174), .S1(n4411), 
        .Y(n2366) );
  MX4X1 U4600 ( .A(\registers[708][3] ), .B(\registers[709][3] ), .C(
        \registers[710][3] ), .D(\registers[711][3] ), .S0(n4174), .S1(n4411), 
        .Y(n2371) );
  MX4X1 U4601 ( .A(\registers[756][3] ), .B(\registers[757][3] ), .C(
        \registers[758][3] ), .D(\registers[759][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2355) );
  MX4X1 U4602 ( .A(\registers[740][3] ), .B(\registers[741][3] ), .C(
        \registers[742][3] ), .D(\registers[743][3] ), .S0(n4174), .S1(n4410), 
        .Y(n2360) );
  MX4X1 U4603 ( .A(\registers[660][3] ), .B(\registers[661][3] ), .C(
        \registers[662][3] ), .D(\registers[663][3] ), .S0(n4175), .S1(n4412), 
        .Y(n2443) );
  MX4X1 U4604 ( .A(\registers[644][3] ), .B(\registers[645][3] ), .C(
        \registers[646][3] ), .D(\registers[647][3] ), .S0(n4176), .S1(n4412), 
        .Y(n2448) );
  MX4X1 U4605 ( .A(\registers[692][3] ), .B(\registers[693][3] ), .C(
        \registers[694][3] ), .D(\registers[695][3] ), .S0(n4175), .S1(n4411), 
        .Y(n2378) );
  MX4X1 U4606 ( .A(\registers[676][3] ), .B(\registers[677][3] ), .C(
        \registers[678][3] ), .D(\registers[679][3] ), .S0(n4175), .S1(n4412), 
        .Y(n2438) );
  MX4X1 U4607 ( .A(\registers[340][4] ), .B(\registers[341][4] ), .C(
        \registers[342][4] ), .D(\registers[343][4] ), .S0(n4203), .S1(n4438), 
        .Y(n2889) );
  MX4X1 U4608 ( .A(\registers[324][4] ), .B(\registers[325][4] ), .C(
        \registers[326][4] ), .D(\registers[327][4] ), .S0(n4204), .S1(n4438), 
        .Y(n2894) );
  MX4X1 U4609 ( .A(\registers[372][4] ), .B(\registers[373][4] ), .C(
        \registers[374][4] ), .D(\registers[375][4] ), .S0(n4203), .S1(n4437), 
        .Y(n2879) );
  MX4X1 U4610 ( .A(\registers[356][4] ), .B(\registers[357][4] ), .C(
        \registers[358][4] ), .D(\registers[359][4] ), .S0(n4203), .S1(n4438), 
        .Y(n2884) );
  MX4X1 U4611 ( .A(\registers[276][4] ), .B(\registers[277][4] ), .C(
        \registers[278][4] ), .D(\registers[279][4] ), .S0(n4205), .S1(n4439), 
        .Y(n2910) );
  MX4X1 U4612 ( .A(\registers[260][4] ), .B(\registers[261][4] ), .C(
        \registers[262][4] ), .D(\registers[263][4] ), .S0(n4205), .S1(n4439), 
        .Y(n2915) );
  MX4X1 U4613 ( .A(\registers[308][4] ), .B(\registers[309][4] ), .C(
        \registers[310][4] ), .D(\registers[311][4] ), .S0(n4204), .S1(n4438), 
        .Y(n2900) );
  MX4X1 U4614 ( .A(\registers[292][4] ), .B(\registers[293][4] ), .C(
        \registers[294][4] ), .D(\registers[295][4] ), .S0(n4204), .S1(n4439), 
        .Y(n2905) );
  MX4X1 U4615 ( .A(\registers[468][4] ), .B(\registers[469][4] ), .C(
        \registers[470][4] ), .D(\registers[471][4] ), .S0(n4201), .S1(n4435), 
        .Y(n2847) );
  MX4X1 U4616 ( .A(\registers[452][4] ), .B(\registers[453][4] ), .C(
        \registers[454][4] ), .D(\registers[455][4] ), .S0(n4201), .S1(n4436), 
        .Y(n2852) );
  MX4X1 U4617 ( .A(\registers[500][4] ), .B(\registers[501][4] ), .C(
        \registers[502][4] ), .D(\registers[503][4] ), .S0(n4200), .S1(n4435), 
        .Y(n2837) );
  MX4X1 U4618 ( .A(\registers[484][4] ), .B(\registers[485][4] ), .C(
        \registers[486][4] ), .D(\registers[487][4] ), .S0(n4200), .S1(n4435), 
        .Y(n2842) );
  MX4X1 U4619 ( .A(\registers[404][4] ), .B(\registers[405][4] ), .C(
        \registers[406][4] ), .D(\registers[407][4] ), .S0(n4202), .S1(n4437), 
        .Y(n2868) );
  MX4X1 U4620 ( .A(\registers[388][4] ), .B(\registers[389][4] ), .C(
        \registers[390][4] ), .D(\registers[391][4] ), .S0(n4202), .S1(n4437), 
        .Y(n2873) );
  MX4X1 U4621 ( .A(\registers[436][4] ), .B(\registers[437][4] ), .C(
        \registers[438][4] ), .D(\registers[439][4] ), .S0(n4201), .S1(n4436), 
        .Y(n2858) );
  MX4X1 U4622 ( .A(\registers[420][4] ), .B(\registers[421][4] ), .C(
        \registers[422][4] ), .D(\registers[423][4] ), .S0(n4202), .S1(n4436), 
        .Y(n2863) );
  MX4X1 U4623 ( .A(\registers[84][4] ), .B(\registers[85][4] ), .C(
        \registers[86][4] ), .D(\registers[87][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2974) );
  MX4X1 U4624 ( .A(\registers[68][4] ), .B(\registers[69][4] ), .C(
        \registers[70][4] ), .D(\registers[71][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2979) );
  MX4X1 U4625 ( .A(\registers[116][4] ), .B(\registers[117][4] ), .C(
        \registers[118][4] ), .D(\registers[119][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2964) );
  MX4X1 U4626 ( .A(\registers[100][4] ), .B(\registers[101][4] ), .C(
        \registers[102][4] ), .D(\registers[103][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2969) );
  MX4X1 U4627 ( .A(\registers[20][4] ), .B(\registers[21][4] ), .C(
        \registers[22][4] ), .D(\registers[23][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2995) );
  MX4X1 U4628 ( .A(\registers[4][4] ), .B(\registers[5][4] ), .C(
        \registers[6][4] ), .D(\registers[7][4] ), .S0(n4210), .S1(n4444), .Y(
        n3000) );
  MX4X1 U4629 ( .A(\registers[52][4] ), .B(\registers[53][4] ), .C(
        \registers[54][4] ), .D(\registers[55][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2985) );
  MX4X1 U4630 ( .A(\registers[36][4] ), .B(\registers[37][4] ), .C(
        \registers[38][4] ), .D(\registers[39][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2990) );
  MX4X1 U4631 ( .A(\registers[212][4] ), .B(\registers[213][4] ), .C(
        \registers[214][4] ), .D(\registers[215][4] ), .S0(n4206), .S1(n4440), 
        .Y(n2932) );
  MX4X1 U4632 ( .A(\registers[196][4] ), .B(\registers[197][4] ), .C(
        \registers[198][4] ), .D(\registers[199][4] ), .S0(n4206), .S1(n4441), 
        .Y(n2937) );
  MX4X1 U4633 ( .A(\registers[244][4] ), .B(\registers[245][4] ), .C(
        \registers[246][4] ), .D(\registers[247][4] ), .S0(n4205), .S1(n4440), 
        .Y(n2922) );
  MX4X1 U4634 ( .A(\registers[228][4] ), .B(\registers[229][4] ), .C(
        \registers[230][4] ), .D(\registers[231][4] ), .S0(n4206), .S1(n4440), 
        .Y(n2927) );
  MX4X1 U4635 ( .A(\registers[148][4] ), .B(\registers[149][4] ), .C(
        \registers[150][4] ), .D(\registers[151][4] ), .S0(n4207), .S1(n4442), 
        .Y(n2953) );
  MX4X1 U4636 ( .A(\registers[132][4] ), .B(\registers[133][4] ), .C(
        \registers[134][4] ), .D(\registers[135][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2958) );
  MX4X1 U4637 ( .A(\registers[180][4] ), .B(\registers[181][4] ), .C(
        \registers[182][4] ), .D(\registers[183][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2943) );
  MX4X1 U4638 ( .A(\registers[164][4] ), .B(\registers[165][4] ), .C(
        \registers[166][4] ), .D(\registers[167][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2948) );
  MX4X1 U4639 ( .A(\registers[852][4] ), .B(\registers[853][4] ), .C(
        \registers[854][4] ), .D(\registers[855][4] ), .S0(n4193), .S1(n4428), 
        .Y(n2719) );
  MX4X1 U4640 ( .A(\registers[836][4] ), .B(\registers[837][4] ), .C(
        \registers[838][4] ), .D(\registers[839][4] ), .S0(n4193), .S1(n4428), 
        .Y(n2724) );
  MX4X1 U4641 ( .A(\registers[884][4] ), .B(\registers[885][4] ), .C(
        \registers[886][4] ), .D(\registers[887][4] ), .S0(n4192), .S1(n4427), 
        .Y(n2709) );
  MX4X1 U4642 ( .A(\registers[868][4] ), .B(\registers[869][4] ), .C(
        \registers[870][4] ), .D(\registers[871][4] ), .S0(n4192), .S1(n4428), 
        .Y(n2714) );
  MX4X1 U4643 ( .A(\registers[788][4] ), .B(\registers[789][4] ), .C(
        \registers[790][4] ), .D(\registers[791][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2740) );
  MX4X1 U4644 ( .A(\registers[772][4] ), .B(\registers[773][4] ), .C(
        \registers[774][4] ), .D(\registers[775][4] ), .S0(n4194), .S1(n4430), 
        .Y(n2745) );
  MX4X1 U4645 ( .A(\registers[820][4] ), .B(\registers[821][4] ), .C(
        \registers[822][4] ), .D(\registers[823][4] ), .S0(n4193), .S1(n4429), 
        .Y(n2730) );
  MX4X1 U4646 ( .A(\registers[804][4] ), .B(\registers[805][4] ), .C(
        \registers[806][4] ), .D(\registers[807][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2735) );
  MX4X1 U4647 ( .A(\registers[980][4] ), .B(\registers[981][4] ), .C(
        \registers[982][4] ), .D(\registers[983][4] ), .S0(n4190), .S1(n4426), 
        .Y(n2677) );
  MX4X1 U4648 ( .A(\registers[964][4] ), .B(\registers[965][4] ), .C(
        \registers[966][4] ), .D(\registers[967][4] ), .S0(n4190), .S1(n4426), 
        .Y(n2682) );
  MX4X1 U4649 ( .A(\registers[1012][4] ), .B(\registers[1013][4] ), .C(
        \registers[1014][4] ), .D(\registers[1015][4] ), .S0(n4189), .S1(n4425), .Y(n2667) );
  MX4X1 U4650 ( .A(\registers[996][4] ), .B(\registers[997][4] ), .C(
        \registers[998][4] ), .D(\registers[999][4] ), .S0(n4190), .S1(n4425), 
        .Y(n2672) );
  MX4X1 U4651 ( .A(\registers[916][4] ), .B(\registers[917][4] ), .C(
        \registers[918][4] ), .D(\registers[919][4] ), .S0(n4191), .S1(n4427), 
        .Y(n2698) );
  MX4X1 U4652 ( .A(\registers[900][4] ), .B(\registers[901][4] ), .C(
        \registers[902][4] ), .D(\registers[903][4] ), .S0(n4192), .S1(n4427), 
        .Y(n2703) );
  MX4X1 U4653 ( .A(\registers[948][4] ), .B(\registers[949][4] ), .C(
        \registers[950][4] ), .D(\registers[951][4] ), .S0(n4191), .S1(n4426), 
        .Y(n2688) );
  MX4X1 U4654 ( .A(\registers[932][4] ), .B(\registers[933][4] ), .C(
        \registers[934][4] ), .D(\registers[935][4] ), .S0(n4191), .S1(n4426), 
        .Y(n2693) );
  MX4X1 U4655 ( .A(\registers[596][4] ), .B(\registers[597][4] ), .C(
        \registers[598][4] ), .D(\registers[599][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2804) );
  MX4X1 U4656 ( .A(\registers[580][4] ), .B(\registers[581][4] ), .C(
        \registers[582][4] ), .D(\registers[583][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2809) );
  MX4X1 U4657 ( .A(\registers[628][4] ), .B(\registers[629][4] ), .C(
        \registers[630][4] ), .D(\registers[631][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2794) );
  MX4X1 U4658 ( .A(\registers[612][4] ), .B(\registers[613][4] ), .C(
        \registers[614][4] ), .D(\registers[615][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2799) );
  MX4X1 U4659 ( .A(\registers[532][4] ), .B(\registers[533][4] ), .C(
        \registers[534][4] ), .D(\registers[535][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2825) );
  MX4X1 U4660 ( .A(\registers[516][4] ), .B(\registers[517][4] ), .C(
        \registers[518][4] ), .D(\registers[519][4] ), .S0(n4200), .S1(n4434), 
        .Y(n2830) );
  MX4X1 U4661 ( .A(\registers[564][4] ), .B(\registers[565][4] ), .C(
        \registers[566][4] ), .D(\registers[567][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2815) );
  MX4X1 U4662 ( .A(\registers[548][4] ), .B(\registers[549][4] ), .C(
        \registers[550][4] ), .D(\registers[551][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2820) );
  MX4X1 U4663 ( .A(\registers[724][4] ), .B(\registers[725][4] ), .C(
        \registers[726][4] ), .D(\registers[727][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2762) );
  MX4X1 U4664 ( .A(\registers[708][4] ), .B(\registers[709][4] ), .C(
        \registers[710][4] ), .D(\registers[711][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2767) );
  MX4X1 U4665 ( .A(\registers[756][4] ), .B(\registers[757][4] ), .C(
        \registers[758][4] ), .D(\registers[759][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2752) );
  MX4X1 U4666 ( .A(\registers[740][4] ), .B(\registers[741][4] ), .C(
        \registers[742][4] ), .D(\registers[743][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2757) );
  MX4X1 U4667 ( .A(\registers[660][4] ), .B(\registers[661][4] ), .C(
        \registers[662][4] ), .D(\registers[663][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2783) );
  MX4X1 U4668 ( .A(\registers[644][4] ), .B(\registers[645][4] ), .C(
        \registers[646][4] ), .D(\registers[647][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2788) );
  MX4X1 U4669 ( .A(\registers[692][4] ), .B(\registers[693][4] ), .C(
        \registers[694][4] ), .D(\registers[695][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2773) );
  MX4X1 U4670 ( .A(\registers[676][4] ), .B(\registers[677][4] ), .C(
        \registers[678][4] ), .D(\registers[679][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2778) );
  MX4X1 U4671 ( .A(\registers[340][5] ), .B(\registers[341][5] ), .C(
        \registers[342][5] ), .D(\registers[343][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3229) );
  MX4X1 U4672 ( .A(\registers[324][5] ), .B(\registers[325][5] ), .C(
        \registers[326][5] ), .D(\registers[327][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3234) );
  MX4X1 U4673 ( .A(\registers[372][5] ), .B(\registers[373][5] ), .C(
        \registers[374][5] ), .D(\registers[375][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3219) );
  MX4X1 U4674 ( .A(\registers[356][5] ), .B(\registers[357][5] ), .C(
        \registers[358][5] ), .D(\registers[359][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3224) );
  MX4X1 U4675 ( .A(\registers[276][5] ), .B(\registers[277][5] ), .C(
        \registers[278][5] ), .D(\registers[279][5] ), .S0(n4226), .S1(n4459), 
        .Y(n3250) );
  MX4X1 U4676 ( .A(\registers[260][5] ), .B(\registers[261][5] ), .C(
        \registers[262][5] ), .D(\registers[263][5] ), .S0(n4226), .S1(n4459), 
        .Y(n3255) );
  MX4X1 U4677 ( .A(\registers[308][5] ), .B(\registers[309][5] ), .C(
        \registers[310][5] ), .D(\registers[311][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3240) );
  MX4X1 U4678 ( .A(\registers[292][5] ), .B(\registers[293][5] ), .C(
        \registers[294][5] ), .D(\registers[295][5] ), .S0(n4226), .S1(n4458), 
        .Y(n3245) );
  MX4X1 U4679 ( .A(\registers[468][5] ), .B(\registers[469][5] ), .C(
        \registers[470][5] ), .D(\registers[471][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3187) );
  MX4X1 U4680 ( .A(\registers[452][5] ), .B(\registers[453][5] ), .C(
        \registers[454][5] ), .D(\registers[455][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3192) );
  MX4X1 U4681 ( .A(\registers[500][5] ), .B(\registers[501][5] ), .C(
        \registers[502][5] ), .D(\registers[503][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3177) );
  MX4X1 U4682 ( .A(\registers[484][5] ), .B(\registers[485][5] ), .C(
        \registers[486][5] ), .D(\registers[487][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3182) );
  MX4X1 U4683 ( .A(\registers[404][5] ), .B(\registers[405][5] ), .C(
        \registers[406][5] ), .D(\registers[407][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3208) );
  MX4X1 U4684 ( .A(\registers[388][5] ), .B(\registers[389][5] ), .C(
        \registers[390][5] ), .D(\registers[391][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3213) );
  MX4X1 U4685 ( .A(\registers[436][5] ), .B(\registers[437][5] ), .C(
        \registers[438][5] ), .D(\registers[439][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3198) );
  MX4X1 U4686 ( .A(\registers[420][5] ), .B(\registers[421][5] ), .C(
        \registers[422][5] ), .D(\registers[423][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3203) );
  MX4X1 U4687 ( .A(\registers[84][5] ), .B(\registers[85][5] ), .C(
        \registers[86][5] ), .D(\registers[87][5] ), .S0(n4230), .S1(n4462), 
        .Y(n3314) );
  MX4X1 U4688 ( .A(\registers[68][5] ), .B(\registers[69][5] ), .C(
        \registers[70][5] ), .D(\registers[71][5] ), .S0(n4230), .S1(n4463), 
        .Y(n3319) );
  MX4X1 U4689 ( .A(\registers[116][5] ), .B(\registers[117][5] ), .C(
        \registers[118][5] ), .D(\registers[119][5] ), .S0(n4229), .S1(n4462), 
        .Y(n3304) );
  MX4X1 U4690 ( .A(\registers[100][5] ), .B(\registers[101][5] ), .C(
        \registers[102][5] ), .D(\registers[103][5] ), .S0(n4230), .S1(n4462), 
        .Y(n3309) );
  MX4X1 U4691 ( .A(\registers[20][5] ), .B(\registers[21][5] ), .C(
        \registers[22][5] ), .D(\registers[23][5] ), .S0(n4231), .S1(n4464), 
        .Y(n3335) );
  MX4X1 U4692 ( .A(\registers[4][5] ), .B(\registers[5][5] ), .C(
        \registers[6][5] ), .D(\registers[7][5] ), .S0(n4232), .S1(n4464), .Y(
        n3340) );
  MX4X1 U4693 ( .A(\registers[52][5] ), .B(\registers[53][5] ), .C(
        \registers[54][5] ), .D(\registers[55][5] ), .S0(n4231), .S1(n4463), 
        .Y(n3325) );
  MX4X1 U4694 ( .A(\registers[36][5] ), .B(\registers[37][5] ), .C(
        \registers[38][5] ), .D(\registers[39][5] ), .S0(n4231), .S1(n4463), 
        .Y(n3330) );
  MX4X1 U4695 ( .A(\registers[212][5] ), .B(\registers[213][5] ), .C(
        \registers[214][5] ), .D(\registers[215][5] ), .S0(n4227), .S1(n4460), 
        .Y(n3272) );
  MX4X1 U4696 ( .A(\registers[196][5] ), .B(\registers[197][5] ), .C(
        \registers[198][5] ), .D(\registers[199][5] ), .S0(n4228), .S1(n4460), 
        .Y(n3277) );
  MX4X1 U4697 ( .A(\registers[244][5] ), .B(\registers[245][5] ), .C(
        \registers[246][5] ), .D(\registers[247][5] ), .S0(n4227), .S1(n4459), 
        .Y(n3262) );
  MX4X1 U4698 ( .A(\registers[228][5] ), .B(\registers[229][5] ), .C(
        \registers[230][5] ), .D(\registers[231][5] ), .S0(n4227), .S1(n4460), 
        .Y(n3267) );
  MX4X1 U4699 ( .A(\registers[148][5] ), .B(\registers[149][5] ), .C(
        \registers[150][5] ), .D(\registers[151][5] ), .S0(n4229), .S1(n4461), 
        .Y(n3293) );
  MX4X1 U4700 ( .A(\registers[132][5] ), .B(\registers[133][5] ), .C(
        \registers[134][5] ), .D(\registers[135][5] ), .S0(n4229), .S1(n4462), 
        .Y(n3298) );
  MX4X1 U4701 ( .A(\registers[180][5] ), .B(\registers[181][5] ), .C(
        \registers[182][5] ), .D(\registers[183][5] ), .S0(n4228), .S1(n4461), 
        .Y(n3283) );
  MX4X1 U4702 ( .A(\registers[164][5] ), .B(\registers[165][5] ), .C(
        \registers[166][5] ), .D(\registers[167][5] ), .S0(n4228), .S1(n4461), 
        .Y(n3288) );
  MX4X1 U4703 ( .A(\registers[852][5] ), .B(\registers[853][5] ), .C(
        \registers[854][5] ), .D(\registers[855][5] ), .S0(n4214), .S1(n4448), 
        .Y(n3059) );
  MX4X1 U4704 ( .A(\registers[836][5] ), .B(\registers[837][5] ), .C(
        \registers[838][5] ), .D(\registers[839][5] ), .S0(n4214), .S1(n4448), 
        .Y(n3064) );
  MX4X1 U4705 ( .A(\registers[884][5] ), .B(\registers[885][5] ), .C(
        \registers[886][5] ), .D(\registers[887][5] ), .S0(n4213), .S1(n4447), 
        .Y(n3049) );
  MX4X1 U4706 ( .A(\registers[868][5] ), .B(\registers[869][5] ), .C(
        \registers[870][5] ), .D(\registers[871][5] ), .S0(n4214), .S1(n4447), 
        .Y(n3054) );
  MX4X1 U4707 ( .A(\registers[788][5] ), .B(\registers[789][5] ), .C(
        \registers[790][5] ), .D(\registers[791][5] ), .S0(n4215), .S1(n4449), 
        .Y(n3080) );
  MX4X1 U4708 ( .A(\registers[772][5] ), .B(\registers[773][5] ), .C(
        \registers[774][5] ), .D(\registers[775][5] ), .S0(n4216), .S1(n4449), 
        .Y(n3085) );
  MX4X1 U4709 ( .A(\registers[820][5] ), .B(\registers[821][5] ), .C(
        \registers[822][5] ), .D(\registers[823][5] ), .S0(n4215), .S1(n4448), 
        .Y(n3070) );
  MX4X1 U4710 ( .A(\registers[804][5] ), .B(\registers[805][5] ), .C(
        \registers[806][5] ), .D(\registers[807][5] ), .S0(n4215), .S1(n4449), 
        .Y(n3075) );
  MX4X1 U4711 ( .A(\registers[980][5] ), .B(\registers[981][5] ), .C(
        \registers[982][5] ), .D(\registers[983][5] ), .S0(n4211), .S1(n4445), 
        .Y(n3017) );
  MX4X1 U4712 ( .A(\registers[964][5] ), .B(\registers[965][5] ), .C(
        \registers[966][5] ), .D(\registers[967][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3022) );
  MX4X1 U4713 ( .A(\registers[1012][5] ), .B(\registers[1013][5] ), .C(
        \registers[1014][5] ), .D(\registers[1015][5] ), .S0(n4211), .S1(n4445), .Y(n3007) );
  MX4X1 U4714 ( .A(\registers[996][5] ), .B(\registers[997][5] ), .C(
        \registers[998][5] ), .D(\registers[999][5] ), .S0(n4211), .S1(n4445), 
        .Y(n3012) );
  MX4X1 U4715 ( .A(\registers[916][5] ), .B(\registers[917][5] ), .C(
        \registers[918][5] ), .D(\registers[919][5] ), .S0(n4213), .S1(n4446), 
        .Y(n3038) );
  MX4X1 U4716 ( .A(\registers[900][5] ), .B(\registers[901][5] ), .C(
        \registers[902][5] ), .D(\registers[903][5] ), .S0(n4213), .S1(n4447), 
        .Y(n3043) );
  MX4X1 U4717 ( .A(\registers[948][5] ), .B(\registers[949][5] ), .C(
        \registers[950][5] ), .D(\registers[951][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3028) );
  MX4X1 U4718 ( .A(\registers[932][5] ), .B(\registers[933][5] ), .C(
        \registers[934][5] ), .D(\registers[935][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3033) );
  MX4X1 U4719 ( .A(\registers[596][5] ), .B(\registers[597][5] ), .C(
        \registers[598][5] ), .D(\registers[599][5] ), .S0(n4219), .S1(n4453), 
        .Y(n3144) );
  MX4X1 U4720 ( .A(\registers[580][5] ), .B(\registers[581][5] ), .C(
        \registers[582][5] ), .D(\registers[583][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3149) );
  MX4X1 U4721 ( .A(\registers[628][5] ), .B(\registers[629][5] ), .C(
        \registers[630][5] ), .D(\registers[631][5] ), .S0(n4219), .S1(n4452), 
        .Y(n3134) );
  MX4X1 U4722 ( .A(\registers[612][5] ), .B(\registers[613][5] ), .C(
        \registers[614][5] ), .D(\registers[615][5] ), .S0(n4219), .S1(n4452), 
        .Y(n3139) );
  MX4X1 U4723 ( .A(\registers[532][5] ), .B(\registers[533][5] ), .C(
        \registers[534][5] ), .D(\registers[535][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3165) );
  MX4X1 U4724 ( .A(\registers[516][5] ), .B(\registers[517][5] ), .C(
        \registers[518][5] ), .D(\registers[519][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3170) );
  MX4X1 U4725 ( .A(\registers[564][5] ), .B(\registers[565][5] ), .C(
        \registers[566][5] ), .D(\registers[567][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3155) );
  MX4X1 U4726 ( .A(\registers[548][5] ), .B(\registers[549][5] ), .C(
        \registers[550][5] ), .D(\registers[551][5] ), .S0(n4220), .S1(n4454), 
        .Y(n3160) );
  MX4X1 U4727 ( .A(\registers[724][5] ), .B(\registers[725][5] ), .C(
        \registers[726][5] ), .D(\registers[727][5] ), .S0(n4217), .S1(n4450), 
        .Y(n3102) );
  MX4X1 U4728 ( .A(\registers[708][5] ), .B(\registers[709][5] ), .C(
        \registers[710][5] ), .D(\registers[711][5] ), .S0(n4217), .S1(n4450), 
        .Y(n3107) );
  MX4X1 U4729 ( .A(\registers[756][5] ), .B(\registers[757][5] ), .C(
        \registers[758][5] ), .D(\registers[759][5] ), .S0(n4216), .S1(n4450), 
        .Y(n3092) );
  MX4X1 U4730 ( .A(\registers[740][5] ), .B(\registers[741][5] ), .C(
        \registers[742][5] ), .D(\registers[743][5] ), .S0(n4216), .S1(n4450), 
        .Y(n3097) );
  MX4X1 U4731 ( .A(\registers[660][5] ), .B(\registers[661][5] ), .C(
        \registers[662][5] ), .D(\registers[663][5] ), .S0(n4218), .S1(n4451), 
        .Y(n3123) );
  MX4X1 U4732 ( .A(\registers[644][5] ), .B(\registers[645][5] ), .C(
        \registers[646][5] ), .D(\registers[647][5] ), .S0(n4218), .S1(n4452), 
        .Y(n3128) );
  MX4X1 U4733 ( .A(\registers[692][5] ), .B(\registers[693][5] ), .C(
        \registers[694][5] ), .D(\registers[695][5] ), .S0(n4217), .S1(n4451), 
        .Y(n3113) );
  MX4X1 U4734 ( .A(\registers[676][5] ), .B(\registers[677][5] ), .C(
        \registers[678][5] ), .D(\registers[679][5] ), .S0(n4218), .S1(n4451), 
        .Y(n3118) );
  MX4X1 U4735 ( .A(\registers[340][6] ), .B(\registers[341][6] ), .C(
        \registers[342][6] ), .D(\registers[343][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3569) );
  MX4X1 U4736 ( .A(\registers[324][6] ), .B(\registers[325][6] ), .C(
        \registers[326][6] ), .D(\registers[327][6] ), .S0(n4246), .S1(n4478), 
        .Y(n3574) );
  MX4X1 U4737 ( .A(\registers[372][6] ), .B(\registers[373][6] ), .C(
        \registers[374][6] ), .D(\registers[375][6] ), .S0(n4245), .S1(n4477), 
        .Y(n3559) );
  MX4X1 U4738 ( .A(\registers[356][6] ), .B(\registers[357][6] ), .C(
        \registers[358][6] ), .D(\registers[359][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3564) );
  MX4X1 U4739 ( .A(\registers[276][6] ), .B(\registers[277][6] ), .C(
        \registers[278][6] ), .D(\registers[279][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3590) );
  MX4X1 U4740 ( .A(\registers[260][6] ), .B(\registers[261][6] ), .C(
        \registers[262][6] ), .D(\registers[263][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3595) );
  MX4X1 U4741 ( .A(\registers[308][6] ), .B(\registers[309][6] ), .C(
        \registers[310][6] ), .D(\registers[311][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3580) );
  MX4X1 U4742 ( .A(\registers[292][6] ), .B(\registers[293][6] ), .C(
        \registers[294][6] ), .D(\registers[295][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3585) );
  MX4X1 U4743 ( .A(\registers[468][6] ), .B(\registers[469][6] ), .C(
        \registers[470][6] ), .D(\registers[471][6] ), .S0(n4243), .S1(n4475), 
        .Y(n3527) );
  MX4X1 U4744 ( .A(\registers[452][6] ), .B(\registers[453][6] ), .C(
        \registers[454][6] ), .D(\registers[455][6] ), .S0(n4244), .S1(n4475), 
        .Y(n3532) );
  MX4X1 U4745 ( .A(\registers[500][6] ), .B(\registers[501][6] ), .C(
        \registers[502][6] ), .D(\registers[503][6] ), .S0(n4243), .S1(n4474), 
        .Y(n3517) );
  MX4X1 U4746 ( .A(\registers[484][6] ), .B(\registers[485][6] ), .C(
        \registers[486][6] ), .D(\registers[487][6] ), .S0(n4243), .S1(n4474), 
        .Y(n3522) );
  MX4X1 U4747 ( .A(\registers[404][6] ), .B(\registers[405][6] ), .C(
        \registers[406][6] ), .D(\registers[407][6] ), .S0(n4245), .S1(n4476), 
        .Y(n3548) );
  MX4X1 U4748 ( .A(\registers[388][6] ), .B(\registers[389][6] ), .C(
        \registers[390][6] ), .D(\registers[391][6] ), .S0(n4245), .S1(n4476), 
        .Y(n3553) );
  MX4X1 U4749 ( .A(\registers[436][6] ), .B(\registers[437][6] ), .C(
        \registers[438][6] ), .D(\registers[439][6] ), .S0(n4244), .S1(n4475), 
        .Y(n3538) );
  MX4X1 U4750 ( .A(\registers[420][6] ), .B(\registers[421][6] ), .C(
        \registers[422][6] ), .D(\registers[423][6] ), .S0(n4244), .S1(n4476), 
        .Y(n3543) );
  MX4X1 U4751 ( .A(\registers[84][6] ), .B(\registers[85][6] ), .C(
        \registers[86][6] ), .D(\registers[87][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3654) );
  MX4X1 U4752 ( .A(\registers[68][6] ), .B(\registers[69][6] ), .C(
        \registers[70][6] ), .D(\registers[71][6] ), .S0(n4252), .S1(n4482), 
        .Y(n3659) );
  MX4X1 U4753 ( .A(\registers[116][6] ), .B(\registers[117][6] ), .C(
        \registers[118][6] ), .D(\registers[119][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3644) );
  MX4X1 U4754 ( .A(\registers[100][6] ), .B(\registers[101][6] ), .C(
        \registers[102][6] ), .D(\registers[103][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3649) );
  MX4X1 U4755 ( .A(\registers[20][6] ), .B(\registers[21][6] ), .C(
        \registers[22][6] ), .D(\registers[23][6] ), .S0(n4253), .S1(n4483), 
        .Y(n3675) );
  MX4X1 U4756 ( .A(\registers[4][6] ), .B(\registers[5][6] ), .C(
        \registers[6][6] ), .D(\registers[7][6] ), .S0(n4253), .S1(n4484), .Y(
        n3680) );
  MX4X1 U4757 ( .A(\registers[52][6] ), .B(\registers[53][6] ), .C(
        \registers[54][6] ), .D(\registers[55][6] ), .S0(n4252), .S1(n4483), 
        .Y(n3665) );
  MX4X1 U4758 ( .A(\registers[36][6] ), .B(\registers[37][6] ), .C(
        \registers[38][6] ), .D(\registers[39][6] ), .S0(n4252), .S1(n4483), 
        .Y(n3670) );
  MX4X1 U4759 ( .A(\registers[212][6] ), .B(\registers[213][6] ), .C(
        \registers[214][6] ), .D(\registers[215][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3612) );
  MX4X1 U4760 ( .A(\registers[196][6] ), .B(\registers[197][6] ), .C(
        \registers[198][6] ), .D(\registers[199][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3617) );
  MX4X1 U4761 ( .A(\registers[244][6] ), .B(\registers[245][6] ), .C(
        \registers[246][6] ), .D(\registers[247][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3602) );
  MX4X1 U4762 ( .A(\registers[228][6] ), .B(\registers[229][6] ), .C(
        \registers[230][6] ), .D(\registers[231][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3607) );
  MX4X1 U4763 ( .A(\registers[148][6] ), .B(\registers[149][6] ), .C(
        \registers[150][6] ), .D(\registers[151][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3633) );
  MX4X1 U4764 ( .A(\registers[132][6] ), .B(\registers[133][6] ), .C(
        \registers[134][6] ), .D(\registers[135][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3638) );
  MX4X1 U4765 ( .A(\registers[180][6] ), .B(\registers[181][6] ), .C(
        \registers[182][6] ), .D(\registers[183][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3623) );
  MX4X1 U4766 ( .A(\registers[164][6] ), .B(\registers[165][6] ), .C(
        \registers[166][6] ), .D(\registers[167][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3628) );
  MX4X1 U4767 ( .A(\registers[852][6] ), .B(\registers[853][6] ), .C(
        \registers[854][6] ), .D(\registers[855][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3399) );
  MX4X1 U4768 ( .A(\registers[836][6] ), .B(\registers[837][6] ), .C(
        \registers[838][6] ), .D(\registers[839][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3404) );
  MX4X1 U4769 ( .A(\registers[884][6] ), .B(\registers[885][6] ), .C(
        \registers[886][6] ), .D(\registers[887][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3389) );
  MX4X1 U4770 ( .A(\registers[868][6] ), .B(\registers[869][6] ), .C(
        \registers[870][6] ), .D(\registers[871][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3394) );
  MX4X1 U4771 ( .A(\registers[788][6] ), .B(\registers[789][6] ), .C(
        \registers[790][6] ), .D(\registers[791][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3420) );
  MX4X1 U4772 ( .A(\registers[772][6] ), .B(\registers[773][6] ), .C(
        \registers[774][6] ), .D(\registers[775][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3425) );
  MX4X1 U4773 ( .A(\registers[820][6] ), .B(\registers[821][6] ), .C(
        \registers[822][6] ), .D(\registers[823][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3410) );
  MX4X1 U4774 ( .A(\registers[804][6] ), .B(\registers[805][6] ), .C(
        \registers[806][6] ), .D(\registers[807][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3415) );
  MX4X1 U4775 ( .A(\registers[980][6] ), .B(\registers[981][6] ), .C(
        \registers[982][6] ), .D(\registers[983][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3357) );
  MX4X1 U4776 ( .A(\registers[964][6] ), .B(\registers[965][6] ), .C(
        \registers[966][6] ), .D(\registers[967][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3362) );
  MX4X1 U4777 ( .A(\registers[1012][6] ), .B(\registers[1013][6] ), .C(
        \registers[1014][6] ), .D(\registers[1015][6] ), .S0(n4232), .S1(n4464), .Y(n3347) );
  MX4X1 U4778 ( .A(\registers[996][6] ), .B(\registers[997][6] ), .C(
        \registers[998][6] ), .D(\registers[999][6] ), .S0(n4232), .S1(n4465), 
        .Y(n3352) );
  MX4X1 U4779 ( .A(\registers[916][6] ), .B(\registers[917][6] ), .C(
        \registers[918][6] ), .D(\registers[919][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3378) );
  MX4X1 U4780 ( .A(\registers[900][6] ), .B(\registers[901][6] ), .C(
        \registers[902][6] ), .D(\registers[903][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3383) );
  MX4X1 U4781 ( .A(\registers[948][6] ), .B(\registers[949][6] ), .C(
        \registers[950][6] ), .D(\registers[951][6] ), .S0(n4233), .S1(n4466), 
        .Y(n3368) );
  MX4X1 U4782 ( .A(\registers[932][6] ), .B(\registers[933][6] ), .C(
        \registers[934][6] ), .D(\registers[935][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3373) );
  MX4X1 U4783 ( .A(\registers[596][6] ), .B(\registers[597][6] ), .C(
        \registers[598][6] ), .D(\registers[599][6] ), .S0(n4241), .S1(n4472), 
        .Y(n3484) );
  MX4X1 U4784 ( .A(\registers[580][6] ), .B(\registers[581][6] ), .C(
        \registers[582][6] ), .D(\registers[583][6] ), .S0(n4241), .S1(n4473), 
        .Y(n3489) );
  MX4X1 U4785 ( .A(\registers[628][6] ), .B(\registers[629][6] ), .C(
        \registers[630][6] ), .D(\registers[631][6] ), .S0(n4240), .S1(n4472), 
        .Y(n3474) );
  MX4X1 U4786 ( .A(\registers[612][6] ), .B(\registers[613][6] ), .C(
        \registers[614][6] ), .D(\registers[615][6] ), .S0(n4240), .S1(n4472), 
        .Y(n3479) );
  MX4X1 U4787 ( .A(\registers[532][6] ), .B(\registers[533][6] ), .C(
        \registers[534][6] ), .D(\registers[535][6] ), .S0(n4242), .S1(n4474), 
        .Y(n3505) );
  MX4X1 U4788 ( .A(\registers[516][6] ), .B(\registers[517][6] ), .C(
        \registers[518][6] ), .D(\registers[519][6] ), .S0(n4242), .S1(n4474), 
        .Y(n3510) );
  MX4X1 U4789 ( .A(\registers[564][6] ), .B(\registers[565][6] ), .C(
        \registers[566][6] ), .D(\registers[567][6] ), .S0(n4241), .S1(n4473), 
        .Y(n3495) );
  MX4X1 U4790 ( .A(\registers[548][6] ), .B(\registers[549][6] ), .C(
        \registers[550][6] ), .D(\registers[551][6] ), .S0(n4242), .S1(n4473), 
        .Y(n3500) );
  MX4X1 U4791 ( .A(\registers[724][6] ), .B(\registers[725][6] ), .C(
        \registers[726][6] ), .D(\registers[727][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3442) );
  MX4X1 U4792 ( .A(\registers[708][6] ), .B(\registers[709][6] ), .C(
        \registers[710][6] ), .D(\registers[711][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3447) );
  MX4X1 U4793 ( .A(\registers[756][6] ), .B(\registers[757][6] ), .C(
        \registers[758][6] ), .D(\registers[759][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3432) );
  MX4X1 U4794 ( .A(\registers[740][6] ), .B(\registers[741][6] ), .C(
        \registers[742][6] ), .D(\registers[743][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3437) );
  MX4X1 U4795 ( .A(\registers[660][6] ), .B(\registers[661][6] ), .C(
        \registers[662][6] ), .D(\registers[663][6] ), .S0(n4239), .S1(n4471), 
        .Y(n3463) );
  MX4X1 U4796 ( .A(\registers[644][6] ), .B(\registers[645][6] ), .C(
        \registers[646][6] ), .D(\registers[647][6] ), .S0(n4240), .S1(n4471), 
        .Y(n3468) );
  MX4X1 U4797 ( .A(\registers[692][6] ), .B(\registers[693][6] ), .C(
        \registers[694][6] ), .D(\registers[695][6] ), .S0(n4239), .S1(n4470), 
        .Y(n3453) );
  MX4X1 U4798 ( .A(\registers[676][6] ), .B(\registers[677][6] ), .C(
        \registers[678][6] ), .D(\registers[679][6] ), .S0(n4239), .S1(n4471), 
        .Y(n3458) );
  MX4X1 U4799 ( .A(\registers[340][7] ), .B(\registers[341][7] ), .C(
        \registers[342][7] ), .D(\registers[343][7] ), .S0(n4267), .S1(n4459), 
        .Y(n3909) );
  MX4X1 U4800 ( .A(\registers[324][7] ), .B(\registers[325][7] ), .C(
        \registers[326][7] ), .D(\registers[327][7] ), .S0(n4268), .S1(n4469), 
        .Y(n3914) );
  MX4X1 U4801 ( .A(\registers[372][7] ), .B(\registers[373][7] ), .C(
        \registers[374][7] ), .D(\registers[375][7] ), .S0(n4267), .S1(n4496), 
        .Y(n3899) );
  MX4X1 U4802 ( .A(\registers[356][7] ), .B(\registers[357][7] ), .C(
        \registers[358][7] ), .D(\registers[359][7] ), .S0(n4267), .S1(n4481), 
        .Y(n3904) );
  MX4X1 U4803 ( .A(\registers[276][7] ), .B(\registers[277][7] ), .C(
        \registers[278][7] ), .D(\registers[279][7] ), .S0(n4269), .S1(n4497), 
        .Y(n3930) );
  MX4X1 U4804 ( .A(\registers[260][7] ), .B(\registers[261][7] ), .C(
        \registers[262][7] ), .D(\registers[263][7] ), .S0(n4269), .S1(n4497), 
        .Y(n3935) );
  MX4X1 U4805 ( .A(\registers[308][7] ), .B(\registers[309][7] ), .C(
        \registers[310][7] ), .D(\registers[311][7] ), .S0(n4268), .S1(n4497), 
        .Y(n3920) );
  MX4X1 U4806 ( .A(\registers[292][7] ), .B(\registers[293][7] ), .C(
        \registers[294][7] ), .D(\registers[295][7] ), .S0(n4268), .S1(n4497), 
        .Y(n3925) );
  MX4X1 U4807 ( .A(\registers[468][7] ), .B(\registers[469][7] ), .C(
        \registers[470][7] ), .D(\registers[471][7] ), .S0(n4265), .S1(n4494), 
        .Y(n3867) );
  MX4X1 U4808 ( .A(\registers[452][7] ), .B(\registers[453][7] ), .C(
        \registers[454][7] ), .D(\registers[455][7] ), .S0(n4265), .S1(n4495), 
        .Y(n3872) );
  MX4X1 U4809 ( .A(\registers[500][7] ), .B(\registers[501][7] ), .C(
        \registers[502][7] ), .D(\registers[503][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3857) );
  MX4X1 U4810 ( .A(\registers[484][7] ), .B(\registers[485][7] ), .C(
        \registers[486][7] ), .D(\registers[487][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3862) );
  MX4X1 U4811 ( .A(\registers[404][7] ), .B(\registers[405][7] ), .C(
        \registers[406][7] ), .D(\registers[407][7] ), .S0(n4266), .S1(n4496), 
        .Y(n3888) );
  MX4X1 U4812 ( .A(\registers[388][7] ), .B(\registers[389][7] ), .C(
        \registers[390][7] ), .D(\registers[391][7] ), .S0(n4266), .S1(n4496), 
        .Y(n3893) );
  MX4X1 U4813 ( .A(\registers[436][7] ), .B(\registers[437][7] ), .C(
        \registers[438][7] ), .D(\registers[439][7] ), .S0(n4265), .S1(n4495), 
        .Y(n3878) );
  MX4X1 U4814 ( .A(\registers[420][7] ), .B(\registers[421][7] ), .C(
        \registers[422][7] ), .D(\registers[423][7] ), .S0(n4266), .S1(n4495), 
        .Y(n3883) );
  MX4X1 U4815 ( .A(\registers[84][7] ), .B(\registers[85][7] ), .C(
        \registers[86][7] ), .D(\registers[87][7] ), .S0(n4273), .S1(n4468), 
        .Y(n3994) );
  MX4X1 U4816 ( .A(\registers[68][7] ), .B(\registers[69][7] ), .C(
        \registers[70][7] ), .D(\registers[71][7] ), .S0(n4273), .S1(n4452), 
        .Y(n3999) );
  MX4X1 U4817 ( .A(\registers[116][7] ), .B(\registers[117][7] ), .C(
        \registers[118][7] ), .D(\registers[119][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3984) );
  MX4X1 U4818 ( .A(\registers[100][7] ), .B(\registers[101][7] ), .C(
        \registers[102][7] ), .D(\registers[103][7] ), .S0(n4272), .S1(n4461), 
        .Y(n3989) );
  MX4X1 U4819 ( .A(\registers[20][7] ), .B(\registers[21][7] ), .C(
        \registers[22][7] ), .D(\registers[23][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4015) );
  MX4X1 U4820 ( .A(\registers[4][7] ), .B(\registers[5][7] ), .C(
        \registers[6][7] ), .D(\registers[7][7] ), .S0(n4274), .S1(n4501), .Y(
        n4020) );
  MX4X1 U4821 ( .A(\registers[52][7] ), .B(\registers[53][7] ), .C(
        \registers[54][7] ), .D(\registers[55][7] ), .S0(n4273), .S1(n4456), 
        .Y(n4005) );
  MX4X1 U4822 ( .A(\registers[36][7] ), .B(\registers[37][7] ), .C(
        \registers[38][7] ), .D(\registers[39][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4010) );
  MX4X1 U4823 ( .A(\registers[212][7] ), .B(\registers[213][7] ), .C(
        \registers[214][7] ), .D(\registers[215][7] ), .S0(n4270), .S1(n4498), 
        .Y(n3952) );
  MX4X1 U4824 ( .A(\registers[196][7] ), .B(\registers[197][7] ), .C(
        \registers[198][7] ), .D(\registers[199][7] ), .S0(n4270), .S1(n4499), 
        .Y(n3957) );
  MX4X1 U4825 ( .A(\registers[244][7] ), .B(\registers[245][7] ), .C(
        \registers[246][7] ), .D(\registers[247][7] ), .S0(n4269), .S1(n4498), 
        .Y(n3942) );
  MX4X1 U4826 ( .A(\registers[228][7] ), .B(\registers[229][7] ), .C(
        \registers[230][7] ), .D(\registers[231][7] ), .S0(n4270), .S1(n4498), 
        .Y(n3947) );
  MX4X1 U4827 ( .A(\registers[148][7] ), .B(\registers[149][7] ), .C(
        \registers[150][7] ), .D(\registers[151][7] ), .S0(n4271), .S1(n4500), 
        .Y(n3973) );
  MX4X1 U4828 ( .A(\registers[132][7] ), .B(\registers[133][7] ), .C(
        \registers[134][7] ), .D(\registers[135][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3978) );
  MX4X1 U4829 ( .A(\registers[180][7] ), .B(\registers[181][7] ), .C(
        \registers[182][7] ), .D(\registers[183][7] ), .S0(n4271), .S1(n4499), 
        .Y(n3963) );
  MX4X1 U4830 ( .A(\registers[164][7] ), .B(\registers[165][7] ), .C(
        \registers[166][7] ), .D(\registers[167][7] ), .S0(n4271), .S1(n4499), 
        .Y(n3968) );
  MX4X1 U4831 ( .A(\registers[852][7] ), .B(\registers[853][7] ), .C(
        \registers[854][7] ), .D(\registers[855][7] ), .S0(n4257), .S1(n4487), 
        .Y(n3739) );
  MX4X1 U4832 ( .A(\registers[836][7] ), .B(\registers[837][7] ), .C(
        \registers[838][7] ), .D(\registers[839][7] ), .S0(n4257), .S1(n4487), 
        .Y(n3744) );
  MX4X1 U4833 ( .A(\registers[884][7] ), .B(\registers[885][7] ), .C(
        \registers[886][7] ), .D(\registers[887][7] ), .S0(n4256), .S1(n4486), 
        .Y(n3729) );
  MX4X1 U4834 ( .A(\registers[868][7] ), .B(\registers[869][7] ), .C(
        \registers[870][7] ), .D(\registers[871][7] ), .S0(n4256), .S1(n4487), 
        .Y(n3734) );
  MX4X1 U4835 ( .A(\registers[788][7] ), .B(\registers[789][7] ), .C(
        \registers[790][7] ), .D(\registers[791][7] ), .S0(n4258), .S1(n4488), 
        .Y(n3760) );
  MX4X1 U4836 ( .A(\registers[772][7] ), .B(\registers[773][7] ), .C(
        \registers[774][7] ), .D(\registers[775][7] ), .S0(n4258), .S1(n4489), 
        .Y(n3765) );
  MX4X1 U4837 ( .A(\registers[820][7] ), .B(\registers[821][7] ), .C(
        \registers[822][7] ), .D(\registers[823][7] ), .S0(n4257), .S1(n4488), 
        .Y(n3750) );
  MX4X1 U4838 ( .A(\registers[804][7] ), .B(\registers[805][7] ), .C(
        \registers[806][7] ), .D(\registers[807][7] ), .S0(n4258), .S1(n4488), 
        .Y(n3755) );
  MX4X1 U4839 ( .A(\registers[980][7] ), .B(\registers[981][7] ), .C(
        \registers[982][7] ), .D(\registers[983][7] ), .S0(n4254), .S1(n4485), 
        .Y(n3697) );
  MX4X1 U4840 ( .A(\registers[964][7] ), .B(\registers[965][7] ), .C(
        \registers[966][7] ), .D(\registers[967][7] ), .S0(n4254), .S1(n4485), 
        .Y(n3702) );
  MX4X1 U4841 ( .A(\registers[1012][7] ), .B(\registers[1013][7] ), .C(
        \registers[1014][7] ), .D(\registers[1015][7] ), .S0(n4253), .S1(n4484), .Y(n3687) );
  MX4X1 U4842 ( .A(\registers[996][7] ), .B(\registers[997][7] ), .C(
        \registers[998][7] ), .D(\registers[999][7] ), .S0(n4254), .S1(n4484), 
        .Y(n3692) );
  MX4X1 U4843 ( .A(\registers[916][7] ), .B(\registers[917][7] ), .C(
        \registers[918][7] ), .D(\registers[919][7] ), .S0(n4255), .S1(n4486), 
        .Y(n3718) );
  MX4X1 U4844 ( .A(\registers[900][7] ), .B(\registers[901][7] ), .C(
        \registers[902][7] ), .D(\registers[903][7] ), .S0(n4256), .S1(n4486), 
        .Y(n3723) );
  MX4X1 U4845 ( .A(\registers[948][7] ), .B(\registers[949][7] ), .C(
        \registers[950][7] ), .D(\registers[951][7] ), .S0(n4255), .S1(n4485), 
        .Y(n3708) );
  MX4X1 U4846 ( .A(\registers[932][7] ), .B(\registers[933][7] ), .C(
        \registers[934][7] ), .D(\registers[935][7] ), .S0(n4255), .S1(n4486), 
        .Y(n3713) );
  MX4X1 U4847 ( .A(\registers[596][7] ), .B(\registers[597][7] ), .C(
        \registers[598][7] ), .D(\registers[599][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3824) );
  MX4X1 U4848 ( .A(\registers[580][7] ), .B(\registers[581][7] ), .C(
        \registers[582][7] ), .D(\registers[583][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3829) );
  MX4X1 U4849 ( .A(\registers[628][7] ), .B(\registers[629][7] ), .C(
        \registers[630][7] ), .D(\registers[631][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3814) );
  MX4X1 U4850 ( .A(\registers[612][7] ), .B(\registers[613][7] ), .C(
        \registers[614][7] ), .D(\registers[615][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3819) );
  MX4X1 U4851 ( .A(\registers[532][7] ), .B(\registers[533][7] ), .C(
        \registers[534][7] ), .D(\registers[535][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3845) );
  MX4X1 U4852 ( .A(\registers[516][7] ), .B(\registers[517][7] ), .C(
        \registers[518][7] ), .D(\registers[519][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3850) );
  MX4X1 U4853 ( .A(\registers[564][7] ), .B(\registers[565][7] ), .C(
        \registers[566][7] ), .D(\registers[567][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3835) );
  MX4X1 U4854 ( .A(\registers[548][7] ), .B(\registers[549][7] ), .C(
        \registers[550][7] ), .D(\registers[551][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3840) );
  MX4X1 U4855 ( .A(\registers[724][7] ), .B(\registers[725][7] ), .C(
        \registers[726][7] ), .D(\registers[727][7] ), .S0(n4259), .S1(n4490), 
        .Y(n3782) );
  MX4X1 U4856 ( .A(\registers[708][7] ), .B(\registers[709][7] ), .C(
        \registers[710][7] ), .D(\registers[711][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3787) );
  MX4X1 U4857 ( .A(\registers[756][7] ), .B(\registers[757][7] ), .C(
        \registers[758][7] ), .D(\registers[759][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3772) );
  MX4X1 U4858 ( .A(\registers[740][7] ), .B(\registers[741][7] ), .C(
        \registers[742][7] ), .D(\registers[743][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3777) );
  MX4X1 U4859 ( .A(\registers[660][7] ), .B(\registers[661][7] ), .C(
        \registers[662][7] ), .D(\registers[663][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3803) );
  MX4X1 U4860 ( .A(\registers[644][7] ), .B(\registers[645][7] ), .C(
        \registers[646][7] ), .D(\registers[647][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3808) );
  MX4X1 U4861 ( .A(\registers[692][7] ), .B(\registers[693][7] ), .C(
        \registers[694][7] ), .D(\registers[695][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3793) );
  MX4X1 U4862 ( .A(\registers[676][7] ), .B(\registers[677][7] ), .C(
        \registers[678][7] ), .D(\registers[679][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3798) );
  MX4X1 U4863 ( .A(\registers[340][0] ), .B(\registers[341][0] ), .C(
        \registers[342][0] ), .D(\registers[343][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4874) );
  MX4X1 U4864 ( .A(\registers[324][0] ), .B(\registers[325][0] ), .C(
        \registers[326][0] ), .D(\registers[327][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4879) );
  MX4X1 U4865 ( .A(\registers[372][0] ), .B(\registers[373][0] ), .C(
        \registers[374][0] ), .D(\registers[375][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4864) );
  MX4X1 U4866 ( .A(\registers[356][0] ), .B(\registers[357][0] ), .C(
        \registers[358][0] ), .D(\registers[359][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4869) );
  MX4X1 U4867 ( .A(\registers[276][0] ), .B(\registers[277][0] ), .C(
        \registers[278][0] ), .D(\registers[279][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4895) );
  MX4X1 U4868 ( .A(\registers[260][0] ), .B(\registers[261][0] ), .C(
        \registers[262][0] ), .D(\registers[263][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4900) );
  MX4X1 U4869 ( .A(\registers[308][0] ), .B(\registers[309][0] ), .C(
        \registers[310][0] ), .D(\registers[311][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4885) );
  MX4X1 U4870 ( .A(\registers[292][0] ), .B(\registers[293][0] ), .C(
        \registers[294][0] ), .D(\registers[295][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4890) );
  MX4X1 U4871 ( .A(\registers[468][0] ), .B(\registers[469][0] ), .C(
        \registers[470][0] ), .D(\registers[471][0] ), .S0(n7458), .S1(n7701), 
        .Y(n4832) );
  MX4X1 U4872 ( .A(\registers[452][0] ), .B(\registers[453][0] ), .C(
        \registers[454][0] ), .D(\registers[455][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4837) );
  MX4X1 U4873 ( .A(\registers[500][0] ), .B(\registers[501][0] ), .C(
        \registers[502][0] ), .D(\registers[503][0] ), .S0(n7458), .S1(n7700), 
        .Y(n4822) );
  MX4X1 U4874 ( .A(\registers[484][0] ), .B(\registers[485][0] ), .C(
        \registers[486][0] ), .D(\registers[487][0] ), .S0(n7458), .S1(n7700), 
        .Y(n4827) );
  MX4X1 U4875 ( .A(\registers[404][0] ), .B(\registers[405][0] ), .C(
        \registers[406][0] ), .D(\registers[407][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4853) );
  MX4X1 U4876 ( .A(\registers[388][0] ), .B(\registers[389][0] ), .C(
        \registers[390][0] ), .D(\registers[391][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4858) );
  MX4X1 U4877 ( .A(\registers[436][0] ), .B(\registers[437][0] ), .C(
        \registers[438][0] ), .D(\registers[439][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4843) );
  MX4X1 U4878 ( .A(\registers[420][0] ), .B(\registers[421][0] ), .C(
        \registers[422][0] ), .D(\registers[423][0] ), .S0(n7459), .S1(n7702), 
        .Y(n4848) );
  MX4X1 U4879 ( .A(\registers[84][0] ), .B(\registers[85][0] ), .C(
        \registers[86][0] ), .D(\registers[87][0] ), .S0(n7466), .S1(n7708), 
        .Y(n4959) );
  MX4X1 U4880 ( .A(\registers[68][0] ), .B(\registers[69][0] ), .C(
        \registers[70][0] ), .D(\registers[71][0] ), .S0(n7467), .S1(n7708), 
        .Y(n4964) );
  MX4X1 U4881 ( .A(\registers[116][0] ), .B(\registers[117][0] ), .C(
        \registers[118][0] ), .D(\registers[119][0] ), .S0(n7466), .S1(n7707), 
        .Y(n4949) );
  MX4X1 U4882 ( .A(\registers[100][0] ), .B(\registers[101][0] ), .C(
        \registers[102][0] ), .D(\registers[103][0] ), .S0(n7466), .S1(n7708), 
        .Y(n4954) );
  MX4X1 U4883 ( .A(\registers[20][0] ), .B(\registers[21][0] ), .C(
        \registers[22][0] ), .D(\registers[23][0] ), .S0(n7468), .S1(n7709), 
        .Y(n4980) );
  MX4X1 U4884 ( .A(\registers[4][0] ), .B(\registers[5][0] ), .C(
        \registers[6][0] ), .D(\registers[7][0] ), .S0(n7468), .S1(n7710), .Y(
        n4985) );
  MX4X1 U4885 ( .A(\registers[52][0] ), .B(\registers[53][0] ), .C(
        \registers[54][0] ), .D(\registers[55][0] ), .S0(n7467), .S1(n7709), 
        .Y(n4970) );
  MX4X1 U4886 ( .A(\registers[36][0] ), .B(\registers[37][0] ), .C(
        \registers[38][0] ), .D(\registers[39][0] ), .S0(n7467), .S1(n7709), 
        .Y(n4975) );
  MX4X1 U4887 ( .A(\registers[212][0] ), .B(\registers[213][0] ), .C(
        \registers[214][0] ), .D(\registers[215][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4917) );
  MX4X1 U4888 ( .A(\registers[196][0] ), .B(\registers[197][0] ), .C(
        \registers[198][0] ), .D(\registers[199][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4922) );
  MX4X1 U4889 ( .A(\registers[244][0] ), .B(\registers[245][0] ), .C(
        \registers[246][0] ), .D(\registers[247][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4907) );
  MX4X1 U4890 ( .A(\registers[228][0] ), .B(\registers[229][0] ), .C(
        \registers[230][0] ), .D(\registers[231][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4912) );
  MX4X1 U4891 ( .A(\registers[148][0] ), .B(\registers[149][0] ), .C(
        \registers[150][0] ), .D(\registers[151][0] ), .S0(n7465), .S1(n7707), 
        .Y(n4938) );
  MX4X1 U4892 ( .A(\registers[132][0] ), .B(\registers[133][0] ), .C(
        \registers[134][0] ), .D(\registers[135][0] ), .S0(n7465), .S1(n7707), 
        .Y(n4943) );
  MX4X1 U4893 ( .A(\registers[180][0] ), .B(\registers[181][0] ), .C(
        \registers[182][0] ), .D(\registers[183][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4928) );
  MX4X1 U4894 ( .A(\registers[164][0] ), .B(\registers[165][0] ), .C(
        \registers[166][0] ), .D(\registers[167][0] ), .S0(n7465), .S1(n7706), 
        .Y(n4933) );
  MX4X1 U4895 ( .A(\registers[852][0] ), .B(\registers[853][0] ), .C(
        \registers[854][0] ), .D(\registers[855][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4704) );
  MX4X1 U4896 ( .A(\registers[836][0] ), .B(\registers[837][0] ), .C(
        \registers[838][0] ), .D(\registers[839][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4709) );
  MX4X1 U4897 ( .A(\registers[884][0] ), .B(\registers[885][0] ), .C(
        \registers[886][0] ), .D(\registers[887][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4694) );
  MX4X1 U4898 ( .A(\registers[868][0] ), .B(\registers[869][0] ), .C(
        \registers[870][0] ), .D(\registers[871][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4699) );
  MX4X1 U4899 ( .A(\registers[788][0] ), .B(\registers[789][0] ), .C(
        \registers[790][0] ), .D(\registers[791][0] ), .S0(n7452), .S1(n7694), 
        .Y(n4725) );
  MX4X1 U4900 ( .A(\registers[772][0] ), .B(\registers[773][0] ), .C(
        \registers[774][0] ), .D(\registers[775][0] ), .S0(n7452), .S1(n7695), 
        .Y(n4730) );
  MX4X1 U4901 ( .A(\registers[820][0] ), .B(\registers[821][0] ), .C(
        \registers[822][0] ), .D(\registers[823][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4715) );
  MX4X1 U4902 ( .A(\registers[804][0] ), .B(\registers[805][0] ), .C(
        \registers[806][0] ), .D(\registers[807][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4720) );
  MX4X1 U4903 ( .A(\registers[980][0] ), .B(\registers[981][0] ), .C(
        \registers[982][0] ), .D(\registers[983][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4662) );
  MX4X1 U4904 ( .A(\registers[964][0] ), .B(\registers[965][0] ), .C(
        \registers[966][0] ), .D(\registers[967][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4667) );
  MX4X1 U4905 ( .A(\registers[916][0] ), .B(\registers[917][0] ), .C(
        \registers[918][0] ), .D(\registers[919][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4683) );
  MX4X1 U4906 ( .A(\registers[900][0] ), .B(\registers[901][0] ), .C(
        \registers[902][0] ), .D(\registers[903][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4688) );
  MX4X1 U4907 ( .A(\registers[948][0] ), .B(\registers[949][0] ), .C(
        \registers[950][0] ), .D(\registers[951][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4673) );
  MX4X1 U4908 ( .A(\registers[932][0] ), .B(\registers[933][0] ), .C(
        \registers[934][0] ), .D(\registers[935][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4678) );
  MX4X1 U4909 ( .A(\registers[596][0] ), .B(\registers[597][0] ), .C(
        \registers[598][0] ), .D(\registers[599][0] ), .S0(n7456), .S1(n7698), 
        .Y(n4789) );
  MX4X1 U4910 ( .A(\registers[580][0] ), .B(\registers[581][0] ), .C(
        \registers[582][0] ), .D(\registers[583][0] ), .S0(n7456), .S1(n7698), 
        .Y(n4794) );
  MX4X1 U4911 ( .A(\registers[628][0] ), .B(\registers[629][0] ), .C(
        \registers[630][0] ), .D(\registers[631][0] ), .S0(n7455), .S1(n7698), 
        .Y(n4779) );
  MX4X1 U4912 ( .A(\registers[612][0] ), .B(\registers[613][0] ), .C(
        \registers[614][0] ), .D(\registers[615][0] ), .S0(n7455), .S1(n7698), 
        .Y(n4784) );
  MX4X1 U4913 ( .A(\registers[532][0] ), .B(\registers[533][0] ), .C(
        \registers[534][0] ), .D(\registers[535][0] ), .S0(n7457), .S1(n7699), 
        .Y(n4810) );
  MX4X1 U4914 ( .A(\registers[516][0] ), .B(\registers[517][0] ), .C(
        \registers[518][0] ), .D(\registers[519][0] ), .S0(n7457), .S1(n7700), 
        .Y(n4815) );
  MX4X1 U4915 ( .A(\registers[564][0] ), .B(\registers[565][0] ), .C(
        \registers[566][0] ), .D(\registers[567][0] ), .S0(n7456), .S1(n7699), 
        .Y(n4800) );
  MX4X1 U4916 ( .A(\registers[548][0] ), .B(\registers[549][0] ), .C(
        \registers[550][0] ), .D(\registers[551][0] ), .S0(n7457), .S1(n7699), 
        .Y(n4805) );
  MX4X1 U4917 ( .A(\registers[724][0] ), .B(\registers[725][0] ), .C(
        \registers[726][0] ), .D(\registers[727][0] ), .S0(n7453), .S1(n7696), 
        .Y(n4747) );
  MX4X1 U4918 ( .A(\registers[708][0] ), .B(\registers[709][0] ), .C(
        \registers[710][0] ), .D(\registers[711][0] ), .S0(n7453), .S1(n7696), 
        .Y(n4752) );
  MX4X1 U4919 ( .A(\registers[756][0] ), .B(\registers[757][0] ), .C(
        \registers[758][0] ), .D(\registers[759][0] ), .S0(n7452), .S1(n7695), 
        .Y(n4737) );
  MX4X1 U4920 ( .A(\registers[740][0] ), .B(\registers[741][0] ), .C(
        \registers[742][0] ), .D(\registers[743][0] ), .S0(n7453), .S1(n7695), 
        .Y(n4742) );
  MX4X1 U4921 ( .A(\registers[660][0] ), .B(\registers[661][0] ), .C(
        \registers[662][0] ), .D(\registers[663][0] ), .S0(n7454), .S1(n7697), 
        .Y(n4768) );
  MX4X1 U4922 ( .A(\registers[644][0] ), .B(\registers[645][0] ), .C(
        \registers[646][0] ), .D(\registers[647][0] ), .S0(n7455), .S1(n7697), 
        .Y(n4773) );
  MX4X1 U4923 ( .A(\registers[692][0] ), .B(\registers[693][0] ), .C(
        \registers[694][0] ), .D(\registers[695][0] ), .S0(n7454), .S1(n7696), 
        .Y(n4758) );
  MX4X1 U4924 ( .A(\registers[676][0] ), .B(\registers[677][0] ), .C(
        \registers[678][0] ), .D(\registers[679][0] ), .S0(n7454), .S1(n7697), 
        .Y(n4763) );
  MX4X1 U4925 ( .A(\registers[340][1] ), .B(\registers[341][1] ), .C(
        \registers[342][1] ), .D(\registers[343][1] ), .S0(n7482), .S1(n7723), 
        .Y(n5214) );
  MX4X1 U4926 ( .A(\registers[324][1] ), .B(\registers[325][1] ), .C(
        \registers[326][1] ), .D(\registers[327][1] ), .S0(n7483), .S1(n7723), 
        .Y(n5219) );
  MX4X1 U4927 ( .A(\registers[372][1] ), .B(\registers[373][1] ), .C(
        \registers[374][1] ), .D(\registers[375][1] ), .S0(n7482), .S1(n7722), 
        .Y(n5204) );
  MX4X1 U4928 ( .A(\registers[356][1] ), .B(\registers[357][1] ), .C(
        \registers[358][1] ), .D(\registers[359][1] ), .S0(n7482), .S1(n7722), 
        .Y(n5209) );
  MX4X1 U4929 ( .A(\registers[276][1] ), .B(\registers[277][1] ), .C(
        \registers[278][1] ), .D(\registers[279][1] ), .S0(n7484), .S1(n7724), 
        .Y(n5235) );
  MX4X1 U4930 ( .A(\registers[260][1] ), .B(\registers[261][1] ), .C(
        \registers[262][1] ), .D(\registers[263][1] ), .S0(n7484), .S1(n7724), 
        .Y(n5240) );
  MX4X1 U4931 ( .A(\registers[308][1] ), .B(\registers[309][1] ), .C(
        \registers[310][1] ), .D(\registers[311][1] ), .S0(n7483), .S1(n7723), 
        .Y(n5225) );
  MX4X1 U4932 ( .A(\registers[292][1] ), .B(\registers[293][1] ), .C(
        \registers[294][1] ), .D(\registers[295][1] ), .S0(n7483), .S1(n7724), 
        .Y(n5230) );
  MX4X1 U4933 ( .A(\registers[468][1] ), .B(\registers[469][1] ), .C(
        \registers[470][1] ), .D(\registers[471][1] ), .S0(n7480), .S1(n7720), 
        .Y(n5172) );
  MX4X1 U4934 ( .A(\registers[452][1] ), .B(\registers[453][1] ), .C(
        \registers[454][1] ), .D(\registers[455][1] ), .S0(n7480), .S1(n7721), 
        .Y(n5177) );
  MX4X1 U4935 ( .A(\registers[500][1] ), .B(\registers[501][1] ), .C(
        \registers[502][1] ), .D(\registers[503][1] ), .S0(n7479), .S1(n7720), 
        .Y(n5162) );
  MX4X1 U4936 ( .A(\registers[484][1] ), .B(\registers[485][1] ), .C(
        \registers[486][1] ), .D(\registers[487][1] ), .S0(n7479), .S1(n7720), 
        .Y(n5167) );
  MX4X1 U4937 ( .A(\registers[404][1] ), .B(\registers[405][1] ), .C(
        \registers[406][1] ), .D(\registers[407][1] ), .S0(n7481), .S1(n7722), 
        .Y(n5193) );
  MX4X1 U4938 ( .A(\registers[388][1] ), .B(\registers[389][1] ), .C(
        \registers[390][1] ), .D(\registers[391][1] ), .S0(n7481), .S1(n7722), 
        .Y(n5198) );
  MX4X1 U4939 ( .A(\registers[436][1] ), .B(\registers[437][1] ), .C(
        \registers[438][1] ), .D(\registers[439][1] ), .S0(n7480), .S1(n7721), 
        .Y(n5183) );
  MX4X1 U4940 ( .A(\registers[420][1] ), .B(\registers[421][1] ), .C(
        \registers[422][1] ), .D(\registers[423][1] ), .S0(n7481), .S1(n7721), 
        .Y(n5188) );
  MX4X1 U4941 ( .A(\registers[84][1] ), .B(\registers[85][1] ), .C(
        \registers[86][1] ), .D(\registers[87][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5299) );
  MX4X1 U4942 ( .A(\registers[68][1] ), .B(\registers[69][1] ), .C(
        \registers[70][1] ), .D(\registers[71][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5304) );
  MX4X1 U4943 ( .A(\registers[116][1] ), .B(\registers[117][1] ), .C(
        \registers[118][1] ), .D(\registers[119][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5289) );
  MX4X1 U4944 ( .A(\registers[100][1] ), .B(\registers[101][1] ), .C(
        \registers[102][1] ), .D(\registers[103][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5294) );
  MX4X1 U4945 ( .A(\registers[20][1] ), .B(\registers[21][1] ), .C(
        \registers[22][1] ), .D(\registers[23][1] ), .S0(n7489), .S1(n7729), 
        .Y(n5320) );
  MX4X1 U4946 ( .A(\registers[4][1] ), .B(\registers[5][1] ), .C(
        \registers[6][1] ), .D(\registers[7][1] ), .S0(n7489), .S1(n7729), .Y(
        n5325) );
  MX4X1 U4947 ( .A(\registers[52][1] ), .B(\registers[53][1] ), .C(
        \registers[54][1] ), .D(\registers[55][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5310) );
  MX4X1 U4948 ( .A(\registers[36][1] ), .B(\registers[37][1] ), .C(
        \registers[38][1] ), .D(\registers[39][1] ), .S0(n7489), .S1(n7729), 
        .Y(n5315) );
  MX4X1 U4949 ( .A(\registers[212][1] ), .B(\registers[213][1] ), .C(
        \registers[214][1] ), .D(\registers[215][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5257) );
  MX4X1 U4950 ( .A(\registers[196][1] ), .B(\registers[197][1] ), .C(
        \registers[198][1] ), .D(\registers[199][1] ), .S0(n7485), .S1(n7726), 
        .Y(n5262) );
  MX4X1 U4951 ( .A(\registers[244][1] ), .B(\registers[245][1] ), .C(
        \registers[246][1] ), .D(\registers[247][1] ), .S0(n7484), .S1(n7725), 
        .Y(n5247) );
  MX4X1 U4952 ( .A(\registers[228][1] ), .B(\registers[229][1] ), .C(
        \registers[230][1] ), .D(\registers[231][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5252) );
  MX4X1 U4953 ( .A(\registers[148][1] ), .B(\registers[149][1] ), .C(
        \registers[150][1] ), .D(\registers[151][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5278) );
  MX4X1 U4954 ( .A(\registers[132][1] ), .B(\registers[133][1] ), .C(
        \registers[134][1] ), .D(\registers[135][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5283) );
  MX4X1 U4955 ( .A(\registers[180][1] ), .B(\registers[181][1] ), .C(
        \registers[182][1] ), .D(\registers[183][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5268) );
  MX4X1 U4956 ( .A(\registers[164][1] ), .B(\registers[165][1] ), .C(
        \registers[166][1] ), .D(\registers[167][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5273) );
  MX4X1 U4957 ( .A(\registers[852][1] ), .B(\registers[853][1] ), .C(
        \registers[854][1] ), .D(\registers[855][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5044) );
  MX4X1 U4958 ( .A(\registers[836][1] ), .B(\registers[837][1] ), .C(
        \registers[838][1] ), .D(\registers[839][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5049) );
  MX4X1 U4959 ( .A(\registers[884][1] ), .B(\registers[885][1] ), .C(
        \registers[886][1] ), .D(\registers[887][1] ), .S0(n7471), .S1(n7712), 
        .Y(n5034) );
  MX4X1 U4960 ( .A(\registers[868][1] ), .B(\registers[869][1] ), .C(
        \registers[870][1] ), .D(\registers[871][1] ), .S0(n7471), .S1(n7713), 
        .Y(n5039) );
  MX4X1 U4961 ( .A(\registers[788][1] ), .B(\registers[789][1] ), .C(
        \registers[790][1] ), .D(\registers[791][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5065) );
  MX4X1 U4962 ( .A(\registers[772][1] ), .B(\registers[773][1] ), .C(
        \registers[774][1] ), .D(\registers[775][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5070) );
  MX4X1 U4963 ( .A(\registers[820][1] ), .B(\registers[821][1] ), .C(
        \registers[822][1] ), .D(\registers[823][1] ), .S0(n7472), .S1(n7714), 
        .Y(n5055) );
  MX4X1 U4964 ( .A(\registers[804][1] ), .B(\registers[805][1] ), .C(
        \registers[806][1] ), .D(\registers[807][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5060) );
  MX4X1 U4965 ( .A(\registers[980][1] ), .B(\registers[981][1] ), .C(
        \registers[982][1] ), .D(\registers[983][1] ), .S0(n7469), .S1(n7710), 
        .Y(n5002) );
  MX4X1 U4966 ( .A(\registers[964][1] ), .B(\registers[965][1] ), .C(
        \registers[966][1] ), .D(\registers[967][1] ), .S0(n7469), .S1(n7711), 
        .Y(n5007) );
  MX4X1 U4967 ( .A(\registers[1012][1] ), .B(\registers[1013][1] ), .C(
        \registers[1014][1] ), .D(\registers[1015][1] ), .S0(n7468), .S1(n7710), .Y(n4992) );
  MX4X1 U4968 ( .A(\registers[996][1] ), .B(\registers[997][1] ), .C(
        \registers[998][1] ), .D(\registers[999][1] ), .S0(n7469), .S1(n7710), 
        .Y(n4997) );
  MX4X1 U4969 ( .A(\registers[916][1] ), .B(\registers[917][1] ), .C(
        \registers[918][1] ), .D(\registers[919][1] ), .S0(n7470), .S1(n7712), 
        .Y(n5023) );
  MX4X1 U4970 ( .A(\registers[900][1] ), .B(\registers[901][1] ), .C(
        \registers[902][1] ), .D(\registers[903][1] ), .S0(n7471), .S1(n7712), 
        .Y(n5028) );
  MX4X1 U4971 ( .A(\registers[948][1] ), .B(\registers[949][1] ), .C(
        \registers[950][1] ), .D(\registers[951][1] ), .S0(n7470), .S1(n7711), 
        .Y(n5013) );
  MX4X1 U4972 ( .A(\registers[932][1] ), .B(\registers[933][1] ), .C(
        \registers[934][1] ), .D(\registers[935][1] ), .S0(n7470), .S1(n7711), 
        .Y(n5018) );
  MX4X1 U4973 ( .A(\registers[596][1] ), .B(\registers[597][1] ), .C(
        \registers[598][1] ), .D(\registers[599][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5129) );
  MX4X1 U4974 ( .A(\registers[580][1] ), .B(\registers[581][1] ), .C(
        \registers[582][1] ), .D(\registers[583][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5134) );
  MX4X1 U4975 ( .A(\registers[628][1] ), .B(\registers[629][1] ), .C(
        \registers[630][1] ), .D(\registers[631][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5119) );
  MX4X1 U4976 ( .A(\registers[612][1] ), .B(\registers[613][1] ), .C(
        \registers[614][1] ), .D(\registers[615][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5124) );
  MX4X1 U4977 ( .A(\registers[532][1] ), .B(\registers[533][1] ), .C(
        \registers[534][1] ), .D(\registers[535][1] ), .S0(n7478), .S1(n7719), 
        .Y(n5150) );
  MX4X1 U4978 ( .A(\registers[516][1] ), .B(\registers[517][1] ), .C(
        \registers[518][1] ), .D(\registers[519][1] ), .S0(n7479), .S1(n7719), 
        .Y(n5155) );
  MX4X1 U4979 ( .A(\registers[564][1] ), .B(\registers[565][1] ), .C(
        \registers[566][1] ), .D(\registers[567][1] ), .S0(n7478), .S1(n7718), 
        .Y(n5140) );
  MX4X1 U4980 ( .A(\registers[548][1] ), .B(\registers[549][1] ), .C(
        \registers[550][1] ), .D(\registers[551][1] ), .S0(n7478), .S1(n7719), 
        .Y(n5145) );
  MX4X1 U4981 ( .A(\registers[724][1] ), .B(\registers[725][1] ), .C(
        \registers[726][1] ), .D(\registers[727][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5087) );
  MX4X1 U4982 ( .A(\registers[708][1] ), .B(\registers[709][1] ), .C(
        \registers[710][1] ), .D(\registers[711][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5092) );
  MX4X1 U4983 ( .A(\registers[756][1] ), .B(\registers[757][1] ), .C(
        \registers[758][1] ), .D(\registers[759][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5077) );
  MX4X1 U4984 ( .A(\registers[740][1] ), .B(\registers[741][1] ), .C(
        \registers[742][1] ), .D(\registers[743][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5082) );
  MX4X1 U4985 ( .A(\registers[660][1] ), .B(\registers[661][1] ), .C(
        \registers[662][1] ), .D(\registers[663][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5108) );
  MX4X1 U4986 ( .A(\registers[644][1] ), .B(\registers[645][1] ), .C(
        \registers[646][1] ), .D(\registers[647][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5113) );
  MX4X1 U4987 ( .A(\registers[692][1] ), .B(\registers[693][1] ), .C(
        \registers[694][1] ), .D(\registers[695][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5098) );
  MX4X1 U4988 ( .A(\registers[676][1] ), .B(\registers[677][1] ), .C(
        \registers[678][1] ), .D(\registers[679][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5103) );
  MX4X1 U4989 ( .A(\registers[340][2] ), .B(\registers[341][2] ), .C(
        \registers[342][2] ), .D(\registers[343][2] ), .S0(n7504), .S1(n7742), 
        .Y(n5554) );
  MX4X1 U4990 ( .A(\registers[324][2] ), .B(\registers[325][2] ), .C(
        \registers[326][2] ), .D(\registers[327][2] ), .S0(n7504), .S1(n7743), 
        .Y(n5559) );
  MX4X1 U4991 ( .A(\registers[372][2] ), .B(\registers[373][2] ), .C(
        \registers[374][2] ), .D(\registers[375][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5544) );
  MX4X1 U4992 ( .A(\registers[356][2] ), .B(\registers[357][2] ), .C(
        \registers[358][2] ), .D(\registers[359][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5549) );
  MX4X1 U4993 ( .A(\registers[276][2] ), .B(\registers[277][2] ), .C(
        \registers[278][2] ), .D(\registers[279][2] ), .S0(n7505), .S1(n7744), 
        .Y(n5575) );
  MX4X1 U4994 ( .A(\registers[260][2] ), .B(\registers[261][2] ), .C(
        \registers[262][2] ), .D(\registers[263][2] ), .S0(n7505), .S1(n7744), 
        .Y(n5580) );
  MX4X1 U4995 ( .A(\registers[308][2] ), .B(\registers[309][2] ), .C(
        \registers[310][2] ), .D(\registers[311][2] ), .S0(n7504), .S1(n7743), 
        .Y(n5565) );
  MX4X1 U4996 ( .A(\registers[292][2] ), .B(\registers[293][2] ), .C(
        \registers[294][2] ), .D(\registers[295][2] ), .S0(n7505), .S1(n7743), 
        .Y(n5570) );
  MX4X1 U4997 ( .A(\registers[468][2] ), .B(\registers[469][2] ), .C(
        \registers[470][2] ), .D(\registers[471][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5512) );
  MX4X1 U4998 ( .A(\registers[452][2] ), .B(\registers[453][2] ), .C(
        \registers[454][2] ), .D(\registers[455][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5517) );
  MX4X1 U4999 ( .A(\registers[500][2] ), .B(\registers[501][2] ), .C(
        \registers[502][2] ), .D(\registers[503][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5502) );
  MX4X1 U5000 ( .A(\registers[484][2] ), .B(\registers[485][2] ), .C(
        \registers[486][2] ), .D(\registers[487][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5507) );
  MX4X1 U5001 ( .A(\registers[404][2] ), .B(\registers[405][2] ), .C(
        \registers[406][2] ), .D(\registers[407][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5533) );
  MX4X1 U5002 ( .A(\registers[388][2] ), .B(\registers[389][2] ), .C(
        \registers[390][2] ), .D(\registers[391][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5538) );
  MX4X1 U5003 ( .A(\registers[436][2] ), .B(\registers[437][2] ), .C(
        \registers[438][2] ), .D(\registers[439][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5523) );
  MX4X1 U5004 ( .A(\registers[420][2] ), .B(\registers[421][2] ), .C(
        \registers[422][2] ), .D(\registers[423][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5528) );
  MX4X1 U5005 ( .A(\registers[84][2] ), .B(\registers[85][2] ), .C(
        \registers[86][2] ), .D(\registers[87][2] ), .S0(n7509), .S1(n7747), 
        .Y(n5639) );
  MX4X1 U5006 ( .A(\registers[68][2] ), .B(\registers[69][2] ), .C(
        \registers[70][2] ), .D(\registers[71][2] ), .S0(n7509), .S1(n7748), 
        .Y(n5644) );
  MX4X1 U5007 ( .A(\registers[116][2] ), .B(\registers[117][2] ), .C(
        \registers[118][2] ), .D(\registers[119][2] ), .S0(n7508), .S1(n7747), 
        .Y(n5629) );
  MX4X1 U5008 ( .A(\registers[100][2] ), .B(\registers[101][2] ), .C(
        \registers[102][2] ), .D(\registers[103][2] ), .S0(n7509), .S1(n7747), 
        .Y(n5634) );
  MX4X1 U5009 ( .A(\registers[20][2] ), .B(\registers[21][2] ), .C(
        \registers[22][2] ), .D(\registers[23][2] ), .S0(n7510), .S1(n7749), 
        .Y(n5660) );
  MX4X1 U5010 ( .A(\registers[4][2] ), .B(\registers[5][2] ), .C(
        \registers[6][2] ), .D(\registers[7][2] ), .S0(n7511), .S1(n7749), .Y(
        n5665) );
  MX4X1 U5011 ( .A(\registers[52][2] ), .B(\registers[53][2] ), .C(
        \registers[54][2] ), .D(\registers[55][2] ), .S0(n7510), .S1(n7748), 
        .Y(n5650) );
  MX4X1 U5012 ( .A(\registers[36][2] ), .B(\registers[37][2] ), .C(
        \registers[38][2] ), .D(\registers[39][2] ), .S0(n7510), .S1(n7748), 
        .Y(n5655) );
  MX4X1 U5013 ( .A(\registers[212][2] ), .B(\registers[213][2] ), .C(
        \registers[214][2] ), .D(\registers[215][2] ), .S0(n7506), .S1(n7745), 
        .Y(n5597) );
  MX4X1 U5014 ( .A(\registers[196][2] ), .B(\registers[197][2] ), .C(
        \registers[198][2] ), .D(\registers[199][2] ), .S0(n7507), .S1(n7745), 
        .Y(n5602) );
  MX4X1 U5015 ( .A(\registers[244][2] ), .B(\registers[245][2] ), .C(
        \registers[246][2] ), .D(\registers[247][2] ), .S0(n7506), .S1(n7744), 
        .Y(n5587) );
  MX4X1 U5016 ( .A(\registers[228][2] ), .B(\registers[229][2] ), .C(
        \registers[230][2] ), .D(\registers[231][2] ), .S0(n7506), .S1(n7745), 
        .Y(n5592) );
  MX4X1 U5017 ( .A(\registers[148][2] ), .B(\registers[149][2] ), .C(
        \registers[150][2] ), .D(\registers[151][2] ), .S0(n7508), .S1(n7746), 
        .Y(n5618) );
  MX4X1 U5018 ( .A(\registers[132][2] ), .B(\registers[133][2] ), .C(
        \registers[134][2] ), .D(\registers[135][2] ), .S0(n7508), .S1(n7746), 
        .Y(n5623) );
  MX4X1 U5019 ( .A(\registers[180][2] ), .B(\registers[181][2] ), .C(
        \registers[182][2] ), .D(\registers[183][2] ), .S0(n7507), .S1(n7746), 
        .Y(n5608) );
  MX4X1 U5020 ( .A(\registers[164][2] ), .B(\registers[165][2] ), .C(
        \registers[166][2] ), .D(\registers[167][2] ), .S0(n7507), .S1(n7746), 
        .Y(n5613) );
  MX4X1 U5021 ( .A(\registers[852][2] ), .B(\registers[853][2] ), .C(
        \registers[854][2] ), .D(\registers[855][2] ), .S0(n7493), .S1(n7733), 
        .Y(n5384) );
  MX4X1 U5022 ( .A(\registers[836][2] ), .B(\registers[837][2] ), .C(
        \registers[838][2] ), .D(\registers[839][2] ), .S0(n7493), .S1(n7733), 
        .Y(n5389) );
  MX4X1 U5023 ( .A(\registers[884][2] ), .B(\registers[885][2] ), .C(
        \registers[886][2] ), .D(\registers[887][2] ), .S0(n7492), .S1(n7732), 
        .Y(n5374) );
  MX4X1 U5024 ( .A(\registers[868][2] ), .B(\registers[869][2] ), .C(
        \registers[870][2] ), .D(\registers[871][2] ), .S0(n7493), .S1(n7732), 
        .Y(n5379) );
  MX4X1 U5025 ( .A(\registers[788][2] ), .B(\registers[789][2] ), .C(
        \registers[790][2] ), .D(\registers[791][2] ), .S0(n7494), .S1(n7734), 
        .Y(n5405) );
  MX4X1 U5026 ( .A(\registers[772][2] ), .B(\registers[773][2] ), .C(
        \registers[774][2] ), .D(\registers[775][2] ), .S0(n7495), .S1(n7734), 
        .Y(n5410) );
  MX4X1 U5027 ( .A(\registers[820][2] ), .B(\registers[821][2] ), .C(
        \registers[822][2] ), .D(\registers[823][2] ), .S0(n7494), .S1(n7733), 
        .Y(n5395) );
  MX4X1 U5028 ( .A(\registers[804][2] ), .B(\registers[805][2] ), .C(
        \registers[806][2] ), .D(\registers[807][2] ), .S0(n7494), .S1(n7734), 
        .Y(n5400) );
  MX4X1 U5029 ( .A(\registers[980][2] ), .B(\registers[981][2] ), .C(
        \registers[982][2] ), .D(\registers[983][2] ), .S0(n7490), .S1(n7730), 
        .Y(n5342) );
  MX4X1 U5030 ( .A(\registers[964][2] ), .B(\registers[965][2] ), .C(
        \registers[966][2] ), .D(\registers[967][2] ), .S0(n7491), .S1(n7730), 
        .Y(n5347) );
  MX4X1 U5031 ( .A(\registers[1012][2] ), .B(\registers[1013][2] ), .C(
        \registers[1014][2] ), .D(\registers[1015][2] ), .S0(n7490), .S1(n7730), .Y(n5332) );
  MX4X1 U5032 ( .A(\registers[996][2] ), .B(\registers[997][2] ), .C(
        \registers[998][2] ), .D(\registers[999][2] ), .S0(n7490), .S1(n7730), 
        .Y(n5337) );
  MX4X1 U5033 ( .A(\registers[916][2] ), .B(\registers[917][2] ), .C(
        \registers[918][2] ), .D(\registers[919][2] ), .S0(n7492), .S1(n7731), 
        .Y(n5363) );
  MX4X1 U5034 ( .A(\registers[900][2] ), .B(\registers[901][2] ), .C(
        \registers[902][2] ), .D(\registers[903][2] ), .S0(n7492), .S1(n7732), 
        .Y(n5368) );
  MX4X1 U5035 ( .A(\registers[948][2] ), .B(\registers[949][2] ), .C(
        \registers[950][2] ), .D(\registers[951][2] ), .S0(n7491), .S1(n7731), 
        .Y(n5353) );
  MX4X1 U5036 ( .A(\registers[932][2] ), .B(\registers[933][2] ), .C(
        \registers[934][2] ), .D(\registers[935][2] ), .S0(n7491), .S1(n7731), 
        .Y(n5358) );
  MX4X1 U5037 ( .A(\registers[596][2] ), .B(\registers[597][2] ), .C(
        \registers[598][2] ), .D(\registers[599][2] ), .S0(n7498), .S1(n7738), 
        .Y(n5469) );
  MX4X1 U5038 ( .A(\registers[580][2] ), .B(\registers[581][2] ), .C(
        \registers[582][2] ), .D(\registers[583][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5474) );
  MX4X1 U5039 ( .A(\registers[628][2] ), .B(\registers[629][2] ), .C(
        \registers[630][2] ), .D(\registers[631][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5459) );
  MX4X1 U5040 ( .A(\registers[612][2] ), .B(\registers[613][2] ), .C(
        \registers[614][2] ), .D(\registers[615][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5464) );
  MX4X1 U5041 ( .A(\registers[532][2] ), .B(\registers[533][2] ), .C(
        \registers[534][2] ), .D(\registers[535][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5490) );
  MX4X1 U5042 ( .A(\registers[516][2] ), .B(\registers[517][2] ), .C(
        \registers[518][2] ), .D(\registers[519][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5495) );
  MX4X1 U5043 ( .A(\registers[564][2] ), .B(\registers[565][2] ), .C(
        \registers[566][2] ), .D(\registers[567][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5480) );
  MX4X1 U5044 ( .A(\registers[548][2] ), .B(\registers[549][2] ), .C(
        \registers[550][2] ), .D(\registers[551][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5485) );
  MX4X1 U5045 ( .A(\registers[724][2] ), .B(\registers[725][2] ), .C(
        \registers[726][2] ), .D(\registers[727][2] ), .S0(n7496), .S1(n7735), 
        .Y(n5427) );
  MX4X1 U5046 ( .A(\registers[708][2] ), .B(\registers[709][2] ), .C(
        \registers[710][2] ), .D(\registers[711][2] ), .S0(n7496), .S1(n7735), 
        .Y(n5432) );
  MX4X1 U5047 ( .A(\registers[756][2] ), .B(\registers[757][2] ), .C(
        \registers[758][2] ), .D(\registers[759][2] ), .S0(n7495), .S1(n7734), 
        .Y(n5417) );
  MX4X1 U5048 ( .A(\registers[740][2] ), .B(\registers[741][2] ), .C(
        \registers[742][2] ), .D(\registers[743][2] ), .S0(n7495), .S1(n7735), 
        .Y(n5422) );
  MX4X1 U5049 ( .A(\registers[660][2] ), .B(\registers[661][2] ), .C(
        \registers[662][2] ), .D(\registers[663][2] ), .S0(n7497), .S1(n7736), 
        .Y(n5448) );
  MX4X1 U5050 ( .A(\registers[644][2] ), .B(\registers[645][2] ), .C(
        \registers[646][2] ), .D(\registers[647][2] ), .S0(n7497), .S1(n7737), 
        .Y(n5453) );
  MX4X1 U5051 ( .A(\registers[692][2] ), .B(\registers[693][2] ), .C(
        \registers[694][2] ), .D(\registers[695][2] ), .S0(n7496), .S1(n7736), 
        .Y(n5438) );
  MX4X1 U5052 ( .A(\registers[676][2] ), .B(\registers[677][2] ), .C(
        \registers[678][2] ), .D(\registers[679][2] ), .S0(n7497), .S1(n7736), 
        .Y(n5443) );
  MX4X1 U5053 ( .A(\registers[340][3] ), .B(\registers[341][3] ), .C(
        \registers[342][3] ), .D(\registers[343][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5894) );
  MX4X1 U5054 ( .A(\registers[324][3] ), .B(\registers[325][3] ), .C(
        \registers[326][3] ), .D(\registers[327][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5899) );
  MX4X1 U5055 ( .A(\registers[372][3] ), .B(\registers[373][3] ), .C(
        \registers[374][3] ), .D(\registers[375][3] ), .S0(n7524), .S1(n7762), 
        .Y(n5884) );
  MX4X1 U5056 ( .A(\registers[356][3] ), .B(\registers[357][3] ), .C(
        \registers[358][3] ), .D(\registers[359][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5889) );
  MX4X1 U5057 ( .A(\registers[276][3] ), .B(\registers[277][3] ), .C(
        \registers[278][3] ), .D(\registers[279][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5915) );
  MX4X1 U5058 ( .A(\registers[260][3] ), .B(\registers[261][3] ), .C(
        \registers[262][3] ), .D(\registers[263][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5920) );
  MX4X1 U5059 ( .A(\registers[308][3] ), .B(\registers[309][3] ), .C(
        \registers[310][3] ), .D(\registers[311][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5905) );
  MX4X1 U5060 ( .A(\registers[292][3] ), .B(\registers[293][3] ), .C(
        \registers[294][3] ), .D(\registers[295][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5910) );
  MX4X1 U5061 ( .A(\registers[468][3] ), .B(\registers[469][3] ), .C(
        \registers[470][3] ), .D(\registers[471][3] ), .S0(n7522), .S1(n7760), 
        .Y(n5852) );
  MX4X1 U5062 ( .A(\registers[452][3] ), .B(\registers[453][3] ), .C(
        \registers[454][3] ), .D(\registers[455][3] ), .S0(n7523), .S1(n7760), 
        .Y(n5857) );
  MX4X1 U5063 ( .A(\registers[500][3] ), .B(\registers[501][3] ), .C(
        \registers[502][3] ), .D(\registers[503][3] ), .S0(n7522), .S1(n7759), 
        .Y(n5842) );
  MX4X1 U5064 ( .A(\registers[484][3] ), .B(\registers[485][3] ), .C(
        \registers[486][3] ), .D(\registers[487][3] ), .S0(n7522), .S1(n7759), 
        .Y(n5847) );
  MX4X1 U5065 ( .A(\registers[404][3] ), .B(\registers[405][3] ), .C(
        \registers[406][3] ), .D(\registers[407][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5873) );
  MX4X1 U5066 ( .A(\registers[388][3] ), .B(\registers[389][3] ), .C(
        \registers[390][3] ), .D(\registers[391][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5878) );
  MX4X1 U5067 ( .A(\registers[436][3] ), .B(\registers[437][3] ), .C(
        \registers[438][3] ), .D(\registers[439][3] ), .S0(n7523), .S1(n7760), 
        .Y(n5863) );
  MX4X1 U5068 ( .A(\registers[420][3] ), .B(\registers[421][3] ), .C(
        \registers[422][3] ), .D(\registers[423][3] ), .S0(n7523), .S1(n7761), 
        .Y(n5868) );
  MX4X1 U5069 ( .A(\registers[84][3] ), .B(\registers[85][3] ), .C(
        \registers[86][3] ), .D(\registers[87][3] ), .S0(n7530), .S1(n7767), 
        .Y(n5979) );
  MX4X1 U5070 ( .A(\registers[68][3] ), .B(\registers[69][3] ), .C(
        \registers[70][3] ), .D(\registers[71][3] ), .S0(n7531), .S1(n7767), 
        .Y(n5984) );
  MX4X1 U5071 ( .A(\registers[116][3] ), .B(\registers[117][3] ), .C(
        \registers[118][3] ), .D(\registers[119][3] ), .S0(n7530), .S1(n7766), 
        .Y(n5969) );
  MX4X1 U5072 ( .A(\registers[100][3] ), .B(\registers[101][3] ), .C(
        \registers[102][3] ), .D(\registers[103][3] ), .S0(n7530), .S1(n7767), 
        .Y(n5974) );
  MX4X1 U5073 ( .A(\registers[20][3] ), .B(\registers[21][3] ), .C(
        \registers[22][3] ), .D(\registers[23][3] ), .S0(n7532), .S1(n7768), 
        .Y(n6000) );
  MX4X1 U5074 ( .A(\registers[4][3] ), .B(\registers[5][3] ), .C(
        \registers[6][3] ), .D(\registers[7][3] ), .S0(n7532), .S1(n7769), .Y(
        n6005) );
  MX4X1 U5075 ( .A(\registers[52][3] ), .B(\registers[53][3] ), .C(
        \registers[54][3] ), .D(\registers[55][3] ), .S0(n7531), .S1(n7768), 
        .Y(n5990) );
  MX4X1 U5076 ( .A(\registers[36][3] ), .B(\registers[37][3] ), .C(
        \registers[38][3] ), .D(\registers[39][3] ), .S0(n7531), .S1(n7768), 
        .Y(n5995) );
  MX4X1 U5077 ( .A(\registers[212][3] ), .B(\registers[213][3] ), .C(
        \registers[214][3] ), .D(\registers[215][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5937) );
  MX4X1 U5078 ( .A(\registers[196][3] ), .B(\registers[197][3] ), .C(
        \registers[198][3] ), .D(\registers[199][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5942) );
  MX4X1 U5079 ( .A(\registers[244][3] ), .B(\registers[245][3] ), .C(
        \registers[246][3] ), .D(\registers[247][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5927) );
  MX4X1 U5080 ( .A(\registers[228][3] ), .B(\registers[229][3] ), .C(
        \registers[230][3] ), .D(\registers[231][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5932) );
  MX4X1 U5081 ( .A(\registers[148][3] ), .B(\registers[149][3] ), .C(
        \registers[150][3] ), .D(\registers[151][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5958) );
  MX4X1 U5082 ( .A(\registers[132][3] ), .B(\registers[133][3] ), .C(
        \registers[134][3] ), .D(\registers[135][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5963) );
  MX4X1 U5083 ( .A(\registers[180][3] ), .B(\registers[181][3] ), .C(
        \registers[182][3] ), .D(\registers[183][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5948) );
  MX4X1 U5084 ( .A(\registers[164][3] ), .B(\registers[165][3] ), .C(
        \registers[166][3] ), .D(\registers[167][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5953) );
  MX4X1 U5085 ( .A(\registers[852][3] ), .B(\registers[853][3] ), .C(
        \registers[854][3] ), .D(\registers[855][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5724) );
  MX4X1 U5086 ( .A(\registers[836][3] ), .B(\registers[837][3] ), .C(
        \registers[838][3] ), .D(\registers[839][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5729) );
  MX4X1 U5087 ( .A(\registers[884][3] ), .B(\registers[885][3] ), .C(
        \registers[886][3] ), .D(\registers[887][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5714) );
  MX4X1 U5088 ( .A(\registers[868][3] ), .B(\registers[869][3] ), .C(
        \registers[870][3] ), .D(\registers[871][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5719) );
  MX4X1 U5089 ( .A(\registers[788][3] ), .B(\registers[789][3] ), .C(
        \registers[790][3] ), .D(\registers[791][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5745) );
  MX4X1 U5090 ( .A(\registers[772][3] ), .B(\registers[773][3] ), .C(
        \registers[774][3] ), .D(\registers[775][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5750) );
  MX4X1 U5091 ( .A(\registers[820][3] ), .B(\registers[821][3] ), .C(
        \registers[822][3] ), .D(\registers[823][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5735) );
  MX4X1 U5092 ( .A(\registers[804][3] ), .B(\registers[805][3] ), .C(
        \registers[806][3] ), .D(\registers[807][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5740) );
  MX4X1 U5093 ( .A(\registers[980][3] ), .B(\registers[981][3] ), .C(
        \registers[982][3] ), .D(\registers[983][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5682) );
  MX4X1 U5094 ( .A(\registers[964][3] ), .B(\registers[965][3] ), .C(
        \registers[966][3] ), .D(\registers[967][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5687) );
  MX4X1 U5095 ( .A(\registers[1012][3] ), .B(\registers[1013][3] ), .C(
        \registers[1014][3] ), .D(\registers[1015][3] ), .S0(n7511), .S1(n7749), .Y(n5672) );
  MX4X1 U5096 ( .A(\registers[996][3] ), .B(\registers[997][3] ), .C(
        \registers[998][3] ), .D(\registers[999][3] ), .S0(n7511), .S1(n7750), 
        .Y(n5677) );
  MX4X1 U5097 ( .A(\registers[916][3] ), .B(\registers[917][3] ), .C(
        \registers[918][3] ), .D(\registers[919][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5703) );
  MX4X1 U5098 ( .A(\registers[900][3] ), .B(\registers[901][3] ), .C(
        \registers[902][3] ), .D(\registers[903][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5708) );
  MX4X1 U5099 ( .A(\registers[948][3] ), .B(\registers[949][3] ), .C(
        \registers[950][3] ), .D(\registers[951][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5693) );
  MX4X1 U5100 ( .A(\registers[932][3] ), .B(\registers[933][3] ), .C(
        \registers[934][3] ), .D(\registers[935][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5698) );
  MX4X1 U5101 ( .A(\registers[596][3] ), .B(\registers[597][3] ), .C(
        \registers[598][3] ), .D(\registers[599][3] ), .S0(n7520), .S1(n7757), 
        .Y(n5809) );
  MX4X1 U5102 ( .A(\registers[580][3] ), .B(\registers[581][3] ), .C(
        \registers[582][3] ), .D(\registers[583][3] ), .S0(n7520), .S1(n7758), 
        .Y(n5814) );
  MX4X1 U5103 ( .A(\registers[628][3] ), .B(\registers[629][3] ), .C(
        \registers[630][3] ), .D(\registers[631][3] ), .S0(n7519), .S1(n7757), 
        .Y(n5799) );
  MX4X1 U5104 ( .A(\registers[612][3] ), .B(\registers[613][3] ), .C(
        \registers[614][3] ), .D(\registers[615][3] ), .S0(n7519), .S1(n7757), 
        .Y(n5804) );
  MX4X1 U5105 ( .A(\registers[532][3] ), .B(\registers[533][3] ), .C(
        \registers[534][3] ), .D(\registers[535][3] ), .S0(n7521), .S1(n7758), 
        .Y(n5830) );
  MX4X1 U5106 ( .A(\registers[516][3] ), .B(\registers[517][3] ), .C(
        \registers[518][3] ), .D(\registers[519][3] ), .S0(n7521), .S1(n7759), 
        .Y(n5835) );
  MX4X1 U5107 ( .A(\registers[564][3] ), .B(\registers[565][3] ), .C(
        \registers[566][3] ), .D(\registers[567][3] ), .S0(n7520), .S1(n7758), 
        .Y(n5820) );
  MX4X1 U5108 ( .A(\registers[548][3] ), .B(\registers[549][3] ), .C(
        \registers[550][3] ), .D(\registers[551][3] ), .S0(n7521), .S1(n7758), 
        .Y(n5825) );
  MX4X1 U5109 ( .A(\registers[724][3] ), .B(\registers[725][3] ), .C(
        \registers[726][3] ), .D(\registers[727][3] ), .S0(n7517), .S1(n7755), 
        .Y(n5767) );
  MX4X1 U5110 ( .A(\registers[708][3] ), .B(\registers[709][3] ), .C(
        \registers[710][3] ), .D(\registers[711][3] ), .S0(n7517), .S1(n7755), 
        .Y(n5772) );
  MX4X1 U5111 ( .A(\registers[756][3] ), .B(\registers[757][3] ), .C(
        \registers[758][3] ), .D(\registers[759][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5757) );
  MX4X1 U5112 ( .A(\registers[740][3] ), .B(\registers[741][3] ), .C(
        \registers[742][3] ), .D(\registers[743][3] ), .S0(n7517), .S1(n7754), 
        .Y(n5762) );
  MX4X1 U5113 ( .A(\registers[660][3] ), .B(\registers[661][3] ), .C(
        \registers[662][3] ), .D(\registers[663][3] ), .S0(n7518), .S1(n7756), 
        .Y(n5788) );
  MX4X1 U5114 ( .A(\registers[644][3] ), .B(\registers[645][3] ), .C(
        \registers[646][3] ), .D(\registers[647][3] ), .S0(n7519), .S1(n7756), 
        .Y(n5793) );
  MX4X1 U5115 ( .A(\registers[692][3] ), .B(\registers[693][3] ), .C(
        \registers[694][3] ), .D(\registers[695][3] ), .S0(n7518), .S1(n7755), 
        .Y(n5778) );
  MX4X1 U5116 ( .A(\registers[676][3] ), .B(\registers[677][3] ), .C(
        \registers[678][3] ), .D(\registers[679][3] ), .S0(n7518), .S1(n7756), 
        .Y(n5783) );
  MX4X1 U5117 ( .A(\registers[340][4] ), .B(\registers[341][4] ), .C(
        \registers[342][4] ), .D(\registers[343][4] ), .S0(n7546), .S1(n7782), 
        .Y(n6234) );
  MX4X1 U5118 ( .A(\registers[324][4] ), .B(\registers[325][4] ), .C(
        \registers[326][4] ), .D(\registers[327][4] ), .S0(n7547), .S1(n7782), 
        .Y(n6239) );
  MX4X1 U5119 ( .A(\registers[372][4] ), .B(\registers[373][4] ), .C(
        \registers[374][4] ), .D(\registers[375][4] ), .S0(n7546), .S1(n7781), 
        .Y(n6224) );
  MX4X1 U5120 ( .A(\registers[356][4] ), .B(\registers[357][4] ), .C(
        \registers[358][4] ), .D(\registers[359][4] ), .S0(n7546), .S1(n7782), 
        .Y(n6229) );
  MX4X1 U5121 ( .A(\registers[276][4] ), .B(\registers[277][4] ), .C(
        \registers[278][4] ), .D(\registers[279][4] ), .S0(n7548), .S1(n7783), 
        .Y(n6255) );
  MX4X1 U5122 ( .A(\registers[260][4] ), .B(\registers[261][4] ), .C(
        \registers[262][4] ), .D(\registers[263][4] ), .S0(n7548), .S1(n7783), 
        .Y(n6260) );
  MX4X1 U5123 ( .A(\registers[308][4] ), .B(\registers[309][4] ), .C(
        \registers[310][4] ), .D(\registers[311][4] ), .S0(n7547), .S1(n7782), 
        .Y(n6245) );
  MX4X1 U5124 ( .A(\registers[292][4] ), .B(\registers[293][4] ), .C(
        \registers[294][4] ), .D(\registers[295][4] ), .S0(n7547), .S1(n7783), 
        .Y(n6250) );
  MX4X1 U5125 ( .A(\registers[468][4] ), .B(\registers[469][4] ), .C(
        \registers[470][4] ), .D(\registers[471][4] ), .S0(n7544), .S1(n7779), 
        .Y(n6192) );
  MX4X1 U5126 ( .A(\registers[452][4] ), .B(\registers[453][4] ), .C(
        \registers[454][4] ), .D(\registers[455][4] ), .S0(n7544), .S1(n7780), 
        .Y(n6197) );
  MX4X1 U5127 ( .A(\registers[500][4] ), .B(\registers[501][4] ), .C(
        \registers[502][4] ), .D(\registers[503][4] ), .S0(n7543), .S1(n7779), 
        .Y(n6182) );
  MX4X1 U5128 ( .A(\registers[484][4] ), .B(\registers[485][4] ), .C(
        \registers[486][4] ), .D(\registers[487][4] ), .S0(n7543), .S1(n7779), 
        .Y(n6187) );
  MX4X1 U5129 ( .A(\registers[404][4] ), .B(\registers[405][4] ), .C(
        \registers[406][4] ), .D(\registers[407][4] ), .S0(n7545), .S1(n7781), 
        .Y(n6213) );
  MX4X1 U5130 ( .A(\registers[388][4] ), .B(\registers[389][4] ), .C(
        \registers[390][4] ), .D(\registers[391][4] ), .S0(n7545), .S1(n7781), 
        .Y(n6218) );
  MX4X1 U5131 ( .A(\registers[436][4] ), .B(\registers[437][4] ), .C(
        \registers[438][4] ), .D(\registers[439][4] ), .S0(n7544), .S1(n7780), 
        .Y(n6203) );
  MX4X1 U5132 ( .A(\registers[420][4] ), .B(\registers[421][4] ), .C(
        \registers[422][4] ), .D(\registers[423][4] ), .S0(n7545), .S1(n7780), 
        .Y(n6208) );
  MX4X1 U5133 ( .A(\registers[84][4] ), .B(\registers[85][4] ), .C(
        \registers[86][4] ), .D(\registers[87][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6319) );
  MX4X1 U5134 ( .A(\registers[68][4] ), .B(\registers[69][4] ), .C(
        \registers[70][4] ), .D(\registers[71][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6324) );
  MX4X1 U5135 ( .A(\registers[116][4] ), .B(\registers[117][4] ), .C(
        \registers[118][4] ), .D(\registers[119][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6309) );
  MX4X1 U5136 ( .A(\registers[100][4] ), .B(\registers[101][4] ), .C(
        \registers[102][4] ), .D(\registers[103][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6314) );
  MX4X1 U5137 ( .A(\registers[20][4] ), .B(\registers[21][4] ), .C(
        \registers[22][4] ), .D(\registers[23][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6340) );
  MX4X1 U5138 ( .A(\registers[4][4] ), .B(\registers[5][4] ), .C(
        \registers[6][4] ), .D(\registers[7][4] ), .S0(n7553), .S1(n7788), .Y(
        n6345) );
  MX4X1 U5139 ( .A(\registers[52][4] ), .B(\registers[53][4] ), .C(
        \registers[54][4] ), .D(\registers[55][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6330) );
  MX4X1 U5140 ( .A(\registers[36][4] ), .B(\registers[37][4] ), .C(
        \registers[38][4] ), .D(\registers[39][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6335) );
  MX4X1 U5141 ( .A(\registers[212][4] ), .B(\registers[213][4] ), .C(
        \registers[214][4] ), .D(\registers[215][4] ), .S0(n7549), .S1(n7784), 
        .Y(n6277) );
  MX4X1 U5142 ( .A(\registers[196][4] ), .B(\registers[197][4] ), .C(
        \registers[198][4] ), .D(\registers[199][4] ), .S0(n7549), .S1(n7785), 
        .Y(n6282) );
  MX4X1 U5143 ( .A(\registers[244][4] ), .B(\registers[245][4] ), .C(
        \registers[246][4] ), .D(\registers[247][4] ), .S0(n7548), .S1(n7784), 
        .Y(n6267) );
  MX4X1 U5144 ( .A(\registers[228][4] ), .B(\registers[229][4] ), .C(
        \registers[230][4] ), .D(\registers[231][4] ), .S0(n7549), .S1(n7784), 
        .Y(n6272) );
  MX4X1 U5145 ( .A(\registers[148][4] ), .B(\registers[149][4] ), .C(
        \registers[150][4] ), .D(\registers[151][4] ), .S0(n7550), .S1(n7786), 
        .Y(n6298) );
  MX4X1 U5146 ( .A(\registers[132][4] ), .B(\registers[133][4] ), .C(
        \registers[134][4] ), .D(\registers[135][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6303) );
  MX4X1 U5147 ( .A(\registers[180][4] ), .B(\registers[181][4] ), .C(
        \registers[182][4] ), .D(\registers[183][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6288) );
  MX4X1 U5148 ( .A(\registers[164][4] ), .B(\registers[165][4] ), .C(
        \registers[166][4] ), .D(\registers[167][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6293) );
  MX4X1 U5149 ( .A(\registers[852][4] ), .B(\registers[853][4] ), .C(
        \registers[854][4] ), .D(\registers[855][4] ), .S0(n7536), .S1(n7772), 
        .Y(n6064) );
  MX4X1 U5150 ( .A(\registers[836][4] ), .B(\registers[837][4] ), .C(
        \registers[838][4] ), .D(\registers[839][4] ), .S0(n7536), .S1(n7772), 
        .Y(n6069) );
  MX4X1 U5151 ( .A(\registers[884][4] ), .B(\registers[885][4] ), .C(
        \registers[886][4] ), .D(\registers[887][4] ), .S0(n7535), .S1(n7771), 
        .Y(n6054) );
  MX4X1 U5152 ( .A(\registers[868][4] ), .B(\registers[869][4] ), .C(
        \registers[870][4] ), .D(\registers[871][4] ), .S0(n7535), .S1(n7772), 
        .Y(n6059) );
  MX4X1 U5153 ( .A(\registers[788][4] ), .B(\registers[789][4] ), .C(
        \registers[790][4] ), .D(\registers[791][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6085) );
  MX4X1 U5154 ( .A(\registers[772][4] ), .B(\registers[773][4] ), .C(
        \registers[774][4] ), .D(\registers[775][4] ), .S0(n7537), .S1(n7774), 
        .Y(n6090) );
  MX4X1 U5155 ( .A(\registers[820][4] ), .B(\registers[821][4] ), .C(
        \registers[822][4] ), .D(\registers[823][4] ), .S0(n7536), .S1(n7773), 
        .Y(n6075) );
  MX4X1 U5156 ( .A(\registers[804][4] ), .B(\registers[805][4] ), .C(
        \registers[806][4] ), .D(\registers[807][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6080) );
  MX4X1 U5157 ( .A(\registers[980][4] ), .B(\registers[981][4] ), .C(
        \registers[982][4] ), .D(\registers[983][4] ), .S0(n7533), .S1(n7770), 
        .Y(n6022) );
  MX4X1 U5158 ( .A(\registers[964][4] ), .B(\registers[965][4] ), .C(
        \registers[966][4] ), .D(\registers[967][4] ), .S0(n7533), .S1(n7770), 
        .Y(n6027) );
  MX4X1 U5159 ( .A(\registers[1012][4] ), .B(\registers[1013][4] ), .C(
        \registers[1014][4] ), .D(\registers[1015][4] ), .S0(n7532), .S1(n7769), .Y(n6012) );
  MX4X1 U5160 ( .A(\registers[996][4] ), .B(\registers[997][4] ), .C(
        \registers[998][4] ), .D(\registers[999][4] ), .S0(n7533), .S1(n7769), 
        .Y(n6017) );
  MX4X1 U5161 ( .A(\registers[916][4] ), .B(\registers[917][4] ), .C(
        \registers[918][4] ), .D(\registers[919][4] ), .S0(n7534), .S1(n7771), 
        .Y(n6043) );
  MX4X1 U5162 ( .A(\registers[900][4] ), .B(\registers[901][4] ), .C(
        \registers[902][4] ), .D(\registers[903][4] ), .S0(n7535), .S1(n7771), 
        .Y(n6048) );
  MX4X1 U5163 ( .A(\registers[948][4] ), .B(\registers[949][4] ), .C(
        \registers[950][4] ), .D(\registers[951][4] ), .S0(n7534), .S1(n7770), 
        .Y(n6033) );
  MX4X1 U5164 ( .A(\registers[932][4] ), .B(\registers[933][4] ), .C(
        \registers[934][4] ), .D(\registers[935][4] ), .S0(n7534), .S1(n7770), 
        .Y(n6038) );
  MX4X1 U5165 ( .A(\registers[596][4] ), .B(\registers[597][4] ), .C(
        \registers[598][4] ), .D(\registers[599][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6149) );
  MX4X1 U5166 ( .A(\registers[580][4] ), .B(\registers[581][4] ), .C(
        \registers[582][4] ), .D(\registers[583][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6154) );
  MX4X1 U5167 ( .A(\registers[628][4] ), .B(\registers[629][4] ), .C(
        \registers[630][4] ), .D(\registers[631][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6139) );
  MX4X1 U5168 ( .A(\registers[612][4] ), .B(\registers[613][4] ), .C(
        \registers[614][4] ), .D(\registers[615][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6144) );
  MX4X1 U5169 ( .A(\registers[532][4] ), .B(\registers[533][4] ), .C(
        \registers[534][4] ), .D(\registers[535][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6170) );
  MX4X1 U5170 ( .A(\registers[516][4] ), .B(\registers[517][4] ), .C(
        \registers[518][4] ), .D(\registers[519][4] ), .S0(n7543), .S1(n7778), 
        .Y(n6175) );
  MX4X1 U5171 ( .A(\registers[564][4] ), .B(\registers[565][4] ), .C(
        \registers[566][4] ), .D(\registers[567][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6160) );
  MX4X1 U5172 ( .A(\registers[548][4] ), .B(\registers[549][4] ), .C(
        \registers[550][4] ), .D(\registers[551][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6165) );
  MX4X1 U5173 ( .A(\registers[724][4] ), .B(\registers[725][4] ), .C(
        \registers[726][4] ), .D(\registers[727][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6107) );
  MX4X1 U5174 ( .A(\registers[708][4] ), .B(\registers[709][4] ), .C(
        \registers[710][4] ), .D(\registers[711][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6112) );
  MX4X1 U5175 ( .A(\registers[756][4] ), .B(\registers[757][4] ), .C(
        \registers[758][4] ), .D(\registers[759][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6097) );
  MX4X1 U5176 ( .A(\registers[740][4] ), .B(\registers[741][4] ), .C(
        \registers[742][4] ), .D(\registers[743][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6102) );
  MX4X1 U5177 ( .A(\registers[660][4] ), .B(\registers[661][4] ), .C(
        \registers[662][4] ), .D(\registers[663][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6128) );
  MX4X1 U5178 ( .A(\registers[644][4] ), .B(\registers[645][4] ), .C(
        \registers[646][4] ), .D(\registers[647][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6133) );
  MX4X1 U5179 ( .A(\registers[692][4] ), .B(\registers[693][4] ), .C(
        \registers[694][4] ), .D(\registers[695][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6118) );
  MX4X1 U5180 ( .A(\registers[676][4] ), .B(\registers[677][4] ), .C(
        \registers[678][4] ), .D(\registers[679][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6123) );
  MX4X1 U5181 ( .A(\registers[340][5] ), .B(\registers[341][5] ), .C(
        \registers[342][5] ), .D(\registers[343][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6574) );
  MX4X1 U5182 ( .A(\registers[324][5] ), .B(\registers[325][5] ), .C(
        \registers[326][5] ), .D(\registers[327][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6579) );
  MX4X1 U5183 ( .A(\registers[372][5] ), .B(\registers[373][5] ), .C(
        \registers[374][5] ), .D(\registers[375][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6564) );
  MX4X1 U5184 ( .A(\registers[356][5] ), .B(\registers[357][5] ), .C(
        \registers[358][5] ), .D(\registers[359][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6569) );
  MX4X1 U5185 ( .A(\registers[276][5] ), .B(\registers[277][5] ), .C(
        \registers[278][5] ), .D(\registers[279][5] ), .S0(n7569), .S1(n7803), 
        .Y(n6595) );
  MX4X1 U5186 ( .A(\registers[260][5] ), .B(\registers[261][5] ), .C(
        \registers[262][5] ), .D(\registers[263][5] ), .S0(n7569), .S1(n7803), 
        .Y(n6600) );
  MX4X1 U5187 ( .A(\registers[308][5] ), .B(\registers[309][5] ), .C(
        \registers[310][5] ), .D(\registers[311][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6585) );
  MX4X1 U5188 ( .A(\registers[292][5] ), .B(\registers[293][5] ), .C(
        \registers[294][5] ), .D(\registers[295][5] ), .S0(n7569), .S1(n7802), 
        .Y(n6590) );
  MX4X1 U5189 ( .A(\registers[468][5] ), .B(\registers[469][5] ), .C(
        \registers[470][5] ), .D(\registers[471][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6532) );
  MX4X1 U5190 ( .A(\registers[452][5] ), .B(\registers[453][5] ), .C(
        \registers[454][5] ), .D(\registers[455][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6537) );
  MX4X1 U5191 ( .A(\registers[500][5] ), .B(\registers[501][5] ), .C(
        \registers[502][5] ), .D(\registers[503][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6522) );
  MX4X1 U5192 ( .A(\registers[484][5] ), .B(\registers[485][5] ), .C(
        \registers[486][5] ), .D(\registers[487][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6527) );
  MX4X1 U5193 ( .A(\registers[404][5] ), .B(\registers[405][5] ), .C(
        \registers[406][5] ), .D(\registers[407][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6553) );
  MX4X1 U5194 ( .A(\registers[388][5] ), .B(\registers[389][5] ), .C(
        \registers[390][5] ), .D(\registers[391][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6558) );
  MX4X1 U5195 ( .A(\registers[436][5] ), .B(\registers[437][5] ), .C(
        \registers[438][5] ), .D(\registers[439][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6543) );
  MX4X1 U5196 ( .A(\registers[420][5] ), .B(\registers[421][5] ), .C(
        \registers[422][5] ), .D(\registers[423][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6548) );
  MX4X1 U5197 ( .A(\registers[84][5] ), .B(\registers[85][5] ), .C(
        \registers[86][5] ), .D(\registers[87][5] ), .S0(n7573), .S1(n7805), 
        .Y(n6659) );
  MX4X1 U5198 ( .A(\registers[68][5] ), .B(\registers[69][5] ), .C(
        \registers[70][5] ), .D(\registers[71][5] ), .S0(n7573), .S1(n7806), 
        .Y(n6664) );
  MX4X1 U5199 ( .A(\registers[116][5] ), .B(\registers[117][5] ), .C(
        \registers[118][5] ), .D(\registers[119][5] ), .S0(n7572), .S1(n7805), 
        .Y(n6649) );
  MX4X1 U5200 ( .A(\registers[100][5] ), .B(\registers[101][5] ), .C(
        \registers[102][5] ), .D(\registers[103][5] ), .S0(n7573), .S1(n7805), 
        .Y(n6654) );
  MX4X1 U5201 ( .A(\registers[20][5] ), .B(\registers[21][5] ), .C(
        \registers[22][5] ), .D(\registers[23][5] ), .S0(n7574), .S1(n7807), 
        .Y(n6680) );
  MX4X1 U5202 ( .A(\registers[4][5] ), .B(\registers[5][5] ), .C(
        \registers[6][5] ), .D(\registers[7][5] ), .S0(n7575), .S1(n7807), .Y(
        n6685) );
  MX4X1 U5203 ( .A(\registers[52][5] ), .B(\registers[53][5] ), .C(
        \registers[54][5] ), .D(\registers[55][5] ), .S0(n7574), .S1(n7806), 
        .Y(n6670) );
  MX4X1 U5204 ( .A(\registers[36][5] ), .B(\registers[37][5] ), .C(
        \registers[38][5] ), .D(\registers[39][5] ), .S0(n7574), .S1(n7806), 
        .Y(n6675) );
  MX4X1 U5205 ( .A(\registers[212][5] ), .B(\registers[213][5] ), .C(
        \registers[214][5] ), .D(\registers[215][5] ), .S0(n7570), .S1(n7703), 
        .Y(n6617) );
  MX4X1 U5206 ( .A(\registers[196][5] ), .B(\registers[197][5] ), .C(
        \registers[198][5] ), .D(\registers[199][5] ), .S0(n7571), .S1(n7701), 
        .Y(n6622) );
  MX4X1 U5207 ( .A(\registers[244][5] ), .B(\registers[245][5] ), .C(
        \registers[246][5] ), .D(\registers[247][5] ), .S0(n7570), .S1(n7803), 
        .Y(n6607) );
  MX4X1 U5208 ( .A(\registers[228][5] ), .B(\registers[229][5] ), .C(
        \registers[230][5] ), .D(\registers[231][5] ), .S0(n7570), .S1(n7698), 
        .Y(n6612) );
  MX4X1 U5209 ( .A(\registers[148][5] ), .B(\registers[149][5] ), .C(
        \registers[150][5] ), .D(\registers[151][5] ), .S0(n7572), .S1(n7804), 
        .Y(n6638) );
  MX4X1 U5210 ( .A(\registers[132][5] ), .B(\registers[133][5] ), .C(
        \registers[134][5] ), .D(\registers[135][5] ), .S0(n7572), .S1(n7805), 
        .Y(n6643) );
  MX4X1 U5211 ( .A(\registers[180][5] ), .B(\registers[181][5] ), .C(
        \registers[182][5] ), .D(\registers[183][5] ), .S0(n7571), .S1(n7804), 
        .Y(n6628) );
  MX4X1 U5212 ( .A(\registers[164][5] ), .B(\registers[165][5] ), .C(
        \registers[166][5] ), .D(\registers[167][5] ), .S0(n7571), .S1(n7804), 
        .Y(n6633) );
  MX4X1 U5213 ( .A(\registers[852][5] ), .B(\registers[853][5] ), .C(
        \registers[854][5] ), .D(\registers[855][5] ), .S0(n7557), .S1(n7792), 
        .Y(n6404) );
  MX4X1 U5214 ( .A(\registers[836][5] ), .B(\registers[837][5] ), .C(
        \registers[838][5] ), .D(\registers[839][5] ), .S0(n7557), .S1(n7792), 
        .Y(n6409) );
  MX4X1 U5215 ( .A(\registers[884][5] ), .B(\registers[885][5] ), .C(
        \registers[886][5] ), .D(\registers[887][5] ), .S0(n7556), .S1(n7791), 
        .Y(n6394) );
  MX4X1 U5216 ( .A(\registers[868][5] ), .B(\registers[869][5] ), .C(
        \registers[870][5] ), .D(\registers[871][5] ), .S0(n7557), .S1(n7791), 
        .Y(n6399) );
  MX4X1 U5217 ( .A(\registers[788][5] ), .B(\registers[789][5] ), .C(
        \registers[790][5] ), .D(\registers[791][5] ), .S0(n7558), .S1(n7793), 
        .Y(n6425) );
  MX4X1 U5218 ( .A(\registers[772][5] ), .B(\registers[773][5] ), .C(
        \registers[774][5] ), .D(\registers[775][5] ), .S0(n7559), .S1(n7793), 
        .Y(n6430) );
  MX4X1 U5219 ( .A(\registers[820][5] ), .B(\registers[821][5] ), .C(
        \registers[822][5] ), .D(\registers[823][5] ), .S0(n7558), .S1(n7792), 
        .Y(n6415) );
  MX4X1 U5220 ( .A(\registers[804][5] ), .B(\registers[805][5] ), .C(
        \registers[806][5] ), .D(\registers[807][5] ), .S0(n7558), .S1(n7793), 
        .Y(n6420) );
  MX4X1 U5221 ( .A(\registers[980][5] ), .B(\registers[981][5] ), .C(
        \registers[982][5] ), .D(\registers[983][5] ), .S0(n7554), .S1(n7789), 
        .Y(n6362) );
  MX4X1 U5222 ( .A(\registers[964][5] ), .B(\registers[965][5] ), .C(
        \registers[966][5] ), .D(\registers[967][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6367) );
  MX4X1 U5223 ( .A(\registers[1012][5] ), .B(\registers[1013][5] ), .C(
        \registers[1014][5] ), .D(\registers[1015][5] ), .S0(n7554), .S1(n7789), .Y(n6352) );
  MX4X1 U5224 ( .A(\registers[996][5] ), .B(\registers[997][5] ), .C(
        \registers[998][5] ), .D(\registers[999][5] ), .S0(n7554), .S1(n7789), 
        .Y(n6357) );
  MX4X1 U5225 ( .A(\registers[916][5] ), .B(\registers[917][5] ), .C(
        \registers[918][5] ), .D(\registers[919][5] ), .S0(n7556), .S1(n7790), 
        .Y(n6383) );
  MX4X1 U5226 ( .A(\registers[900][5] ), .B(\registers[901][5] ), .C(
        \registers[902][5] ), .D(\registers[903][5] ), .S0(n7556), .S1(n7791), 
        .Y(n6388) );
  MX4X1 U5227 ( .A(\registers[948][5] ), .B(\registers[949][5] ), .C(
        \registers[950][5] ), .D(\registers[951][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6373) );
  MX4X1 U5228 ( .A(\registers[932][5] ), .B(\registers[933][5] ), .C(
        \registers[934][5] ), .D(\registers[935][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6378) );
  MX4X1 U5229 ( .A(\registers[596][5] ), .B(\registers[597][5] ), .C(
        \registers[598][5] ), .D(\registers[599][5] ), .S0(n7562), .S1(n7797), 
        .Y(n6489) );
  MX4X1 U5230 ( .A(\registers[580][5] ), .B(\registers[581][5] ), .C(
        \registers[582][5] ), .D(\registers[583][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6494) );
  MX4X1 U5231 ( .A(\registers[628][5] ), .B(\registers[629][5] ), .C(
        \registers[630][5] ), .D(\registers[631][5] ), .S0(n7562), .S1(n7796), 
        .Y(n6479) );
  MX4X1 U5232 ( .A(\registers[612][5] ), .B(\registers[613][5] ), .C(
        \registers[614][5] ), .D(\registers[615][5] ), .S0(n7562), .S1(n7796), 
        .Y(n6484) );
  MX4X1 U5233 ( .A(\registers[532][5] ), .B(\registers[533][5] ), .C(
        \registers[534][5] ), .D(\registers[535][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6510) );
  MX4X1 U5234 ( .A(\registers[516][5] ), .B(\registers[517][5] ), .C(
        \registers[518][5] ), .D(\registers[519][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6515) );
  MX4X1 U5235 ( .A(\registers[564][5] ), .B(\registers[565][5] ), .C(
        \registers[566][5] ), .D(\registers[567][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6500) );
  MX4X1 U5236 ( .A(\registers[548][5] ), .B(\registers[549][5] ), .C(
        \registers[550][5] ), .D(\registers[551][5] ), .S0(n7563), .S1(n7798), 
        .Y(n6505) );
  MX4X1 U5237 ( .A(\registers[724][5] ), .B(\registers[725][5] ), .C(
        \registers[726][5] ), .D(\registers[727][5] ), .S0(n7560), .S1(n7794), 
        .Y(n6447) );
  MX4X1 U5238 ( .A(\registers[708][5] ), .B(\registers[709][5] ), .C(
        \registers[710][5] ), .D(\registers[711][5] ), .S0(n7560), .S1(n7794), 
        .Y(n6452) );
  MX4X1 U5239 ( .A(\registers[756][5] ), .B(\registers[757][5] ), .C(
        \registers[758][5] ), .D(\registers[759][5] ), .S0(n7559), .S1(n7794), 
        .Y(n6437) );
  MX4X1 U5240 ( .A(\registers[740][5] ), .B(\registers[741][5] ), .C(
        \registers[742][5] ), .D(\registers[743][5] ), .S0(n7559), .S1(n7794), 
        .Y(n6442) );
  MX4X1 U5241 ( .A(\registers[660][5] ), .B(\registers[661][5] ), .C(
        \registers[662][5] ), .D(\registers[663][5] ), .S0(n7561), .S1(n7795), 
        .Y(n6468) );
  MX4X1 U5242 ( .A(\registers[644][5] ), .B(\registers[645][5] ), .C(
        \registers[646][5] ), .D(\registers[647][5] ), .S0(n7561), .S1(n7796), 
        .Y(n6473) );
  MX4X1 U5243 ( .A(\registers[692][5] ), .B(\registers[693][5] ), .C(
        \registers[694][5] ), .D(\registers[695][5] ), .S0(n7560), .S1(n7795), 
        .Y(n6458) );
  MX4X1 U5244 ( .A(\registers[676][5] ), .B(\registers[677][5] ), .C(
        \registers[678][5] ), .D(\registers[679][5] ), .S0(n7561), .S1(n7795), 
        .Y(n6463) );
  MX4X1 U5245 ( .A(\registers[340][6] ), .B(\registers[341][6] ), .C(
        \registers[342][6] ), .D(\registers[343][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6914) );
  MX4X1 U5246 ( .A(\registers[324][6] ), .B(\registers[325][6] ), .C(
        \registers[326][6] ), .D(\registers[327][6] ), .S0(n7589), .S1(n7821), 
        .Y(n6919) );
  MX4X1 U5247 ( .A(\registers[372][6] ), .B(\registers[373][6] ), .C(
        \registers[374][6] ), .D(\registers[375][6] ), .S0(n7588), .S1(n7820), 
        .Y(n6904) );
  MX4X1 U5248 ( .A(\registers[356][6] ), .B(\registers[357][6] ), .C(
        \registers[358][6] ), .D(\registers[359][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6909) );
  MX4X1 U5249 ( .A(\registers[276][6] ), .B(\registers[277][6] ), .C(
        \registers[278][6] ), .D(\registers[279][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6935) );
  MX4X1 U5250 ( .A(\registers[260][6] ), .B(\registers[261][6] ), .C(
        \registers[262][6] ), .D(\registers[263][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6940) );
  MX4X1 U5251 ( .A(\registers[308][6] ), .B(\registers[309][6] ), .C(
        \registers[310][6] ), .D(\registers[311][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6925) );
  MX4X1 U5252 ( .A(\registers[292][6] ), .B(\registers[293][6] ), .C(
        \registers[294][6] ), .D(\registers[295][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6930) );
  MX4X1 U5253 ( .A(\registers[468][6] ), .B(\registers[469][6] ), .C(
        \registers[470][6] ), .D(\registers[471][6] ), .S0(n7586), .S1(n7818), 
        .Y(n6872) );
  MX4X1 U5254 ( .A(\registers[452][6] ), .B(\registers[453][6] ), .C(
        \registers[454][6] ), .D(\registers[455][6] ), .S0(n7587), .S1(n7818), 
        .Y(n6877) );
  MX4X1 U5255 ( .A(\registers[500][6] ), .B(\registers[501][6] ), .C(
        \registers[502][6] ), .D(\registers[503][6] ), .S0(n7586), .S1(n7817), 
        .Y(n6862) );
  MX4X1 U5256 ( .A(\registers[484][6] ), .B(\registers[485][6] ), .C(
        \registers[486][6] ), .D(\registers[487][6] ), .S0(n7586), .S1(n7817), 
        .Y(n6867) );
  MX4X1 U5257 ( .A(\registers[404][6] ), .B(\registers[405][6] ), .C(
        \registers[406][6] ), .D(\registers[407][6] ), .S0(n7588), .S1(n7819), 
        .Y(n6893) );
  MX4X1 U5258 ( .A(\registers[388][6] ), .B(\registers[389][6] ), .C(
        \registers[390][6] ), .D(\registers[391][6] ), .S0(n7588), .S1(n7819), 
        .Y(n6898) );
  MX4X1 U5259 ( .A(\registers[436][6] ), .B(\registers[437][6] ), .C(
        \registers[438][6] ), .D(\registers[439][6] ), .S0(n7587), .S1(n7818), 
        .Y(n6883) );
  MX4X1 U5260 ( .A(\registers[420][6] ), .B(\registers[421][6] ), .C(
        \registers[422][6] ), .D(\registers[423][6] ), .S0(n7587), .S1(n7819), 
        .Y(n6888) );
  MX4X1 U5261 ( .A(\registers[84][6] ), .B(\registers[85][6] ), .C(
        \registers[86][6] ), .D(\registers[87][6] ), .S0(n7594), .S1(n7825), 
        .Y(n6999) );
  MX4X1 U5262 ( .A(\registers[68][6] ), .B(\registers[69][6] ), .C(
        \registers[70][6] ), .D(\registers[71][6] ), .S0(n7595), .S1(n7825), 
        .Y(n7004) );
  MX4X1 U5263 ( .A(\registers[116][6] ), .B(\registers[117][6] ), .C(
        \registers[118][6] ), .D(\registers[119][6] ), .S0(n7594), .S1(n7825), 
        .Y(n6989) );
  MX4X1 U5264 ( .A(\registers[100][6] ), .B(\registers[101][6] ), .C(
        \registers[102][6] ), .D(\registers[103][6] ), .S0(n7594), .S1(n7825), 
        .Y(n6994) );
  MX4X1 U5265 ( .A(\registers[20][6] ), .B(\registers[21][6] ), .C(
        \registers[22][6] ), .D(\registers[23][6] ), .S0(n7596), .S1(n7826), 
        .Y(n7020) );
  MX4X1 U5266 ( .A(\registers[4][6] ), .B(\registers[5][6] ), .C(
        \registers[6][6] ), .D(\registers[7][6] ), .S0(n7596), .S1(n7827), .Y(
        n7025) );
  MX4X1 U5267 ( .A(\registers[52][6] ), .B(\registers[53][6] ), .C(
        \registers[54][6] ), .D(\registers[55][6] ), .S0(n7595), .S1(n7826), 
        .Y(n7010) );
  MX4X1 U5268 ( .A(\registers[36][6] ), .B(\registers[37][6] ), .C(
        \registers[38][6] ), .D(\registers[39][6] ), .S0(n7595), .S1(n7826), 
        .Y(n7015) );
  MX4X1 U5269 ( .A(\registers[212][6] ), .B(\registers[213][6] ), .C(
        \registers[214][6] ), .D(\registers[215][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6957) );
  MX4X1 U5270 ( .A(\registers[196][6] ), .B(\registers[197][6] ), .C(
        \registers[198][6] ), .D(\registers[199][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6962) );
  MX4X1 U5271 ( .A(\registers[244][6] ), .B(\registers[245][6] ), .C(
        \registers[246][6] ), .D(\registers[247][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6947) );
  MX4X1 U5272 ( .A(\registers[228][6] ), .B(\registers[229][6] ), .C(
        \registers[230][6] ), .D(\registers[231][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6952) );
  MX4X1 U5273 ( .A(\registers[148][6] ), .B(\registers[149][6] ), .C(
        \registers[150][6] ), .D(\registers[151][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6978) );
  MX4X1 U5274 ( .A(\registers[132][6] ), .B(\registers[133][6] ), .C(
        \registers[134][6] ), .D(\registers[135][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6983) );
  MX4X1 U5275 ( .A(\registers[180][6] ), .B(\registers[181][6] ), .C(
        \registers[182][6] ), .D(\registers[183][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6968) );
  MX4X1 U5276 ( .A(\registers[164][6] ), .B(\registers[165][6] ), .C(
        \registers[166][6] ), .D(\registers[167][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6973) );
  MX4X1 U5277 ( .A(\registers[852][6] ), .B(\registers[853][6] ), .C(
        \registers[854][6] ), .D(\registers[855][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6744) );
  MX4X1 U5278 ( .A(\registers[836][6] ), .B(\registers[837][6] ), .C(
        \registers[838][6] ), .D(\registers[839][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6749) );
  MX4X1 U5279 ( .A(\registers[884][6] ), .B(\registers[885][6] ), .C(
        \registers[886][6] ), .D(\registers[887][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6734) );
  MX4X1 U5280 ( .A(\registers[868][6] ), .B(\registers[869][6] ), .C(
        \registers[870][6] ), .D(\registers[871][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6739) );
  MX4X1 U5281 ( .A(\registers[788][6] ), .B(\registers[789][6] ), .C(
        \registers[790][6] ), .D(\registers[791][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6765) );
  MX4X1 U5282 ( .A(\registers[772][6] ), .B(\registers[773][6] ), .C(
        \registers[774][6] ), .D(\registers[775][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6770) );
  MX4X1 U5283 ( .A(\registers[820][6] ), .B(\registers[821][6] ), .C(
        \registers[822][6] ), .D(\registers[823][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6755) );
  MX4X1 U5284 ( .A(\registers[804][6] ), .B(\registers[805][6] ), .C(
        \registers[806][6] ), .D(\registers[807][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6760) );
  MX4X1 U5285 ( .A(\registers[980][6] ), .B(\registers[981][6] ), .C(
        \registers[982][6] ), .D(\registers[983][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6702) );
  MX4X1 U5286 ( .A(\registers[964][6] ), .B(\registers[965][6] ), .C(
        \registers[966][6] ), .D(\registers[967][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6707) );
  MX4X1 U5287 ( .A(\registers[1012][6] ), .B(\registers[1013][6] ), .C(
        \registers[1014][6] ), .D(\registers[1015][6] ), .S0(n7575), .S1(n7807), .Y(n6692) );
  MX4X1 U5288 ( .A(\registers[996][6] ), .B(\registers[997][6] ), .C(
        \registers[998][6] ), .D(\registers[999][6] ), .S0(n7575), .S1(n7808), 
        .Y(n6697) );
  MX4X1 U5289 ( .A(\registers[916][6] ), .B(\registers[917][6] ), .C(
        \registers[918][6] ), .D(\registers[919][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6723) );
  MX4X1 U5290 ( .A(\registers[900][6] ), .B(\registers[901][6] ), .C(
        \registers[902][6] ), .D(\registers[903][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6728) );
  MX4X1 U5291 ( .A(\registers[948][6] ), .B(\registers[949][6] ), .C(
        \registers[950][6] ), .D(\registers[951][6] ), .S0(n7576), .S1(n7809), 
        .Y(n6713) );
  MX4X1 U5292 ( .A(\registers[932][6] ), .B(\registers[933][6] ), .C(
        \registers[934][6] ), .D(\registers[935][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6718) );
  MX4X1 U5293 ( .A(\registers[596][6] ), .B(\registers[597][6] ), .C(
        \registers[598][6] ), .D(\registers[599][6] ), .S0(n7584), .S1(n7815), 
        .Y(n6829) );
  MX4X1 U5294 ( .A(\registers[580][6] ), .B(\registers[581][6] ), .C(
        \registers[582][6] ), .D(\registers[583][6] ), .S0(n7584), .S1(n7816), 
        .Y(n6834) );
  MX4X1 U5295 ( .A(\registers[628][6] ), .B(\registers[629][6] ), .C(
        \registers[630][6] ), .D(\registers[631][6] ), .S0(n7583), .S1(n7815), 
        .Y(n6819) );
  MX4X1 U5296 ( .A(\registers[612][6] ), .B(\registers[613][6] ), .C(
        \registers[614][6] ), .D(\registers[615][6] ), .S0(n7583), .S1(n7815), 
        .Y(n6824) );
  MX4X1 U5297 ( .A(\registers[532][6] ), .B(\registers[533][6] ), .C(
        \registers[534][6] ), .D(\registers[535][6] ), .S0(n7585), .S1(n7817), 
        .Y(n6850) );
  MX4X1 U5298 ( .A(\registers[516][6] ), .B(\registers[517][6] ), .C(
        \registers[518][6] ), .D(\registers[519][6] ), .S0(n7585), .S1(n7817), 
        .Y(n6855) );
  MX4X1 U5299 ( .A(\registers[564][6] ), .B(\registers[565][6] ), .C(
        \registers[566][6] ), .D(\registers[567][6] ), .S0(n7584), .S1(n7816), 
        .Y(n6840) );
  MX4X1 U5300 ( .A(\registers[548][6] ), .B(\registers[549][6] ), .C(
        \registers[550][6] ), .D(\registers[551][6] ), .S0(n7585), .S1(n7816), 
        .Y(n6845) );
  MX4X1 U5301 ( .A(\registers[724][6] ), .B(\registers[725][6] ), .C(
        \registers[726][6] ), .D(\registers[727][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6787) );
  MX4X1 U5302 ( .A(\registers[708][6] ), .B(\registers[709][6] ), .C(
        \registers[710][6] ), .D(\registers[711][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6792) );
  MX4X1 U5303 ( .A(\registers[756][6] ), .B(\registers[757][6] ), .C(
        \registers[758][6] ), .D(\registers[759][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6777) );
  MX4X1 U5304 ( .A(\registers[740][6] ), .B(\registers[741][6] ), .C(
        \registers[742][6] ), .D(\registers[743][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6782) );
  MX4X1 U5305 ( .A(\registers[660][6] ), .B(\registers[661][6] ), .C(
        \registers[662][6] ), .D(\registers[663][6] ), .S0(n7582), .S1(n7814), 
        .Y(n6808) );
  MX4X1 U5306 ( .A(\registers[644][6] ), .B(\registers[645][6] ), .C(
        \registers[646][6] ), .D(\registers[647][6] ), .S0(n7583), .S1(n7814), 
        .Y(n6813) );
  MX4X1 U5307 ( .A(\registers[692][6] ), .B(\registers[693][6] ), .C(
        \registers[694][6] ), .D(\registers[695][6] ), .S0(n7582), .S1(n7813), 
        .Y(n6798) );
  MX4X1 U5308 ( .A(\registers[676][6] ), .B(\registers[677][6] ), .C(
        \registers[678][6] ), .D(\registers[679][6] ), .S0(n7582), .S1(n7814), 
        .Y(n6803) );
  MX4X1 U5309 ( .A(\registers[340][7] ), .B(\registers[341][7] ), .C(
        \registers[342][7] ), .D(\registers[343][7] ), .S0(n7610), .S1(n7840), 
        .Y(n7254) );
  MX4X1 U5310 ( .A(\registers[324][7] ), .B(\registers[325][7] ), .C(
        \registers[326][7] ), .D(\registers[327][7] ), .S0(n7611), .S1(n7840), 
        .Y(n7259) );
  MX4X1 U5311 ( .A(\registers[372][7] ), .B(\registers[373][7] ), .C(
        \registers[374][7] ), .D(\registers[375][7] ), .S0(n7610), .S1(n7839), 
        .Y(n7244) );
  MX4X1 U5312 ( .A(\registers[356][7] ), .B(\registers[357][7] ), .C(
        \registers[358][7] ), .D(\registers[359][7] ), .S0(n7610), .S1(n7840), 
        .Y(n7249) );
  MX4X1 U5313 ( .A(\registers[468][7] ), .B(\registers[469][7] ), .C(
        \registers[470][7] ), .D(\registers[471][7] ), .S0(n7608), .S1(n7837), 
        .Y(n7212) );
  MX4X1 U5314 ( .A(\registers[452][7] ), .B(\registers[453][7] ), .C(
        \registers[454][7] ), .D(\registers[455][7] ), .S0(n7608), .S1(n7838), 
        .Y(n7217) );
  MX4X1 U5315 ( .A(\registers[500][7] ), .B(\registers[501][7] ), .C(
        \registers[502][7] ), .D(\registers[503][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7202) );
  MX4X1 U5316 ( .A(\registers[484][7] ), .B(\registers[485][7] ), .C(
        \registers[486][7] ), .D(\registers[487][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7207) );
  MX4X1 U5317 ( .A(\registers[404][7] ), .B(\registers[405][7] ), .C(
        \registers[406][7] ), .D(\registers[407][7] ), .S0(n7609), .S1(n7839), 
        .Y(n7233) );
  MX4X1 U5318 ( .A(\registers[388][7] ), .B(\registers[389][7] ), .C(
        \registers[390][7] ), .D(\registers[391][7] ), .S0(n7609), .S1(n7839), 
        .Y(n7238) );
  MX4X1 U5319 ( .A(\registers[436][7] ), .B(\registers[437][7] ), .C(
        \registers[438][7] ), .D(\registers[439][7] ), .S0(n7608), .S1(n7838), 
        .Y(n7223) );
  MX4X1 U5320 ( .A(\registers[420][7] ), .B(\registers[421][7] ), .C(
        \registers[422][7] ), .D(\registers[423][7] ), .S0(n7609), .S1(n7838), 
        .Y(n7228) );
  MX4X1 U5321 ( .A(\registers[276][7] ), .B(\registers[277][7] ), .C(
        \registers[278][7] ), .D(\registers[279][7] ), .S0(n7612), .S1(n7841), 
        .Y(n7275) );
  MX4X1 U5322 ( .A(\registers[260][7] ), .B(\registers[261][7] ), .C(
        \registers[262][7] ), .D(\registers[263][7] ), .S0(n7612), .S1(n7841), 
        .Y(n7280) );
  MX4X1 U5323 ( .A(\registers[308][7] ), .B(\registers[309][7] ), .C(
        \registers[310][7] ), .D(\registers[311][7] ), .S0(n7611), .S1(n7841), 
        .Y(n7265) );
  MX4X1 U5324 ( .A(\registers[292][7] ), .B(\registers[293][7] ), .C(
        \registers[294][7] ), .D(\registers[295][7] ), .S0(n7611), .S1(n7841), 
        .Y(n7270) );
  MX4X1 U5325 ( .A(\registers[212][7] ), .B(\registers[213][7] ), .C(
        \registers[214][7] ), .D(\registers[215][7] ), .S0(n7613), .S1(n7842), 
        .Y(n7297) );
  MX4X1 U5326 ( .A(\registers[196][7] ), .B(\registers[197][7] ), .C(
        \registers[198][7] ), .D(\registers[199][7] ), .S0(n7613), .S1(n7843), 
        .Y(n7302) );
  MX4X1 U5327 ( .A(\registers[244][7] ), .B(\registers[245][7] ), .C(
        \registers[246][7] ), .D(\registers[247][7] ), .S0(n7612), .S1(n7842), 
        .Y(n7287) );
  MX4X1 U5328 ( .A(\registers[228][7] ), .B(\registers[229][7] ), .C(
        \registers[230][7] ), .D(\registers[231][7] ), .S0(n7613), .S1(n7842), 
        .Y(n7292) );
  MX4X1 U5329 ( .A(\registers[84][7] ), .B(\registers[85][7] ), .C(
        \registers[86][7] ), .D(\registers[87][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7339) );
  MX4X1 U5330 ( .A(\registers[68][7] ), .B(\registers[69][7] ), .C(
        \registers[70][7] ), .D(\registers[71][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7344) );
  MX4X1 U5331 ( .A(\registers[116][7] ), .B(\registers[117][7] ), .C(
        \registers[118][7] ), .D(\registers[119][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7329) );
  MX4X1 U5332 ( .A(\registers[100][7] ), .B(\registers[101][7] ), .C(
        \registers[102][7] ), .D(\registers[103][7] ), .S0(n7615), .S1(n7845), 
        .Y(n7334) );
  MX4X1 U5333 ( .A(\registers[20][7] ), .B(\registers[21][7] ), .C(
        \registers[22][7] ), .D(\registers[23][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7360) );
  MX4X1 U5334 ( .A(\registers[4][7] ), .B(\registers[5][7] ), .C(
        \registers[6][7] ), .D(\registers[7][7] ), .S0(n7617), .S1(n7846), .Y(
        n7365) );
  MX4X1 U5335 ( .A(\registers[52][7] ), .B(\registers[53][7] ), .C(
        \registers[54][7] ), .D(\registers[55][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7350) );
  MX4X1 U5336 ( .A(\registers[36][7] ), .B(\registers[37][7] ), .C(
        \registers[38][7] ), .D(\registers[39][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7355) );
  MX4X1 U5337 ( .A(\registers[148][7] ), .B(\registers[149][7] ), .C(
        \registers[150][7] ), .D(\registers[151][7] ), .S0(n7614), .S1(n7844), 
        .Y(n7318) );
  MX4X1 U5338 ( .A(\registers[132][7] ), .B(\registers[133][7] ), .C(
        \registers[134][7] ), .D(\registers[135][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7323) );
  MX4X1 U5339 ( .A(\registers[180][7] ), .B(\registers[181][7] ), .C(
        \registers[182][7] ), .D(\registers[183][7] ), .S0(n7614), .S1(n7843), 
        .Y(n7308) );
  MX4X1 U5340 ( .A(\registers[164][7] ), .B(\registers[165][7] ), .C(
        \registers[166][7] ), .D(\registers[167][7] ), .S0(n7614), .S1(n7843), 
        .Y(n7313) );
  MX4X1 U5341 ( .A(\registers[852][7] ), .B(\registers[853][7] ), .C(
        \registers[854][7] ), .D(\registers[855][7] ), .S0(n7600), .S1(n7830), 
        .Y(n7084) );
  MX4X1 U5342 ( .A(\registers[836][7] ), .B(\registers[837][7] ), .C(
        \registers[838][7] ), .D(\registers[839][7] ), .S0(n7600), .S1(n7830), 
        .Y(n7089) );
  MX4X1 U5343 ( .A(\registers[884][7] ), .B(\registers[885][7] ), .C(
        \registers[886][7] ), .D(\registers[887][7] ), .S0(n7599), .S1(n7829), 
        .Y(n7074) );
  MX4X1 U5344 ( .A(\registers[868][7] ), .B(\registers[869][7] ), .C(
        \registers[870][7] ), .D(\registers[871][7] ), .S0(n7599), .S1(n7830), 
        .Y(n7079) );
  MX4X1 U5345 ( .A(\registers[788][7] ), .B(\registers[789][7] ), .C(
        \registers[790][7] ), .D(\registers[791][7] ), .S0(n7601), .S1(n7831), 
        .Y(n7105) );
  MX4X1 U5346 ( .A(\registers[772][7] ), .B(\registers[773][7] ), .C(
        \registers[774][7] ), .D(\registers[775][7] ), .S0(n7601), .S1(n7832), 
        .Y(n7110) );
  MX4X1 U5347 ( .A(\registers[820][7] ), .B(\registers[821][7] ), .C(
        \registers[822][7] ), .D(\registers[823][7] ), .S0(n7600), .S1(n7831), 
        .Y(n7095) );
  MX4X1 U5348 ( .A(\registers[804][7] ), .B(\registers[805][7] ), .C(
        \registers[806][7] ), .D(\registers[807][7] ), .S0(n7601), .S1(n7831), 
        .Y(n7100) );
  MX4X1 U5349 ( .A(\registers[980][7] ), .B(\registers[981][7] ), .C(
        \registers[982][7] ), .D(\registers[983][7] ), .S0(n7597), .S1(n7828), 
        .Y(n7042) );
  MX4X1 U5350 ( .A(\registers[964][7] ), .B(\registers[965][7] ), .C(
        \registers[966][7] ), .D(\registers[967][7] ), .S0(n7597), .S1(n7828), 
        .Y(n7047) );
  MX4X1 U5351 ( .A(\registers[1012][7] ), .B(\registers[1013][7] ), .C(
        \registers[1014][7] ), .D(\registers[1015][7] ), .S0(n7596), .S1(n7827), .Y(n7032) );
  MX4X1 U5352 ( .A(\registers[996][7] ), .B(\registers[997][7] ), .C(
        \registers[998][7] ), .D(\registers[999][7] ), .S0(n7597), .S1(n7827), 
        .Y(n7037) );
  MX4X1 U5353 ( .A(\registers[916][7] ), .B(\registers[917][7] ), .C(
        \registers[918][7] ), .D(\registers[919][7] ), .S0(n7598), .S1(n7829), 
        .Y(n7063) );
  MX4X1 U5354 ( .A(\registers[900][7] ), .B(\registers[901][7] ), .C(
        \registers[902][7] ), .D(\registers[903][7] ), .S0(n7599), .S1(n7829), 
        .Y(n7068) );
  MX4X1 U5355 ( .A(\registers[948][7] ), .B(\registers[949][7] ), .C(
        \registers[950][7] ), .D(\registers[951][7] ), .S0(n7598), .S1(n7828), 
        .Y(n7053) );
  MX4X1 U5356 ( .A(\registers[932][7] ), .B(\registers[933][7] ), .C(
        \registers[934][7] ), .D(\registers[935][7] ), .S0(n7598), .S1(n7829), 
        .Y(n7058) );
  MX4X1 U5357 ( .A(\registers[596][7] ), .B(\registers[597][7] ), .C(
        \registers[598][7] ), .D(\registers[599][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7169) );
  MX4X1 U5358 ( .A(\registers[580][7] ), .B(\registers[581][7] ), .C(
        \registers[582][7] ), .D(\registers[583][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7174) );
  MX4X1 U5359 ( .A(\registers[628][7] ), .B(\registers[629][7] ), .C(
        \registers[630][7] ), .D(\registers[631][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7159) );
  MX4X1 U5360 ( .A(\registers[612][7] ), .B(\registers[613][7] ), .C(
        \registers[614][7] ), .D(\registers[615][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7164) );
  MX4X1 U5361 ( .A(\registers[532][7] ), .B(\registers[533][7] ), .C(
        \registers[534][7] ), .D(\registers[535][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7190) );
  MX4X1 U5362 ( .A(\registers[516][7] ), .B(\registers[517][7] ), .C(
        \registers[518][7] ), .D(\registers[519][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7195) );
  MX4X1 U5363 ( .A(\registers[564][7] ), .B(\registers[565][7] ), .C(
        \registers[566][7] ), .D(\registers[567][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7180) );
  MX4X1 U5364 ( .A(\registers[548][7] ), .B(\registers[549][7] ), .C(
        \registers[550][7] ), .D(\registers[551][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7185) );
  MX4X1 U5365 ( .A(\registers[724][7] ), .B(\registers[725][7] ), .C(
        \registers[726][7] ), .D(\registers[727][7] ), .S0(n7602), .S1(n7833), 
        .Y(n7127) );
  MX4X1 U5366 ( .A(\registers[708][7] ), .B(\registers[709][7] ), .C(
        \registers[710][7] ), .D(\registers[711][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7132) );
  MX4X1 U5367 ( .A(\registers[756][7] ), .B(\registers[757][7] ), .C(
        \registers[758][7] ), .D(\registers[759][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7117) );
  MX4X1 U5368 ( .A(\registers[740][7] ), .B(\registers[741][7] ), .C(
        \registers[742][7] ), .D(\registers[743][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7122) );
  MX4X1 U5369 ( .A(\registers[660][7] ), .B(\registers[661][7] ), .C(
        \registers[662][7] ), .D(\registers[663][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7148) );
  MX4X1 U5370 ( .A(\registers[644][7] ), .B(\registers[645][7] ), .C(
        \registers[646][7] ), .D(\registers[647][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7153) );
  MX4X1 U5371 ( .A(\registers[692][7] ), .B(\registers[693][7] ), .C(
        \registers[694][7] ), .D(\registers[695][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7138) );
  MX4X1 U5372 ( .A(\registers[676][7] ), .B(\registers[677][7] ), .C(
        \registers[678][7] ), .D(\registers[679][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7143) );
  MX4X1 U5373 ( .A(n1426), .B(n1424), .C(n1425), .D(n1423), .S0(n4615), .S1(
        n4528), .Y(n1427) );
  MX4X1 U5374 ( .A(\registers[344][0] ), .B(\registers[345][0] ), .C(
        \registers[346][0] ), .D(\registers[347][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1424) );
  MX4X1 U5375 ( .A(\registers[348][0] ), .B(\registers[349][0] ), .C(
        \registers[350][0] ), .D(\registers[351][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1423) );
  MX4X1 U5376 ( .A(\registers[336][0] ), .B(\registers[337][0] ), .C(
        \registers[338][0] ), .D(\registers[339][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1426) );
  MX4X1 U5377 ( .A(n1449), .B(n1447), .C(n1448), .D(n1446), .S0(n4587), .S1(
        n4529), .Y(n1450) );
  MX4X1 U5378 ( .A(\registers[280][0] ), .B(\registers[281][0] ), .C(
        \registers[282][0] ), .D(\registers[283][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1447) );
  MX4X1 U5379 ( .A(\registers[284][0] ), .B(\registers[285][0] ), .C(
        \registers[286][0] ), .D(\registers[287][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1446) );
  MX4X1 U5380 ( .A(\registers[272][0] ), .B(\registers[273][0] ), .C(
        \registers[274][0] ), .D(\registers[275][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1449) );
  MX4X1 U5381 ( .A(n1382), .B(n1380), .C(n1381), .D(n1379), .S0(n4604), .S1(
        n4528), .Y(n1383) );
  MX4X1 U5382 ( .A(\registers[472][0] ), .B(\registers[473][0] ), .C(
        \registers[474][0] ), .D(\registers[475][0] ), .S0(n4115), .S1(n4357), 
        .Y(n1380) );
  MX4X1 U5383 ( .A(\registers[476][0] ), .B(\registers[477][0] ), .C(
        \registers[478][0] ), .D(\registers[479][0] ), .S0(n4115), .S1(n4356), 
        .Y(n1379) );
  MX4X1 U5384 ( .A(\registers[464][0] ), .B(\registers[465][0] ), .C(
        \registers[466][0] ), .D(\registers[467][0] ), .S0(n4115), .S1(n4357), 
        .Y(n1382) );
  MX4X1 U5385 ( .A(n1405), .B(n1402), .C(n1404), .D(n1400), .S0(n4607), .S1(
        n4528), .Y(n1406) );
  MX4X1 U5386 ( .A(\registers[408][0] ), .B(\registers[409][0] ), .C(
        \registers[410][0] ), .D(\registers[411][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1402) );
  MX4X1 U5387 ( .A(\registers[412][0] ), .B(\registers[413][0] ), .C(
        \registers[414][0] ), .D(\registers[415][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1400) );
  MX4X1 U5388 ( .A(\registers[400][0] ), .B(\registers[401][0] ), .C(
        \registers[402][0] ), .D(\registers[403][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1405) );
  MX4X1 U5389 ( .A(n1517), .B(n1515), .C(n1516), .D(n1514), .S0(n4588), .S1(
        n4530), .Y(n1518) );
  MX4X1 U5390 ( .A(\registers[88][0] ), .B(\registers[89][0] ), .C(
        \registers[90][0] ), .D(\registers[91][0] ), .S0(n4123), .S1(n4364), 
        .Y(n1515) );
  MX4X1 U5391 ( .A(\registers[92][0] ), .B(\registers[93][0] ), .C(
        \registers[94][0] ), .D(\registers[95][0] ), .S0(n4123), .S1(n4364), 
        .Y(n1514) );
  MX4X1 U5392 ( .A(\registers[80][0] ), .B(\registers[81][0] ), .C(
        \registers[82][0] ), .D(\registers[83][0] ), .S0(n4123), .S1(n4364), 
        .Y(n1517) );
  MX4X1 U5393 ( .A(n1540), .B(n1536), .C(n1538), .D(n1535), .S0(n4588), .S1(
        n4530), .Y(n1541) );
  MX4X1 U5394 ( .A(\registers[24][0] ), .B(\registers[25][0] ), .C(
        \registers[26][0] ), .D(\registers[27][0] ), .S0(n4125), .S1(n4365), 
        .Y(n1536) );
  MX4X1 U5395 ( .A(\registers[28][0] ), .B(\registers[29][0] ), .C(
        \registers[30][0] ), .D(\registers[31][0] ), .S0(n4125), .S1(n4365), 
        .Y(n1535) );
  MX4X1 U5396 ( .A(\registers[16][0] ), .B(\registers[17][0] ), .C(
        \registers[18][0] ), .D(\registers[19][0] ), .S0(n4125), .S1(n4365), 
        .Y(n1540) );
  MX4X1 U5397 ( .A(n1473), .B(n1470), .C(n1472), .D(n1468), .S0(n4587), .S1(
        n4529), .Y(n1474) );
  MX4X1 U5398 ( .A(\registers[216][0] ), .B(\registers[217][0] ), .C(
        \registers[218][0] ), .D(\registers[219][0] ), .S0(n4121), .S1(n4361), 
        .Y(n1470) );
  MX4X1 U5399 ( .A(\registers[220][0] ), .B(\registers[221][0] ), .C(
        \registers[222][0] ), .D(\registers[223][0] ), .S0(n4121), .S1(n4361), 
        .Y(n1468) );
  MX4X1 U5400 ( .A(\registers[208][0] ), .B(\registers[209][0] ), .C(
        \registers[210][0] ), .D(\registers[211][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1473) );
  MX4X1 U5401 ( .A(n1494), .B(n1492), .C(n1493), .D(n1491), .S0(n4587), .S1(
        n4529), .Y(n1495) );
  MX4X1 U5402 ( .A(\registers[152][0] ), .B(\registers[153][0] ), .C(
        \registers[154][0] ), .D(\registers[155][0] ), .S0(n4122), .S1(n4363), 
        .Y(n1492) );
  MX4X1 U5403 ( .A(\registers[156][0] ), .B(\registers[157][0] ), .C(
        \registers[158][0] ), .D(\registers[159][0] ), .S0(n4122), .S1(n4363), 
        .Y(n1491) );
  MX4X1 U5404 ( .A(\registers[144][0] ), .B(\registers[145][0] ), .C(
        \registers[146][0] ), .D(\registers[147][0] ), .S0(n4122), .S1(n4363), 
        .Y(n1494) );
  MX4X1 U5405 ( .A(n1100), .B(n1098), .C(n1099), .D(n1097), .S0(n4590), .S1(
        n4526), .Y(n1101) );
  MX4X1 U5406 ( .A(\registers[856][0] ), .B(\registers[857][0] ), .C(
        \registers[858][0] ), .D(\registers[859][0] ), .S0(n4107), .S1(n4474), 
        .Y(n1098) );
  MX4X1 U5407 ( .A(\registers[860][0] ), .B(\registers[861][0] ), .C(
        \registers[862][0] ), .D(\registers[863][0] ), .S0(n4107), .S1(n4454), 
        .Y(n1097) );
  MX4X1 U5408 ( .A(\registers[848][0] ), .B(\registers[849][0] ), .C(
        \registers[850][0] ), .D(\registers[851][0] ), .S0(n4107), .S1(n4476), 
        .Y(n1100) );
  MX4X1 U5409 ( .A(n1163), .B(n1161), .C(n1162), .D(n1160), .S0(n4591), .S1(
        n4526), .Y(n1164) );
  MX4X1 U5410 ( .A(\registers[792][0] ), .B(\registers[793][0] ), .C(
        \registers[794][0] ), .D(\registers[795][0] ), .S0(n4109), .S1(n4366), 
        .Y(n1161) );
  MX4X1 U5411 ( .A(\registers[796][0] ), .B(\registers[797][0] ), .C(
        \registers[798][0] ), .D(\registers[799][0] ), .S0(n4109), .S1(n4385), 
        .Y(n1160) );
  MX4X1 U5412 ( .A(\registers[784][0] ), .B(\registers[785][0] ), .C(
        \registers[786][0] ), .D(\registers[787][0] ), .S0(n4109), .S1(n4351), 
        .Y(n1163) );
  MX4X1 U5413 ( .A(n1336), .B(n1333), .C(n1335), .D(n1331), .S0(n4605), .S1(
        n4527), .Y(n1337) );
  MX4X1 U5414 ( .A(\registers[600][0] ), .B(\registers[601][0] ), .C(
        \registers[602][0] ), .D(\registers[603][0] ), .S0(n4113), .S1(n4354), 
        .Y(n1333) );
  MX4X1 U5415 ( .A(\registers[604][0] ), .B(\registers[605][0] ), .C(
        \registers[606][0] ), .D(\registers[607][0] ), .S0(n4113), .S1(n4354), 
        .Y(n1331) );
  MX4X1 U5416 ( .A(\registers[592][0] ), .B(\registers[593][0] ), .C(
        \registers[594][0] ), .D(\registers[595][0] ), .S0(n4113), .S1(n4354), 
        .Y(n1336) );
  MX4X1 U5417 ( .A(n1357), .B(n1355), .C(n1356), .D(n1354), .S0(n4606), .S1(
        n4527), .Y(n1358) );
  MX4X1 U5418 ( .A(\registers[536][0] ), .B(\registers[537][0] ), .C(
        \registers[538][0] ), .D(\registers[539][0] ), .S0(n4114), .S1(n4355), 
        .Y(n1355) );
  MX4X1 U5419 ( .A(\registers[540][0] ), .B(\registers[541][0] ), .C(
        \registers[542][0] ), .D(\registers[543][0] ), .S0(n4114), .S1(n4355), 
        .Y(n1354) );
  MX4X1 U5420 ( .A(\registers[528][0] ), .B(\registers[529][0] ), .C(
        \registers[530][0] ), .D(\registers[531][0] ), .S0(n4114), .S1(n4355), 
        .Y(n1357) );
  MX4X1 U5421 ( .A(n1195), .B(n1183), .C(n1184), .D(n1182), .S0(n4588), .S1(
        n4527), .Y(n1198) );
  MX4X1 U5422 ( .A(\registers[728][0] ), .B(\registers[729][0] ), .C(
        \registers[730][0] ), .D(\registers[731][0] ), .S0(n4110), .S1(n4352), 
        .Y(n1183) );
  MX4X1 U5423 ( .A(\registers[732][0] ), .B(\registers[733][0] ), .C(
        \registers[734][0] ), .D(\registers[735][0] ), .S0(n4110), .S1(n4352), 
        .Y(n1182) );
  MX4X1 U5424 ( .A(\registers[720][0] ), .B(\registers[721][0] ), .C(
        \registers[722][0] ), .D(\registers[723][0] ), .S0(n4110), .S1(n4352), 
        .Y(n1195) );
  MX4X1 U5425 ( .A(n1295), .B(n1291), .C(n1293), .D(n1289), .S0(n4611), .S1(
        n4527), .Y(n1297) );
  MX4X1 U5426 ( .A(\registers[664][0] ), .B(\registers[665][0] ), .C(
        \registers[666][0] ), .D(\registers[667][0] ), .S0(n4111), .S1(n4353), 
        .Y(n1291) );
  MX4X1 U5427 ( .A(\registers[668][0] ), .B(\registers[669][0] ), .C(
        \registers[670][0] ), .D(\registers[671][0] ), .S0(n4111), .S1(n4353), 
        .Y(n1289) );
  MX4X1 U5428 ( .A(\registers[656][0] ), .B(\registers[657][0] ), .C(
        \registers[658][0] ), .D(\registers[659][0] ), .S0(n4111), .S1(n4353), 
        .Y(n1295) );
  MX4X1 U5429 ( .A(n1784), .B(n1782), .C(n1783), .D(n1781), .S0(n4592), .S1(
        n4533), .Y(n1785) );
  MX4X1 U5430 ( .A(\registers[344][1] ), .B(\registers[345][1] ), .C(
        \registers[346][1] ), .D(\registers[347][1] ), .S0(n4139), .S1(n4379), 
        .Y(n1782) );
  MX4X1 U5431 ( .A(\registers[348][1] ), .B(\registers[349][1] ), .C(
        \registers[350][1] ), .D(\registers[351][1] ), .S0(n4139), .S1(n4379), 
        .Y(n1781) );
  MX4X1 U5432 ( .A(\registers[336][1] ), .B(\registers[337][1] ), .C(
        \registers[338][1] ), .D(\registers[339][1] ), .S0(n4139), .S1(n4379), 
        .Y(n1784) );
  MX4X1 U5433 ( .A(n1805), .B(n1803), .C(n1804), .D(n1802), .S0(n4592), .S1(
        n4534), .Y(n1807) );
  MX4X1 U5434 ( .A(\registers[280][1] ), .B(\registers[281][1] ), .C(
        \registers[282][1] ), .D(\registers[283][1] ), .S0(n4141), .S1(n4380), 
        .Y(n1803) );
  MX4X1 U5435 ( .A(\registers[284][1] ), .B(\registers[285][1] ), .C(
        \registers[286][1] ), .D(\registers[287][1] ), .S0(n4141), .S1(n4380), 
        .Y(n1802) );
  MX4X1 U5436 ( .A(\registers[272][1] ), .B(\registers[273][1] ), .C(
        \registers[274][1] ), .D(\registers[275][1] ), .S0(n4141), .S1(n4380), 
        .Y(n1805) );
  MX4X1 U5437 ( .A(n1741), .B(n1738), .C(n1739), .D(n1737), .S0(n4591), .S1(
        n4533), .Y(n1742) );
  MX4X1 U5438 ( .A(\registers[472][1] ), .B(\registers[473][1] ), .C(
        \registers[474][1] ), .D(\registers[475][1] ), .S0(n4137), .S1(n4376), 
        .Y(n1738) );
  MX4X1 U5439 ( .A(\registers[476][1] ), .B(\registers[477][1] ), .C(
        \registers[478][1] ), .D(\registers[479][1] ), .S0(n4137), .S1(n4376), 
        .Y(n1737) );
  MX4X1 U5440 ( .A(\registers[464][1] ), .B(\registers[465][1] ), .C(
        \registers[466][1] ), .D(\registers[467][1] ), .S0(n4137), .S1(n4376), 
        .Y(n1741) );
  MX4X1 U5441 ( .A(n1762), .B(n1760), .C(n1761), .D(n1759), .S0(n4591), .S1(
        n4533), .Y(n1763) );
  MX4X1 U5442 ( .A(\registers[408][1] ), .B(\registers[409][1] ), .C(
        \registers[410][1] ), .D(\registers[411][1] ), .S0(n4138), .S1(n4377), 
        .Y(n1760) );
  MX4X1 U5443 ( .A(\registers[412][1] ), .B(\registers[413][1] ), .C(
        \registers[414][1] ), .D(\registers[415][1] ), .S0(n4138), .S1(n4377), 
        .Y(n1759) );
  MX4X1 U5444 ( .A(\registers[400][1] ), .B(\registers[401][1] ), .C(
        \registers[402][1] ), .D(\registers[403][1] ), .S0(n4138), .S1(n4378), 
        .Y(n1762) );
  MX4X1 U5445 ( .A(n1872), .B(n1869), .C(n1870), .D(n1868), .S0(n4593), .S1(
        n4535), .Y(n1874) );
  MX4X1 U5446 ( .A(\registers[88][1] ), .B(\registers[89][1] ), .C(
        \registers[90][1] ), .D(\registers[91][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1869) );
  MX4X1 U5447 ( .A(\registers[92][1] ), .B(\registers[93][1] ), .C(
        \registers[94][1] ), .D(\registers[95][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1868) );
  MX4X1 U5448 ( .A(\registers[80][1] ), .B(\registers[81][1] ), .C(
        \registers[82][1] ), .D(\registers[83][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1872) );
  MX4X1 U5449 ( .A(n1894), .B(n1892), .C(n1893), .D(n1891), .S0(n4593), .S1(
        n4535), .Y(n1895) );
  MX4X1 U5450 ( .A(\registers[24][1] ), .B(\registers[25][1] ), .C(
        \registers[26][1] ), .D(\registers[27][1] ), .S0(n4146), .S1(n4385), 
        .Y(n1892) );
  MX4X1 U5451 ( .A(\registers[28][1] ), .B(\registers[29][1] ), .C(
        \registers[30][1] ), .D(\registers[31][1] ), .S0(n4146), .S1(n4385), 
        .Y(n1891) );
  MX4X1 U5452 ( .A(\registers[16][1] ), .B(\registers[17][1] ), .C(
        \registers[18][1] ), .D(\registers[19][1] ), .S0(n4146), .S1(n4385), 
        .Y(n1894) );
  MX4X1 U5453 ( .A(n1828), .B(n1826), .C(n1827), .D(n1825), .S0(n4592), .S1(
        n4534), .Y(n1829) );
  MX4X1 U5454 ( .A(\registers[216][1] ), .B(\registers[217][1] ), .C(
        \registers[218][1] ), .D(\registers[219][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1826) );
  MX4X1 U5455 ( .A(\registers[220][1] ), .B(\registers[221][1] ), .C(
        \registers[222][1] ), .D(\registers[223][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1825) );
  MX4X1 U5456 ( .A(\registers[208][1] ), .B(\registers[209][1] ), .C(
        \registers[210][1] ), .D(\registers[211][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1828) );
  MX4X1 U5457 ( .A(n1850), .B(n1848), .C(n1849), .D(n1847), .S0(n4593), .S1(
        n4534), .Y(n1851) );
  MX4X1 U5458 ( .A(\registers[152][1] ), .B(\registers[153][1] ), .C(
        \registers[154][1] ), .D(\registers[155][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1848) );
  MX4X1 U5459 ( .A(\registers[156][1] ), .B(\registers[157][1] ), .C(
        \registers[158][1] ), .D(\registers[159][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1847) );
  MX4X1 U5460 ( .A(\registers[144][1] ), .B(\registers[145][1] ), .C(
        \registers[146][1] ), .D(\registers[147][1] ), .S0(n4143), .S1(n4383), 
        .Y(n1850) );
  MX4X1 U5461 ( .A(n1609), .B(n1604), .C(n1607), .D(n1603), .S0(n4589), .S1(
        n4531), .Y(n1610) );
  MX4X1 U5462 ( .A(\registers[856][1] ), .B(\registers[857][1] ), .C(
        \registers[858][1] ), .D(\registers[859][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1604) );
  MX4X1 U5463 ( .A(\registers[860][1] ), .B(\registers[861][1] ), .C(
        \registers[862][1] ), .D(\registers[863][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1603) );
  MX4X1 U5464 ( .A(\registers[848][1] ), .B(\registers[849][1] ), .C(
        \registers[850][1] ), .D(\registers[851][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1609) );
  MX4X1 U5465 ( .A(n1630), .B(n1628), .C(n1629), .D(n1627), .S0(n4589), .S1(
        n4531), .Y(n1631) );
  MX4X1 U5466 ( .A(\registers[792][1] ), .B(\registers[793][1] ), .C(
        \registers[794][1] ), .D(\registers[795][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1628) );
  MX4X1 U5467 ( .A(\registers[796][1] ), .B(\registers[797][1] ), .C(
        \registers[798][1] ), .D(\registers[799][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1627) );
  MX4X1 U5468 ( .A(\registers[784][1] ), .B(\registers[785][1] ), .C(
        \registers[786][1] ), .D(\registers[787][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1630) );
  MX4X1 U5469 ( .A(n1562), .B(n1560), .C(n1561), .D(n1559), .S0(n4588), .S1(
        n4530), .Y(n1563) );
  MX4X1 U5470 ( .A(\registers[984][1] ), .B(\registers[985][1] ), .C(
        \registers[986][1] ), .D(\registers[987][1] ), .S0(n4126), .S1(n4366), 
        .Y(n1560) );
  MX4X1 U5471 ( .A(\registers[988][1] ), .B(\registers[989][1] ), .C(
        \registers[990][1] ), .D(\registers[991][1] ), .S0(n4126), .S1(n4366), 
        .Y(n1559) );
  MX4X1 U5472 ( .A(\registers[976][1] ), .B(\registers[977][1] ), .C(
        \registers[978][1] ), .D(\registers[979][1] ), .S0(n4126), .S1(n4367), 
        .Y(n1562) );
  MX4X1 U5473 ( .A(n1585), .B(n1583), .C(n1584), .D(n1582), .S0(n4589), .S1(
        n4531), .Y(n1586) );
  MX4X1 U5474 ( .A(\registers[920][1] ), .B(\registers[921][1] ), .C(
        \registers[922][1] ), .D(\registers[923][1] ), .S0(n4127), .S1(n4368), 
        .Y(n1583) );
  MX4X1 U5475 ( .A(\registers[924][1] ), .B(\registers[925][1] ), .C(
        \registers[926][1] ), .D(\registers[927][1] ), .S0(n4127), .S1(n4368), 
        .Y(n1582) );
  MX4X1 U5476 ( .A(\registers[912][1] ), .B(\registers[913][1] ), .C(
        \registers[914][1] ), .D(\registers[915][1] ), .S0(n4127), .S1(n4368), 
        .Y(n1585) );
  MX4X1 U5477 ( .A(n1696), .B(n1694), .C(n1695), .D(n1693), .S0(n4590), .S1(
        n4532), .Y(n1697) );
  MX4X1 U5478 ( .A(\registers[600][1] ), .B(\registers[601][1] ), .C(
        \registers[602][1] ), .D(\registers[603][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1694) );
  MX4X1 U5479 ( .A(\registers[604][1] ), .B(\registers[605][1] ), .C(
        \registers[606][1] ), .D(\registers[607][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1693) );
  MX4X1 U5480 ( .A(\registers[592][1] ), .B(\registers[593][1] ), .C(
        \registers[594][1] ), .D(\registers[595][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1696) );
  MX4X1 U5481 ( .A(n1718), .B(n1716), .C(n1717), .D(n1715), .S0(n4591), .S1(
        n4532), .Y(n1719) );
  MX4X1 U5482 ( .A(\registers[536][1] ), .B(\registers[537][1] ), .C(
        \registers[538][1] ), .D(\registers[539][1] ), .S0(n4135), .S1(n4375), 
        .Y(n1716) );
  MX4X1 U5483 ( .A(\registers[540][1] ), .B(\registers[541][1] ), .C(
        \registers[542][1] ), .D(\registers[543][1] ), .S0(n4135), .S1(n4375), 
        .Y(n1715) );
  MX4X1 U5484 ( .A(\registers[528][1] ), .B(\registers[529][1] ), .C(
        \registers[530][1] ), .D(\registers[531][1] ), .S0(n4135), .S1(n4375), 
        .Y(n1718) );
  MX4X1 U5485 ( .A(n1653), .B(n1651), .C(n1652), .D(n1650), .S0(n4590), .S1(
        n4531), .Y(n1654) );
  MX4X1 U5486 ( .A(\registers[728][1] ), .B(\registers[729][1] ), .C(
        \registers[730][1] ), .D(\registers[731][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1651) );
  MX4X1 U5487 ( .A(\registers[732][1] ), .B(\registers[733][1] ), .C(
        \registers[734][1] ), .D(\registers[735][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1650) );
  MX4X1 U5488 ( .A(\registers[720][1] ), .B(\registers[721][1] ), .C(
        \registers[722][1] ), .D(\registers[723][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1653) );
  MX4X1 U5489 ( .A(n1675), .B(n1672), .C(n1673), .D(n1671), .S0(n4590), .S1(
        n4532), .Y(n1676) );
  MX4X1 U5490 ( .A(\registers[664][1] ), .B(\registers[665][1] ), .C(
        \registers[666][1] ), .D(\registers[667][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1672) );
  MX4X1 U5491 ( .A(\registers[668][1] ), .B(\registers[669][1] ), .C(
        \registers[670][1] ), .D(\registers[671][1] ), .S0(n4133), .S1(n4372), 
        .Y(n1671) );
  MX4X1 U5492 ( .A(\registers[656][1] ), .B(\registers[657][1] ), .C(
        \registers[658][1] ), .D(\registers[659][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1675) );
  MX4X1 U5493 ( .A(n2135), .B(n2133), .C(n2134), .D(n2132), .S0(n4597), .S1(
        n4538), .Y(n2137) );
  MX4X1 U5494 ( .A(\registers[344][2] ), .B(\registers[345][2] ), .C(
        \registers[346][2] ), .D(\registers[347][2] ), .S0(n4161), .S1(n4398), 
        .Y(n2133) );
  MX4X1 U5495 ( .A(\registers[348][2] ), .B(\registers[349][2] ), .C(
        \registers[350][2] ), .D(\registers[351][2] ), .S0(n4161), .S1(n4398), 
        .Y(n2132) );
  MX4X1 U5496 ( .A(\registers[336][2] ), .B(\registers[337][2] ), .C(
        \registers[338][2] ), .D(\registers[339][2] ), .S0(n4161), .S1(n4399), 
        .Y(n2135) );
  MX4X1 U5497 ( .A(n2158), .B(n2156), .C(n2157), .D(n2155), .S0(n4597), .S1(
        n4539), .Y(n2159) );
  MX4X1 U5498 ( .A(\registers[280][2] ), .B(\registers[281][2] ), .C(
        \registers[282][2] ), .D(\registers[283][2] ), .S0(n4162), .S1(n4400), 
        .Y(n2156) );
  MX4X1 U5499 ( .A(\registers[284][2] ), .B(\registers[285][2] ), .C(
        \registers[286][2] ), .D(\registers[287][2] ), .S0(n4162), .S1(n4400), 
        .Y(n2155) );
  MX4X1 U5500 ( .A(\registers[272][2] ), .B(\registers[273][2] ), .C(
        \registers[274][2] ), .D(\registers[275][2] ), .S0(n4162), .S1(n4400), 
        .Y(n2158) );
  MX4X1 U5501 ( .A(n2092), .B(n2090), .C(n2091), .D(n2089), .S0(n4596), .S1(
        n4538), .Y(n2093) );
  MX4X1 U5502 ( .A(\registers[472][2] ), .B(\registers[473][2] ), .C(
        \registers[474][2] ), .D(\registers[475][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2090) );
  MX4X1 U5503 ( .A(\registers[476][2] ), .B(\registers[477][2] ), .C(
        \registers[478][2] ), .D(\registers[479][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2089) );
  MX4X1 U5504 ( .A(\registers[464][2] ), .B(\registers[465][2] ), .C(
        \registers[466][2] ), .D(\registers[467][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2092) );
  MX4X1 U5505 ( .A(n2114), .B(n2112), .C(n2113), .D(n2111), .S0(n4597), .S1(
        n4538), .Y(n2115) );
  MX4X1 U5506 ( .A(\registers[408][2] ), .B(\registers[409][2] ), .C(
        \registers[410][2] ), .D(\registers[411][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2112) );
  MX4X1 U5507 ( .A(\registers[412][2] ), .B(\registers[413][2] ), .C(
        \registers[414][2] ), .D(\registers[415][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2111) );
  MX4X1 U5508 ( .A(\registers[400][2] ), .B(\registers[401][2] ), .C(
        \registers[402][2] ), .D(\registers[403][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2114) );
  MX4X1 U5509 ( .A(n2224), .B(n2222), .C(n2223), .D(n2221), .S0(n4598), .S1(
        n4539), .Y(n2225) );
  MX4X1 U5510 ( .A(\registers[88][2] ), .B(\registers[89][2] ), .C(
        \registers[90][2] ), .D(\registers[91][2] ), .S0(n4166), .S1(n4403), 
        .Y(n2222) );
  MX4X1 U5511 ( .A(\registers[92][2] ), .B(\registers[93][2] ), .C(
        \registers[94][2] ), .D(\registers[95][2] ), .S0(n4166), .S1(n4403), 
        .Y(n2221) );
  MX4X1 U5512 ( .A(\registers[80][2] ), .B(\registers[81][2] ), .C(
        \registers[82][2] ), .D(\registers[83][2] ), .S0(n4166), .S1(n4403), 
        .Y(n2224) );
  MX4X1 U5513 ( .A(n2246), .B(n2244), .C(n2245), .D(n2243), .S0(n4599), .S1(
        n4540), .Y(n2247) );
  MX4X1 U5514 ( .A(\registers[24][2] ), .B(\registers[25][2] ), .C(
        \registers[26][2] ), .D(\registers[27][2] ), .S0(n4167), .S1(n4405), 
        .Y(n2244) );
  MX4X1 U5515 ( .A(\registers[28][2] ), .B(\registers[29][2] ), .C(
        \registers[30][2] ), .D(\registers[31][2] ), .S0(n4167), .S1(n4404), 
        .Y(n2243) );
  MX4X1 U5516 ( .A(\registers[16][2] ), .B(\registers[17][2] ), .C(
        \registers[18][2] ), .D(\registers[19][2] ), .S0(n4167), .S1(n4405), 
        .Y(n2246) );
  MX4X1 U5517 ( .A(n2181), .B(n2179), .C(n2180), .D(n2178), .S0(n4598), .S1(
        n4539), .Y(n2182) );
  MX4X1 U5518 ( .A(\registers[216][2] ), .B(\registers[217][2] ), .C(
        \registers[218][2] ), .D(\registers[219][2] ), .S0(n4163), .S1(n4401), 
        .Y(n2179) );
  MX4X1 U5519 ( .A(\registers[220][2] ), .B(\registers[221][2] ), .C(
        \registers[222][2] ), .D(\registers[223][2] ), .S0(n4163), .S1(n4401), 
        .Y(n2178) );
  MX4X1 U5520 ( .A(\registers[208][2] ), .B(\registers[209][2] ), .C(
        \registers[210][2] ), .D(\registers[211][2] ), .S0(n4163), .S1(n4401), 
        .Y(n2181) );
  MX4X1 U5521 ( .A(n2202), .B(n2200), .C(n2201), .D(n2199), .S0(n4598), .S1(
        n4539), .Y(n2203) );
  MX4X1 U5522 ( .A(\registers[152][2] ), .B(\registers[153][2] ), .C(
        \registers[154][2] ), .D(\registers[155][2] ), .S0(n4165), .S1(n4402), 
        .Y(n2200) );
  MX4X1 U5523 ( .A(\registers[156][2] ), .B(\registers[157][2] ), .C(
        \registers[158][2] ), .D(\registers[159][2] ), .S0(n4165), .S1(n4402), 
        .Y(n2199) );
  MX4X1 U5524 ( .A(\registers[144][2] ), .B(\registers[145][2] ), .C(
        \registers[146][2] ), .D(\registers[147][2] ), .S0(n4165), .S1(n4402), 
        .Y(n2202) );
  MX4X1 U5525 ( .A(n1960), .B(n1958), .C(n1959), .D(n1957), .S0(n4594), .S1(
        n4536), .Y(n1961) );
  MX4X1 U5526 ( .A(\registers[856][2] ), .B(\registers[857][2] ), .C(
        \registers[858][2] ), .D(\registers[859][2] ), .S0(n4150), .S1(n4389), 
        .Y(n1958) );
  MX4X1 U5527 ( .A(\registers[860][2] ), .B(\registers[861][2] ), .C(
        \registers[862][2] ), .D(\registers[863][2] ), .S0(n4150), .S1(n4388), 
        .Y(n1957) );
  MX4X1 U5528 ( .A(\registers[848][2] ), .B(\registers[849][2] ), .C(
        \registers[850][2] ), .D(\registers[851][2] ), .S0(n4150), .S1(n4389), 
        .Y(n1960) );
  MX4X1 U5529 ( .A(n1982), .B(n1980), .C(n1981), .D(n1979), .S0(n4595), .S1(
        n4536), .Y(n1983) );
  MX4X1 U5530 ( .A(\registers[792][2] ), .B(\registers[793][2] ), .C(
        \registers[794][2] ), .D(\registers[795][2] ), .S0(n4151), .S1(n4390), 
        .Y(n1980) );
  MX4X1 U5531 ( .A(\registers[796][2] ), .B(\registers[797][2] ), .C(
        \registers[798][2] ), .D(\registers[799][2] ), .S0(n4151), .S1(n4390), 
        .Y(n1979) );
  MX4X1 U5532 ( .A(\registers[784][2] ), .B(\registers[785][2] ), .C(
        \registers[786][2] ), .D(\registers[787][2] ), .S0(n4151), .S1(n4390), 
        .Y(n1982) );
  MX4X1 U5533 ( .A(n1917), .B(n1915), .C(n1916), .D(n1914), .S0(n4594), .S1(
        n4535), .Y(n1918) );
  MX4X1 U5534 ( .A(\registers[984][2] ), .B(\registers[985][2] ), .C(
        \registers[986][2] ), .D(\registers[987][2] ), .S0(n4147), .S1(n4386), 
        .Y(n1915) );
  MX4X1 U5535 ( .A(\registers[988][2] ), .B(\registers[989][2] ), .C(
        \registers[990][2] ), .D(\registers[991][2] ), .S0(n4147), .S1(n4386), 
        .Y(n1914) );
  MX4X1 U5536 ( .A(\registers[976][2] ), .B(\registers[977][2] ), .C(
        \registers[978][2] ), .D(\registers[979][2] ), .S0(n4147), .S1(n4386), 
        .Y(n1917) );
  MX4X1 U5537 ( .A(n1938), .B(n1936), .C(n1937), .D(n1935), .S0(n4594), .S1(
        n4535), .Y(n1940) );
  MX4X1 U5538 ( .A(\registers[920][2] ), .B(\registers[921][2] ), .C(
        \registers[922][2] ), .D(\registers[923][2] ), .S0(n4149), .S1(n4387), 
        .Y(n1936) );
  MX4X1 U5539 ( .A(\registers[924][2] ), .B(\registers[925][2] ), .C(
        \registers[926][2] ), .D(\registers[927][2] ), .S0(n4149), .S1(n4387), 
        .Y(n1935) );
  MX4X1 U5540 ( .A(\registers[912][2] ), .B(\registers[913][2] ), .C(
        \registers[914][2] ), .D(\registers[915][2] ), .S0(n4149), .S1(n4387), 
        .Y(n1938) );
  MX4X1 U5541 ( .A(n2048), .B(n2046), .C(n2047), .D(n2045), .S0(n4596), .S1(
        n4537), .Y(n2049) );
  MX4X1 U5542 ( .A(\registers[600][2] ), .B(\registers[601][2] ), .C(
        \registers[602][2] ), .D(\registers[603][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2046) );
  MX4X1 U5543 ( .A(\registers[604][2] ), .B(\registers[605][2] ), .C(
        \registers[606][2] ), .D(\registers[607][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2045) );
  MX4X1 U5544 ( .A(\registers[592][2] ), .B(\registers[593][2] ), .C(
        \registers[594][2] ), .D(\registers[595][2] ), .S0(n4155), .S1(n4394), 
        .Y(n2048) );
  MX4X1 U5545 ( .A(n2069), .B(n2067), .C(n2068), .D(n2066), .S0(n4596), .S1(
        n4537), .Y(n2070) );
  MX4X1 U5546 ( .A(\registers[536][2] ), .B(\registers[537][2] ), .C(
        \registers[538][2] ), .D(\registers[539][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2067) );
  MX4X1 U5547 ( .A(\registers[540][2] ), .B(\registers[541][2] ), .C(
        \registers[542][2] ), .D(\registers[543][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2066) );
  MX4X1 U5548 ( .A(\registers[528][2] ), .B(\registers[529][2] ), .C(
        \registers[530][2] ), .D(\registers[531][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2069) );
  MX4X1 U5549 ( .A(n2004), .B(n2002), .C(n2003), .D(n2001), .S0(n4595), .S1(
        n4536), .Y(n2006) );
  MX4X1 U5550 ( .A(\registers[728][2] ), .B(\registers[729][2] ), .C(
        \registers[730][2] ), .D(\registers[731][2] ), .S0(n4153), .S1(n4391), 
        .Y(n2002) );
  MX4X1 U5551 ( .A(\registers[732][2] ), .B(\registers[733][2] ), .C(
        \registers[734][2] ), .D(\registers[735][2] ), .S0(n4153), .S1(n4391), 
        .Y(n2001) );
  MX4X1 U5552 ( .A(\registers[720][2] ), .B(\registers[721][2] ), .C(
        \registers[722][2] ), .D(\registers[723][2] ), .S0(n4153), .S1(n4391), 
        .Y(n2004) );
  MX4X1 U5553 ( .A(n2026), .B(n2024), .C(n2025), .D(n2023), .S0(n4595), .S1(
        n4537), .Y(n2027) );
  MX4X1 U5554 ( .A(\registers[664][2] ), .B(\registers[665][2] ), .C(
        \registers[666][2] ), .D(\registers[667][2] ), .S0(n4154), .S1(n4392), 
        .Y(n2024) );
  MX4X1 U5555 ( .A(\registers[668][2] ), .B(\registers[669][2] ), .C(
        \registers[670][2] ), .D(\registers[671][2] ), .S0(n4154), .S1(n4392), 
        .Y(n2023) );
  MX4X1 U5556 ( .A(\registers[656][2] ), .B(\registers[657][2] ), .C(
        \registers[658][2] ), .D(\registers[659][2] ), .S0(n4154), .S1(n4392), 
        .Y(n2026) );
  MX4X1 U5557 ( .A(n2550), .B(n2548), .C(n2549), .D(n2547), .S0(n4602), .S1(
        n4543), .Y(n2551) );
  MX4X1 U5558 ( .A(\registers[344][3] ), .B(\registers[345][3] ), .C(
        \registers[346][3] ), .D(\registers[347][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2548) );
  MX4X1 U5559 ( .A(\registers[348][3] ), .B(\registers[349][3] ), .C(
        \registers[350][3] ), .D(\registers[351][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2547) );
  MX4X1 U5560 ( .A(\registers[336][3] ), .B(\registers[337][3] ), .C(
        \registers[338][3] ), .D(\registers[339][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2550) );
  MX4X1 U5561 ( .A(n2571), .B(n2569), .C(n2570), .D(n2568), .S0(n4603), .S1(
        n4543), .Y(n2572) );
  MX4X1 U5562 ( .A(\registers[280][3] ), .B(\registers[281][3] ), .C(
        \registers[282][3] ), .D(\registers[283][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2569) );
  MX4X1 U5563 ( .A(\registers[284][3] ), .B(\registers[285][3] ), .C(
        \registers[286][3] ), .D(\registers[287][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2568) );
  MX4X1 U5564 ( .A(\registers[272][3] ), .B(\registers[273][3] ), .C(
        \registers[274][3] ), .D(\registers[275][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2571) );
  MX4X1 U5565 ( .A(n2508), .B(n2506), .C(n2507), .D(n2505), .S0(n4602), .S1(
        n4543), .Y(n2509) );
  MX4X1 U5566 ( .A(\registers[472][3] ), .B(\registers[473][3] ), .C(
        \registers[474][3] ), .D(\registers[475][3] ), .S0(n4179), .S1(n4416), 
        .Y(n2506) );
  MX4X1 U5567 ( .A(\registers[476][3] ), .B(\registers[477][3] ), .C(
        \registers[478][3] ), .D(\registers[479][3] ), .S0(n4179), .S1(n4416), 
        .Y(n2505) );
  MX4X1 U5568 ( .A(\registers[464][3] ), .B(\registers[465][3] ), .C(
        \registers[466][3] ), .D(\registers[467][3] ), .S0(n4179), .S1(n4416), 
        .Y(n2508) );
  MX4X1 U5569 ( .A(n2529), .B(n2527), .C(n2528), .D(n2526), .S0(n4602), .S1(
        n4543), .Y(n2530) );
  MX4X1 U5570 ( .A(\registers[408][3] ), .B(\registers[409][3] ), .C(
        \registers[410][3] ), .D(\registers[411][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2527) );
  MX4X1 U5571 ( .A(\registers[412][3] ), .B(\registers[413][3] ), .C(
        \registers[414][3] ), .D(\registers[415][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2526) );
  MX4X1 U5572 ( .A(\registers[400][3] ), .B(\registers[401][3] ), .C(
        \registers[402][3] ), .D(\registers[403][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2529) );
  MX4X1 U5573 ( .A(n2635), .B(n2633), .C(n2634), .D(n2632), .S0(n4604), .S1(
        n4539), .Y(n2636) );
  MX4X1 U5574 ( .A(\registers[88][3] ), .B(\registers[89][3] ), .C(
        \registers[90][3] ), .D(\registers[91][3] ), .S0(n4187), .S1(n4423), 
        .Y(n2633) );
  MX4X1 U5575 ( .A(\registers[92][3] ), .B(\registers[93][3] ), .C(
        \registers[94][3] ), .D(\registers[95][3] ), .S0(n4187), .S1(n4423), 
        .Y(n2632) );
  MX4X1 U5576 ( .A(\registers[80][3] ), .B(\registers[81][3] ), .C(
        \registers[82][3] ), .D(\registers[83][3] ), .S0(n4187), .S1(n4423), 
        .Y(n2635) );
  MX4X1 U5577 ( .A(n2656), .B(n2654), .C(n2655), .D(n2653), .S0(n4604), .S1(
        n4544), .Y(n2657) );
  MX4X1 U5578 ( .A(\registers[24][3] ), .B(\registers[25][3] ), .C(
        \registers[26][3] ), .D(\registers[27][3] ), .S0(n4189), .S1(n4424), 
        .Y(n2654) );
  MX4X1 U5579 ( .A(\registers[28][3] ), .B(\registers[29][3] ), .C(
        \registers[30][3] ), .D(\registers[31][3] ), .S0(n4189), .S1(n4424), 
        .Y(n2653) );
  MX4X1 U5580 ( .A(\registers[16][3] ), .B(\registers[17][3] ), .C(
        \registers[18][3] ), .D(\registers[19][3] ), .S0(n4189), .S1(n4424), 
        .Y(n2656) );
  MX4X1 U5581 ( .A(n2593), .B(n2591), .C(n2592), .D(n2590), .S0(n4603), .S1(
        n4535), .Y(n2594) );
  MX4X1 U5582 ( .A(\registers[216][3] ), .B(\registers[217][3] ), .C(
        \registers[218][3] ), .D(\registers[219][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2591) );
  MX4X1 U5583 ( .A(\registers[220][3] ), .B(\registers[221][3] ), .C(
        \registers[222][3] ), .D(\registers[223][3] ), .S0(n4185), .S1(n4420), 
        .Y(n2590) );
  MX4X1 U5584 ( .A(\registers[208][3] ), .B(\registers[209][3] ), .C(
        \registers[210][3] ), .D(\registers[211][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2593) );
  MX4X1 U5585 ( .A(n2614), .B(n2612), .C(n2613), .D(n2611), .S0(n4603), .S1(
        n4541), .Y(n2615) );
  MX4X1 U5586 ( .A(\registers[152][3] ), .B(\registers[153][3] ), .C(
        \registers[154][3] ), .D(\registers[155][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2612) );
  MX4X1 U5587 ( .A(\registers[156][3] ), .B(\registers[157][3] ), .C(
        \registers[158][3] ), .D(\registers[159][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2611) );
  MX4X1 U5588 ( .A(\registers[144][3] ), .B(\registers[145][3] ), .C(
        \registers[146][3] ), .D(\registers[147][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2614) );
  MX4X1 U5589 ( .A(n2312), .B(n2310), .C(n2311), .D(n2309), .S0(n4600), .S1(
        n4541), .Y(n2313) );
  MX4X1 U5590 ( .A(\registers[856][3] ), .B(\registers[857][3] ), .C(
        \registers[858][3] ), .D(\registers[859][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2310) );
  MX4X1 U5591 ( .A(\registers[860][3] ), .B(\registers[861][3] ), .C(
        \registers[862][3] ), .D(\registers[863][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2309) );
  MX4X1 U5592 ( .A(\registers[848][3] ), .B(\registers[849][3] ), .C(
        \registers[850][3] ), .D(\registers[851][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2312) );
  MX4X1 U5593 ( .A(n2333), .B(n2331), .C(n2332), .D(n2330), .S0(n4600), .S1(
        n4541), .Y(n2334) );
  MX4X1 U5594 ( .A(\registers[792][3] ), .B(\registers[793][3] ), .C(
        \registers[794][3] ), .D(\registers[795][3] ), .S0(n4173), .S1(n4409), 
        .Y(n2331) );
  MX4X1 U5595 ( .A(\registers[796][3] ), .B(\registers[797][3] ), .C(
        \registers[798][3] ), .D(\registers[799][3] ), .S0(n4173), .S1(n4409), 
        .Y(n2330) );
  MX4X1 U5596 ( .A(\registers[784][3] ), .B(\registers[785][3] ), .C(
        \registers[786][3] ), .D(\registers[787][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2333) );
  MX4X1 U5597 ( .A(n2268), .B(n2266), .C(n2267), .D(n2265), .S0(n4599), .S1(
        n4540), .Y(n2269) );
  MX4X1 U5598 ( .A(\registers[984][3] ), .B(\registers[985][3] ), .C(
        \registers[986][3] ), .D(\registers[987][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2266) );
  MX4X1 U5599 ( .A(\registers[988][3] ), .B(\registers[989][3] ), .C(
        \registers[990][3] ), .D(\registers[991][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2265) );
  MX4X1 U5600 ( .A(\registers[976][3] ), .B(\registers[977][3] ), .C(
        \registers[978][3] ), .D(\registers[979][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2268) );
  MX4X1 U5601 ( .A(n2290), .B(n2288), .C(n2289), .D(n2287), .S0(n4599), .S1(
        n4540), .Y(n2291) );
  MX4X1 U5602 ( .A(\registers[920][3] ), .B(\registers[921][3] ), .C(
        \registers[922][3] ), .D(\registers[923][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2288) );
  MX4X1 U5603 ( .A(\registers[924][3] ), .B(\registers[925][3] ), .C(
        \registers[926][3] ), .D(\registers[927][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2287) );
  MX4X1 U5604 ( .A(\registers[912][3] ), .B(\registers[913][3] ), .C(
        \registers[914][3] ), .D(\registers[915][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2290) );
  MX4X1 U5605 ( .A(n2465), .B(n2463), .C(n2464), .D(n2462), .S0(n4601), .S1(
        n4542), .Y(n2466) );
  MX4X1 U5606 ( .A(\registers[600][3] ), .B(\registers[601][3] ), .C(
        \registers[602][3] ), .D(\registers[603][3] ), .S0(n4177), .S1(n4413), 
        .Y(n2463) );
  MX4X1 U5607 ( .A(\registers[604][3] ), .B(\registers[605][3] ), .C(
        \registers[606][3] ), .D(\registers[607][3] ), .S0(n4177), .S1(n4413), 
        .Y(n2462) );
  MX4X1 U5608 ( .A(\registers[592][3] ), .B(\registers[593][3] ), .C(
        \registers[594][3] ), .D(\registers[595][3] ), .S0(n4177), .S1(n4413), 
        .Y(n2465) );
  MX4X1 U5609 ( .A(n2486), .B(n2484), .C(n2485), .D(n2483), .S0(n4601), .S1(
        n4542), .Y(n2487) );
  MX4X1 U5610 ( .A(\registers[536][3] ), .B(\registers[537][3] ), .C(
        \registers[538][3] ), .D(\registers[539][3] ), .S0(n4178), .S1(n4414), 
        .Y(n2484) );
  MX4X1 U5611 ( .A(\registers[540][3] ), .B(\registers[541][3] ), .C(
        \registers[542][3] ), .D(\registers[543][3] ), .S0(n4178), .S1(n4414), 
        .Y(n2483) );
  MX4X1 U5612 ( .A(\registers[528][3] ), .B(\registers[529][3] ), .C(
        \registers[530][3] ), .D(\registers[531][3] ), .S0(n4178), .S1(n4415), 
        .Y(n2486) );
  MX4X1 U5613 ( .A(n2367), .B(n2365), .C(n2366), .D(n2364), .S0(n4600), .S1(
        n4541), .Y(n2368) );
  MX4X1 U5614 ( .A(\registers[728][3] ), .B(\registers[729][3] ), .C(
        \registers[730][3] ), .D(\registers[731][3] ), .S0(n4174), .S1(n4411), 
        .Y(n2365) );
  MX4X1 U5615 ( .A(\registers[732][3] ), .B(\registers[733][3] ), .C(
        \registers[734][3] ), .D(\registers[735][3] ), .S0(n4174), .S1(n4411), 
        .Y(n2364) );
  MX4X1 U5616 ( .A(\registers[720][3] ), .B(\registers[721][3] ), .C(
        \registers[722][3] ), .D(\registers[723][3] ), .S0(n4174), .S1(n4411), 
        .Y(n2367) );
  MX4X1 U5617 ( .A(n2444), .B(n2442), .C(n2443), .D(n2441), .S0(n4601), .S1(
        n4542), .Y(n2445) );
  MX4X1 U5618 ( .A(\registers[664][3] ), .B(\registers[665][3] ), .C(
        \registers[666][3] ), .D(\registers[667][3] ), .S0(n4175), .S1(n4412), 
        .Y(n2442) );
  MX4X1 U5619 ( .A(\registers[668][3] ), .B(\registers[669][3] ), .C(
        \registers[670][3] ), .D(\registers[671][3] ), .S0(n4175), .S1(n4412), 
        .Y(n2441) );
  MX4X1 U5620 ( .A(\registers[656][3] ), .B(\registers[657][3] ), .C(
        \registers[658][3] ), .D(\registers[659][3] ), .S0(n4175), .S1(n4412), 
        .Y(n2444) );
  MX4X1 U5621 ( .A(n2890), .B(n2888), .C(n2889), .D(n2887), .S0(n4608), .S1(
        n4547), .Y(n2891) );
  MX4X1 U5622 ( .A(\registers[344][4] ), .B(\registers[345][4] ), .C(
        \registers[346][4] ), .D(\registers[347][4] ), .S0(n4203), .S1(n4438), 
        .Y(n2888) );
  MX4X1 U5623 ( .A(\registers[348][4] ), .B(\registers[349][4] ), .C(
        \registers[350][4] ), .D(\registers[351][4] ), .S0(n4203), .S1(n4438), 
        .Y(n2887) );
  MX4X1 U5624 ( .A(\registers[336][4] ), .B(\registers[337][4] ), .C(
        \registers[338][4] ), .D(\registers[339][4] ), .S0(n4203), .S1(n4438), 
        .Y(n2890) );
  MX4X1 U5625 ( .A(n2911), .B(n2909), .C(n2910), .D(n2908), .S0(n4608), .S1(
        n4547), .Y(n2912) );
  MX4X1 U5626 ( .A(\registers[280][4] ), .B(\registers[281][4] ), .C(
        \registers[282][4] ), .D(\registers[283][4] ), .S0(n4205), .S1(n4439), 
        .Y(n2909) );
  MX4X1 U5627 ( .A(\registers[284][4] ), .B(\registers[285][4] ), .C(
        \registers[286][4] ), .D(\registers[287][4] ), .S0(n4205), .S1(n4439), 
        .Y(n2908) );
  MX4X1 U5628 ( .A(\registers[272][4] ), .B(\registers[273][4] ), .C(
        \registers[274][4] ), .D(\registers[275][4] ), .S0(n4205), .S1(n4439), 
        .Y(n2911) );
  MX4X1 U5629 ( .A(n2848), .B(n2846), .C(n2847), .D(n2845), .S0(n4607), .S1(
        n4546), .Y(n2849) );
  MX4X1 U5630 ( .A(\registers[472][4] ), .B(\registers[473][4] ), .C(
        \registers[474][4] ), .D(\registers[475][4] ), .S0(n4201), .S1(n4435), 
        .Y(n2846) );
  MX4X1 U5631 ( .A(\registers[476][4] ), .B(\registers[477][4] ), .C(
        \registers[478][4] ), .D(\registers[479][4] ), .S0(n4201), .S1(n4435), 
        .Y(n2845) );
  MX4X1 U5632 ( .A(\registers[464][4] ), .B(\registers[465][4] ), .C(
        \registers[466][4] ), .D(\registers[467][4] ), .S0(n4201), .S1(n4435), 
        .Y(n2848) );
  MX4X1 U5633 ( .A(n2869), .B(n2867), .C(n2868), .D(n2866), .S0(n4607), .S1(
        n4547), .Y(n2870) );
  MX4X1 U5634 ( .A(\registers[408][4] ), .B(\registers[409][4] ), .C(
        \registers[410][4] ), .D(\registers[411][4] ), .S0(n4202), .S1(n4437), 
        .Y(n2867) );
  MX4X1 U5635 ( .A(\registers[412][4] ), .B(\registers[413][4] ), .C(
        \registers[414][4] ), .D(\registers[415][4] ), .S0(n4202), .S1(n4436), 
        .Y(n2866) );
  MX4X1 U5636 ( .A(\registers[400][4] ), .B(\registers[401][4] ), .C(
        \registers[402][4] ), .D(\registers[403][4] ), .S0(n4202), .S1(n4437), 
        .Y(n2869) );
  MX4X1 U5637 ( .A(n2975), .B(n2973), .C(n2974), .D(n2972), .S0(n4609), .S1(
        n4548), .Y(n2976) );
  MX4X1 U5638 ( .A(\registers[88][4] ), .B(\registers[89][4] ), .C(
        \registers[90][4] ), .D(\registers[91][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2973) );
  MX4X1 U5639 ( .A(\registers[92][4] ), .B(\registers[93][4] ), .C(
        \registers[94][4] ), .D(\registers[95][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2972) );
  MX4X1 U5640 ( .A(\registers[80][4] ), .B(\registers[81][4] ), .C(
        \registers[82][4] ), .D(\registers[83][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2975) );
  MX4X1 U5641 ( .A(n2996), .B(n2994), .C(n2995), .D(n2993), .S0(n4609), .S1(
        n4549), .Y(n2997) );
  MX4X1 U5642 ( .A(\registers[24][4] ), .B(\registers[25][4] ), .C(
        \registers[26][4] ), .D(\registers[27][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2994) );
  MX4X1 U5643 ( .A(\registers[28][4] ), .B(\registers[29][4] ), .C(
        \registers[30][4] ), .D(\registers[31][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2993) );
  MX4X1 U5644 ( .A(\registers[16][4] ), .B(\registers[17][4] ), .C(
        \registers[18][4] ), .D(\registers[19][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2996) );
  MX4X1 U5645 ( .A(n2933), .B(n2931), .C(n2932), .D(n2930), .S0(n4608), .S1(
        n4548), .Y(n2934) );
  MX4X1 U5646 ( .A(\registers[216][4] ), .B(\registers[217][4] ), .C(
        \registers[218][4] ), .D(\registers[219][4] ), .S0(n4206), .S1(n4440), 
        .Y(n2931) );
  MX4X1 U5647 ( .A(\registers[220][4] ), .B(\registers[221][4] ), .C(
        \registers[222][4] ), .D(\registers[223][4] ), .S0(n4206), .S1(n4440), 
        .Y(n2930) );
  MX4X1 U5648 ( .A(\registers[208][4] ), .B(\registers[209][4] ), .C(
        \registers[210][4] ), .D(\registers[211][4] ), .S0(n4206), .S1(n4440), 
        .Y(n2933) );
  MX4X1 U5649 ( .A(n2954), .B(n2952), .C(n2953), .D(n2951), .S0(n4609), .S1(
        n4548), .Y(n2955) );
  MX4X1 U5650 ( .A(\registers[152][4] ), .B(\registers[153][4] ), .C(
        \registers[154][4] ), .D(\registers[155][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2952) );
  MX4X1 U5651 ( .A(\registers[156][4] ), .B(\registers[157][4] ), .C(
        \registers[158][4] ), .D(\registers[159][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2951) );
  MX4X1 U5652 ( .A(\registers[144][4] ), .B(\registers[145][4] ), .C(
        \registers[146][4] ), .D(\registers[147][4] ), .S0(n4207), .S1(n4442), 
        .Y(n2954) );
  MX4X1 U5653 ( .A(n2720), .B(n2718), .C(n2719), .D(n2717), .S0(n4605), .S1(
        n4545), .Y(n2721) );
  MX4X1 U5654 ( .A(\registers[856][4] ), .B(\registers[857][4] ), .C(
        \registers[858][4] ), .D(\registers[859][4] ), .S0(n4193), .S1(n4428), 
        .Y(n2718) );
  MX4X1 U5655 ( .A(\registers[860][4] ), .B(\registers[861][4] ), .C(
        \registers[862][4] ), .D(\registers[863][4] ), .S0(n4193), .S1(n4428), 
        .Y(n2717) );
  MX4X1 U5656 ( .A(\registers[848][4] ), .B(\registers[849][4] ), .C(
        \registers[850][4] ), .D(\registers[851][4] ), .S0(n4193), .S1(n4428), 
        .Y(n2720) );
  MX4X1 U5657 ( .A(n2741), .B(n2739), .C(n2740), .D(n2738), .S0(n4605), .S1(
        n4545), .Y(n2742) );
  MX4X1 U5658 ( .A(\registers[792][4] ), .B(\registers[793][4] ), .C(
        \registers[794][4] ), .D(\registers[795][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2739) );
  MX4X1 U5659 ( .A(\registers[796][4] ), .B(\registers[797][4] ), .C(
        \registers[798][4] ), .D(\registers[799][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2738) );
  MX4X1 U5660 ( .A(\registers[784][4] ), .B(\registers[785][4] ), .C(
        \registers[786][4] ), .D(\registers[787][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2741) );
  MX4X1 U5661 ( .A(n2678), .B(n2676), .C(n2677), .D(n2675), .S0(n4604), .S1(
        n4544), .Y(n2679) );
  MX4X1 U5662 ( .A(\registers[984][4] ), .B(\registers[985][4] ), .C(
        \registers[986][4] ), .D(\registers[987][4] ), .S0(n4190), .S1(n4425), 
        .Y(n2676) );
  MX4X1 U5663 ( .A(\registers[988][4] ), .B(\registers[989][4] ), .C(
        \registers[990][4] ), .D(\registers[991][4] ), .S0(n4190), .S1(n4425), 
        .Y(n2675) );
  MX4X1 U5664 ( .A(\registers[976][4] ), .B(\registers[977][4] ), .C(
        \registers[978][4] ), .D(\registers[979][4] ), .S0(n4190), .S1(n4426), 
        .Y(n2678) );
  MX4X1 U5665 ( .A(n2699), .B(n2697), .C(n2698), .D(n2696), .S0(n4605), .S1(
        n4544), .Y(n2700) );
  MX4X1 U5666 ( .A(\registers[920][4] ), .B(\registers[921][4] ), .C(
        \registers[922][4] ), .D(\registers[923][4] ), .S0(n4191), .S1(n4427), 
        .Y(n2697) );
  MX4X1 U5667 ( .A(\registers[924][4] ), .B(\registers[925][4] ), .C(
        \registers[926][4] ), .D(\registers[927][4] ), .S0(n4191), .S1(n4427), 
        .Y(n2696) );
  MX4X1 U5668 ( .A(\registers[912][4] ), .B(\registers[913][4] ), .C(
        \registers[914][4] ), .D(\registers[915][4] ), .S0(n4191), .S1(n4427), 
        .Y(n2699) );
  MX4X1 U5669 ( .A(n2805), .B(n2803), .C(n2804), .D(n2802), .S0(n4606), .S1(
        n4546), .Y(n2806) );
  MX4X1 U5670 ( .A(\registers[600][4] ), .B(\registers[601][4] ), .C(
        \registers[602][4] ), .D(\registers[603][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2803) );
  MX4X1 U5671 ( .A(\registers[604][4] ), .B(\registers[605][4] ), .C(
        \registers[606][4] ), .D(\registers[607][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2802) );
  MX4X1 U5672 ( .A(\registers[592][4] ), .B(\registers[593][4] ), .C(
        \registers[594][4] ), .D(\registers[595][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2805) );
  MX4X1 U5673 ( .A(n2826), .B(n2824), .C(n2825), .D(n2823), .S0(n4607), .S1(
        n4546), .Y(n2827) );
  MX4X1 U5674 ( .A(\registers[536][4] ), .B(\registers[537][4] ), .C(
        \registers[538][4] ), .D(\registers[539][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2824) );
  MX4X1 U5675 ( .A(\registers[540][4] ), .B(\registers[541][4] ), .C(
        \registers[542][4] ), .D(\registers[543][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2823) );
  MX4X1 U5676 ( .A(\registers[528][4] ), .B(\registers[529][4] ), .C(
        \registers[530][4] ), .D(\registers[531][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2826) );
  MX4X1 U5677 ( .A(n2763), .B(n2761), .C(n2762), .D(n2760), .S0(n4606), .S1(
        n4545), .Y(n2764) );
  MX4X1 U5678 ( .A(\registers[728][4] ), .B(\registers[729][4] ), .C(
        \registers[730][4] ), .D(\registers[731][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2761) );
  MX4X1 U5679 ( .A(\registers[732][4] ), .B(\registers[733][4] ), .C(
        \registers[734][4] ), .D(\registers[735][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2760) );
  MX4X1 U5680 ( .A(\registers[720][4] ), .B(\registers[721][4] ), .C(
        \registers[722][4] ), .D(\registers[723][4] ), .S0(n4195), .S1(n4431), 
        .Y(n2763) );
  MX4X1 U5681 ( .A(n2784), .B(n2782), .C(n2783), .D(n2781), .S0(n4606), .S1(
        n4546), .Y(n2785) );
  MX4X1 U5682 ( .A(\registers[664][4] ), .B(\registers[665][4] ), .C(
        \registers[666][4] ), .D(\registers[667][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2782) );
  MX4X1 U5683 ( .A(\registers[668][4] ), .B(\registers[669][4] ), .C(
        \registers[670][4] ), .D(\registers[671][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2781) );
  MX4X1 U5684 ( .A(\registers[656][4] ), .B(\registers[657][4] ), .C(
        \registers[658][4] ), .D(\registers[659][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2784) );
  MX4X1 U5685 ( .A(n3230), .B(n3228), .C(n3229), .D(n3227), .S0(n4613), .S1(
        n4552), .Y(n3231) );
  MX4X1 U5686 ( .A(\registers[344][5] ), .B(\registers[345][5] ), .C(
        \registers[346][5] ), .D(\registers[347][5] ), .S0(n4225), .S1(n4457), 
        .Y(n3228) );
  MX4X1 U5687 ( .A(\registers[348][5] ), .B(\registers[349][5] ), .C(
        \registers[350][5] ), .D(\registers[351][5] ), .S0(n4225), .S1(n4457), 
        .Y(n3227) );
  MX4X1 U5688 ( .A(\registers[336][5] ), .B(\registers[337][5] ), .C(
        \registers[338][5] ), .D(\registers[339][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3230) );
  MX4X1 U5689 ( .A(n3251), .B(n3249), .C(n3250), .D(n3248), .S0(n4613), .S1(
        n4552), .Y(n3252) );
  MX4X1 U5690 ( .A(\registers[280][5] ), .B(\registers[281][5] ), .C(
        \registers[282][5] ), .D(\registers[283][5] ), .S0(n4226), .S1(n4459), 
        .Y(n3249) );
  MX4X1 U5691 ( .A(\registers[284][5] ), .B(\registers[285][5] ), .C(
        \registers[286][5] ), .D(\registers[287][5] ), .S0(n4226), .S1(n4459), 
        .Y(n3248) );
  MX4X1 U5692 ( .A(\registers[272][5] ), .B(\registers[273][5] ), .C(
        \registers[274][5] ), .D(\registers[275][5] ), .S0(n4226), .S1(n4459), 
        .Y(n3251) );
  MX4X1 U5693 ( .A(n3188), .B(n3186), .C(n3187), .D(n3185), .S0(n4612), .S1(
        n4551), .Y(n3189) );
  MX4X1 U5694 ( .A(\registers[472][5] ), .B(\registers[473][5] ), .C(
        \registers[474][5] ), .D(\registers[475][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3186) );
  MX4X1 U5695 ( .A(\registers[476][5] ), .B(\registers[477][5] ), .C(
        \registers[478][5] ), .D(\registers[479][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3185) );
  MX4X1 U5696 ( .A(\registers[464][5] ), .B(\registers[465][5] ), .C(
        \registers[466][5] ), .D(\registers[467][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3188) );
  MX4X1 U5697 ( .A(n3209), .B(n3207), .C(n3208), .D(n3206), .S0(n4613), .S1(
        n4552), .Y(n3210) );
  MX4X1 U5698 ( .A(\registers[408][5] ), .B(\registers[409][5] ), .C(
        \registers[410][5] ), .D(\registers[411][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3207) );
  MX4X1 U5699 ( .A(\registers[412][5] ), .B(\registers[413][5] ), .C(
        \registers[414][5] ), .D(\registers[415][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3206) );
  MX4X1 U5700 ( .A(\registers[400][5] ), .B(\registers[401][5] ), .C(
        \registers[402][5] ), .D(\registers[403][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3209) );
  MX4X1 U5701 ( .A(n3315), .B(n3313), .C(n3314), .D(n3312), .S0(n4614), .S1(
        n4553), .Y(n3316) );
  MX4X1 U5702 ( .A(\registers[88][5] ), .B(\registers[89][5] ), .C(
        \registers[90][5] ), .D(\registers[91][5] ), .S0(n4230), .S1(n4462), 
        .Y(n3313) );
  MX4X1 U5703 ( .A(\registers[92][5] ), .B(\registers[93][5] ), .C(
        \registers[94][5] ), .D(\registers[95][5] ), .S0(n4230), .S1(n4462), 
        .Y(n3312) );
  MX4X1 U5704 ( .A(\registers[80][5] ), .B(\registers[81][5] ), .C(
        \registers[82][5] ), .D(\registers[83][5] ), .S0(n4230), .S1(n4463), 
        .Y(n3315) );
  MX4X1 U5705 ( .A(n3336), .B(n3334), .C(n3335), .D(n3333), .S0(n4615), .S1(
        n4554), .Y(n3337) );
  MX4X1 U5706 ( .A(\registers[24][5] ), .B(\registers[25][5] ), .C(
        \registers[26][5] ), .D(\registers[27][5] ), .S0(n4231), .S1(n4464), 
        .Y(n3334) );
  MX4X1 U5707 ( .A(\registers[28][5] ), .B(\registers[29][5] ), .C(
        \registers[30][5] ), .D(\registers[31][5] ), .S0(n4231), .S1(n4464), 
        .Y(n3333) );
  MX4X1 U5708 ( .A(\registers[16][5] ), .B(\registers[17][5] ), .C(
        \registers[18][5] ), .D(\registers[19][5] ), .S0(n4231), .S1(n4464), 
        .Y(n3336) );
  MX4X1 U5709 ( .A(n3273), .B(n3271), .C(n3272), .D(n3270), .S0(n4614), .S1(
        n4553), .Y(n3274) );
  MX4X1 U5710 ( .A(\registers[216][5] ), .B(\registers[217][5] ), .C(
        \registers[218][5] ), .D(\registers[219][5] ), .S0(n4227), .S1(n4460), 
        .Y(n3271) );
  MX4X1 U5711 ( .A(\registers[220][5] ), .B(\registers[221][5] ), .C(
        \registers[222][5] ), .D(\registers[223][5] ), .S0(n4227), .S1(n4460), 
        .Y(n3270) );
  MX4X1 U5712 ( .A(\registers[208][5] ), .B(\registers[209][5] ), .C(
        \registers[210][5] ), .D(\registers[211][5] ), .S0(n4227), .S1(n4460), 
        .Y(n3273) );
  MX4X1 U5713 ( .A(n3294), .B(n3292), .C(n3293), .D(n3291), .S0(n4614), .S1(
        n4553), .Y(n3295) );
  MX4X1 U5714 ( .A(\registers[152][5] ), .B(\registers[153][5] ), .C(
        \registers[154][5] ), .D(\registers[155][5] ), .S0(n4229), .S1(n4461), 
        .Y(n3292) );
  MX4X1 U5715 ( .A(\registers[156][5] ), .B(\registers[157][5] ), .C(
        \registers[158][5] ), .D(\registers[159][5] ), .S0(n4229), .S1(n4461), 
        .Y(n3291) );
  MX4X1 U5716 ( .A(\registers[144][5] ), .B(\registers[145][5] ), .C(
        \registers[146][5] ), .D(\registers[147][5] ), .S0(n4229), .S1(n4461), 
        .Y(n3294) );
  MX4X1 U5717 ( .A(n3060), .B(n3058), .C(n3059), .D(n3057), .S0(n4610), .S1(
        n4550), .Y(n3061) );
  MX4X1 U5718 ( .A(\registers[856][5] ), .B(\registers[857][5] ), .C(
        \registers[858][5] ), .D(\registers[859][5] ), .S0(n4214), .S1(n4448), 
        .Y(n3058) );
  MX4X1 U5719 ( .A(\registers[860][5] ), .B(\registers[861][5] ), .C(
        \registers[862][5] ), .D(\registers[863][5] ), .S0(n4214), .S1(n4448), 
        .Y(n3057) );
  MX4X1 U5720 ( .A(\registers[848][5] ), .B(\registers[849][5] ), .C(
        \registers[850][5] ), .D(\registers[851][5] ), .S0(n4214), .S1(n4448), 
        .Y(n3060) );
  MX4X1 U5721 ( .A(n3081), .B(n3079), .C(n3080), .D(n3078), .S0(n4611), .S1(
        n4550), .Y(n3082) );
  MX4X1 U5722 ( .A(\registers[792][5] ), .B(\registers[793][5] ), .C(
        \registers[794][5] ), .D(\registers[795][5] ), .S0(n4215), .S1(n4449), 
        .Y(n3079) );
  MX4X1 U5723 ( .A(\registers[796][5] ), .B(\registers[797][5] ), .C(
        \registers[798][5] ), .D(\registers[799][5] ), .S0(n4215), .S1(n4449), 
        .Y(n3078) );
  MX4X1 U5724 ( .A(\registers[784][5] ), .B(\registers[785][5] ), .C(
        \registers[786][5] ), .D(\registers[787][5] ), .S0(n4215), .S1(n4449), 
        .Y(n3081) );
  MX4X1 U5725 ( .A(n3018), .B(n3016), .C(n3017), .D(n3015), .S0(n4610), .S1(
        n4549), .Y(n3019) );
  MX4X1 U5726 ( .A(\registers[984][5] ), .B(\registers[985][5] ), .C(
        \registers[986][5] ), .D(\registers[987][5] ), .S0(n4211), .S1(n4445), 
        .Y(n3016) );
  MX4X1 U5727 ( .A(\registers[988][5] ), .B(\registers[989][5] ), .C(
        \registers[990][5] ), .D(\registers[991][5] ), .S0(n4211), .S1(n4445), 
        .Y(n3015) );
  MX4X1 U5728 ( .A(\registers[976][5] ), .B(\registers[977][5] ), .C(
        \registers[978][5] ), .D(\registers[979][5] ), .S0(n4211), .S1(n4445), 
        .Y(n3018) );
  MX4X1 U5729 ( .A(n3039), .B(n3037), .C(n3038), .D(n3036), .S0(n4610), .S1(
        n4549), .Y(n3040) );
  MX4X1 U5730 ( .A(\registers[920][5] ), .B(\registers[921][5] ), .C(
        \registers[922][5] ), .D(\registers[923][5] ), .S0(n4213), .S1(n4446), 
        .Y(n3037) );
  MX4X1 U5731 ( .A(\registers[924][5] ), .B(\registers[925][5] ), .C(
        \registers[926][5] ), .D(\registers[927][5] ), .S0(n4213), .S1(n4446), 
        .Y(n3036) );
  MX4X1 U5732 ( .A(\registers[912][5] ), .B(\registers[913][5] ), .C(
        \registers[914][5] ), .D(\registers[915][5] ), .S0(n4213), .S1(n4447), 
        .Y(n3039) );
  MX4X1 U5733 ( .A(n3145), .B(n3143), .C(n3144), .D(n3142), .S0(n4612), .S1(
        n4551), .Y(n3146) );
  MX4X1 U5734 ( .A(\registers[600][5] ), .B(\registers[601][5] ), .C(
        \registers[602][5] ), .D(\registers[603][5] ), .S0(n4219), .S1(n4453), 
        .Y(n3143) );
  MX4X1 U5735 ( .A(\registers[604][5] ), .B(\registers[605][5] ), .C(
        \registers[606][5] ), .D(\registers[607][5] ), .S0(n4219), .S1(n4452), 
        .Y(n3142) );
  MX4X1 U5736 ( .A(\registers[592][5] ), .B(\registers[593][5] ), .C(
        \registers[594][5] ), .D(\registers[595][5] ), .S0(n4219), .S1(n4453), 
        .Y(n3145) );
  MX4X1 U5737 ( .A(n3166), .B(n3164), .C(n3165), .D(n3163), .S0(n4612), .S1(
        n4551), .Y(n3167) );
  MX4X1 U5738 ( .A(\registers[536][5] ), .B(\registers[537][5] ), .C(
        \registers[538][5] ), .D(\registers[539][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3164) );
  MX4X1 U5739 ( .A(\registers[540][5] ), .B(\registers[541][5] ), .C(
        \registers[542][5] ), .D(\registers[543][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3163) );
  MX4X1 U5740 ( .A(\registers[528][5] ), .B(\registers[529][5] ), .C(
        \registers[530][5] ), .D(\registers[531][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3166) );
  MX4X1 U5741 ( .A(n3103), .B(n3101), .C(n3102), .D(n3100), .S0(n4611), .S1(
        n4550), .Y(n3104) );
  MX4X1 U5742 ( .A(\registers[728][5] ), .B(\registers[729][5] ), .C(
        \registers[730][5] ), .D(\registers[731][5] ), .S0(n4217), .S1(n4450), 
        .Y(n3101) );
  MX4X1 U5743 ( .A(\registers[732][5] ), .B(\registers[733][5] ), .C(
        \registers[734][5] ), .D(\registers[735][5] ), .S0(n4217), .S1(n4450), 
        .Y(n3100) );
  MX4X1 U5744 ( .A(\registers[720][5] ), .B(\registers[721][5] ), .C(
        \registers[722][5] ), .D(\registers[723][5] ), .S0(n4217), .S1(n4450), 
        .Y(n3103) );
  MX4X1 U5745 ( .A(n3124), .B(n3122), .C(n3123), .D(n3121), .S0(n4611), .S1(
        n4550), .Y(n3125) );
  MX4X1 U5746 ( .A(\registers[664][5] ), .B(\registers[665][5] ), .C(
        \registers[666][5] ), .D(\registers[667][5] ), .S0(n4218), .S1(n4451), 
        .Y(n3122) );
  MX4X1 U5747 ( .A(\registers[668][5] ), .B(\registers[669][5] ), .C(
        \registers[670][5] ), .D(\registers[671][5] ), .S0(n4218), .S1(n4451), 
        .Y(n3121) );
  MX4X1 U5748 ( .A(\registers[656][5] ), .B(\registers[657][5] ), .C(
        \registers[658][5] ), .D(\registers[659][5] ), .S0(n4218), .S1(n4451), 
        .Y(n3124) );
  MX4X1 U5749 ( .A(n3570), .B(n3568), .C(n3569), .D(n3567), .S0(n4618), .S1(
        n4557), .Y(n3571) );
  MX4X1 U5750 ( .A(\registers[344][6] ), .B(\registers[345][6] ), .C(
        \registers[346][6] ), .D(\registers[347][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3568) );
  MX4X1 U5751 ( .A(\registers[348][6] ), .B(\registers[349][6] ), .C(
        \registers[350][6] ), .D(\registers[351][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3567) );
  MX4X1 U5752 ( .A(\registers[336][6] ), .B(\registers[337][6] ), .C(
        \registers[338][6] ), .D(\registers[339][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3570) );
  MX4X1 U5753 ( .A(n3591), .B(n3589), .C(n3590), .D(n3588), .S0(n4619), .S1(
        n4557), .Y(n3592) );
  MX4X1 U5754 ( .A(\registers[280][6] ), .B(\registers[281][6] ), .C(
        \registers[282][6] ), .D(\registers[283][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3589) );
  MX4X1 U5755 ( .A(\registers[284][6] ), .B(\registers[285][6] ), .C(
        \registers[286][6] ), .D(\registers[287][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3588) );
  MX4X1 U5756 ( .A(\registers[272][6] ), .B(\registers[273][6] ), .C(
        \registers[274][6] ), .D(\registers[275][6] ), .S0(n4247), .S1(n4479), 
        .Y(n3591) );
  MX4X1 U5757 ( .A(n3528), .B(n3526), .C(n3527), .D(n3525), .S0(n4618), .S1(
        n4556), .Y(n3529) );
  MX4X1 U5758 ( .A(\registers[472][6] ), .B(\registers[473][6] ), .C(
        \registers[474][6] ), .D(\registers[475][6] ), .S0(n4243), .S1(n4475), 
        .Y(n3526) );
  MX4X1 U5759 ( .A(\registers[476][6] ), .B(\registers[477][6] ), .C(
        \registers[478][6] ), .D(\registers[479][6] ), .S0(n4243), .S1(n4475), 
        .Y(n3525) );
  MX4X1 U5760 ( .A(\registers[464][6] ), .B(\registers[465][6] ), .C(
        \registers[466][6] ), .D(\registers[467][6] ), .S0(n4243), .S1(n4475), 
        .Y(n3528) );
  MX4X1 U5761 ( .A(n3549), .B(n3547), .C(n3548), .D(n3546), .S0(n4618), .S1(
        n4557), .Y(n3550) );
  MX4X1 U5762 ( .A(\registers[408][6] ), .B(\registers[409][6] ), .C(
        \registers[410][6] ), .D(\registers[411][6] ), .S0(n4245), .S1(n4476), 
        .Y(n3547) );
  MX4X1 U5763 ( .A(\registers[412][6] ), .B(\registers[413][6] ), .C(
        \registers[414][6] ), .D(\registers[415][6] ), .S0(n4245), .S1(n4476), 
        .Y(n3546) );
  MX4X1 U5764 ( .A(\registers[400][6] ), .B(\registers[401][6] ), .C(
        \registers[402][6] ), .D(\registers[403][6] ), .S0(n4245), .S1(n4476), 
        .Y(n3549) );
  MX4X1 U5765 ( .A(n3655), .B(n3653), .C(n3654), .D(n3652), .S0(n4620), .S1(
        n4532), .Y(n3656) );
  MX4X1 U5766 ( .A(\registers[88][6] ), .B(\registers[89][6] ), .C(
        \registers[90][6] ), .D(\registers[91][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3653) );
  MX4X1 U5767 ( .A(\registers[92][6] ), .B(\registers[93][6] ), .C(
        \registers[94][6] ), .D(\registers[95][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3652) );
  MX4X1 U5768 ( .A(\registers[80][6] ), .B(\registers[81][6] ), .C(
        \registers[82][6] ), .D(\registers[83][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3655) );
  MX4X1 U5769 ( .A(n3676), .B(n3674), .C(n3675), .D(n3673), .S0(n4620), .S1(
        N70), .Y(n3677) );
  MX4X1 U5770 ( .A(\registers[24][6] ), .B(\registers[25][6] ), .C(
        \registers[26][6] ), .D(\registers[27][6] ), .S0(n4253), .S1(n4483), 
        .Y(n3674) );
  MX4X1 U5771 ( .A(\registers[28][6] ), .B(\registers[29][6] ), .C(
        \registers[30][6] ), .D(\registers[31][6] ), .S0(n4253), .S1(n4483), 
        .Y(n3673) );
  MX4X1 U5772 ( .A(\registers[16][6] ), .B(\registers[17][6] ), .C(
        \registers[18][6] ), .D(\registers[19][6] ), .S0(n4253), .S1(n4483), 
        .Y(n3676) );
  MX4X1 U5773 ( .A(n3613), .B(n3611), .C(n3612), .D(n3610), .S0(n4619), .S1(
        n4527), .Y(n3614) );
  MX4X1 U5774 ( .A(\registers[216][6] ), .B(\registers[217][6] ), .C(
        \registers[218][6] ), .D(\registers[219][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3611) );
  MX4X1 U5775 ( .A(\registers[220][6] ), .B(\registers[221][6] ), .C(
        \registers[222][6] ), .D(\registers[223][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3610) );
  MX4X1 U5776 ( .A(\registers[208][6] ), .B(\registers[209][6] ), .C(
        \registers[210][6] ), .D(\registers[211][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3613) );
  MX4X1 U5777 ( .A(n3634), .B(n3632), .C(n3633), .D(n3631), .S0(n4619), .S1(
        N70), .Y(n3635) );
  MX4X1 U5778 ( .A(\registers[152][6] ), .B(\registers[153][6] ), .C(
        \registers[154][6] ), .D(\registers[155][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3632) );
  MX4X1 U5779 ( .A(\registers[156][6] ), .B(\registers[157][6] ), .C(
        \registers[158][6] ), .D(\registers[159][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3631) );
  MX4X1 U5780 ( .A(\registers[144][6] ), .B(\registers[145][6] ), .C(
        \registers[146][6] ), .D(\registers[147][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3634) );
  MX4X1 U5781 ( .A(n3400), .B(n3398), .C(n3399), .D(n3397), .S0(n4616), .S1(
        n4554), .Y(n3401) );
  MX4X1 U5782 ( .A(\registers[856][6] ), .B(\registers[857][6] ), .C(
        \registers[858][6] ), .D(\registers[859][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3398) );
  MX4X1 U5783 ( .A(\registers[860][6] ), .B(\registers[861][6] ), .C(
        \registers[862][6] ), .D(\registers[863][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3397) );
  MX4X1 U5784 ( .A(\registers[848][6] ), .B(\registers[849][6] ), .C(
        \registers[850][6] ), .D(\registers[851][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3400) );
  MX4X1 U5785 ( .A(n3421), .B(n3419), .C(n3420), .D(n3418), .S0(n4616), .S1(
        n4555), .Y(n3422) );
  MX4X1 U5786 ( .A(\registers[792][6] ), .B(\registers[793][6] ), .C(
        \registers[794][6] ), .D(\registers[795][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3419) );
  MX4X1 U5787 ( .A(\registers[796][6] ), .B(\registers[797][6] ), .C(
        \registers[798][6] ), .D(\registers[799][6] ), .S0(n4237), .S1(n4468), 
        .Y(n3418) );
  MX4X1 U5788 ( .A(\registers[784][6] ), .B(\registers[785][6] ), .C(
        \registers[786][6] ), .D(\registers[787][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3421) );
  MX4X1 U5789 ( .A(n3358), .B(n3356), .C(n3357), .D(n3355), .S0(n4615), .S1(
        n4554), .Y(n3359) );
  MX4X1 U5790 ( .A(\registers[984][6] ), .B(\registers[985][6] ), .C(
        \registers[986][6] ), .D(\registers[987][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3356) );
  MX4X1 U5791 ( .A(\registers[988][6] ), .B(\registers[989][6] ), .C(
        \registers[990][6] ), .D(\registers[991][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3355) );
  MX4X1 U5792 ( .A(\registers[976][6] ), .B(\registers[977][6] ), .C(
        \registers[978][6] ), .D(\registers[979][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3358) );
  MX4X1 U5793 ( .A(n3379), .B(n3377), .C(n3378), .D(n3376), .S0(n4615), .S1(
        n4554), .Y(n3380) );
  MX4X1 U5794 ( .A(\registers[920][6] ), .B(\registers[921][6] ), .C(
        \registers[922][6] ), .D(\registers[923][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3377) );
  MX4X1 U5795 ( .A(\registers[924][6] ), .B(\registers[925][6] ), .C(
        \registers[926][6] ), .D(\registers[927][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3376) );
  MX4X1 U5796 ( .A(\registers[912][6] ), .B(\registers[913][6] ), .C(
        \registers[914][6] ), .D(\registers[915][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3379) );
  MX4X1 U5797 ( .A(n3485), .B(n3483), .C(n3484), .D(n3482), .S0(n4617), .S1(
        n4556), .Y(n3486) );
  MX4X1 U5798 ( .A(\registers[600][6] ), .B(\registers[601][6] ), .C(
        \registers[602][6] ), .D(\registers[603][6] ), .S0(n4241), .S1(n4472), 
        .Y(n3483) );
  MX4X1 U5799 ( .A(\registers[604][6] ), .B(\registers[605][6] ), .C(
        \registers[606][6] ), .D(\registers[607][6] ), .S0(n4241), .S1(n4472), 
        .Y(n3482) );
  MX4X1 U5800 ( .A(\registers[592][6] ), .B(\registers[593][6] ), .C(
        \registers[594][6] ), .D(\registers[595][6] ), .S0(n4241), .S1(n4472), 
        .Y(n3485) );
  MX4X1 U5801 ( .A(n3506), .B(n3504), .C(n3505), .D(n3503), .S0(n4617), .S1(
        n4556), .Y(n3507) );
  MX4X1 U5802 ( .A(\registers[536][6] ), .B(\registers[537][6] ), .C(
        \registers[538][6] ), .D(\registers[539][6] ), .S0(n4242), .S1(n4473), 
        .Y(n3504) );
  MX4X1 U5803 ( .A(\registers[540][6] ), .B(\registers[541][6] ), .C(
        \registers[542][6] ), .D(\registers[543][6] ), .S0(n4242), .S1(n4473), 
        .Y(n3503) );
  MX4X1 U5804 ( .A(\registers[528][6] ), .B(\registers[529][6] ), .C(
        \registers[530][6] ), .D(\registers[531][6] ), .S0(n4242), .S1(n4474), 
        .Y(n3506) );
  MX4X1 U5805 ( .A(n3443), .B(n3441), .C(n3442), .D(n3440), .S0(n4616), .S1(
        n4555), .Y(n3444) );
  MX4X1 U5806 ( .A(\registers[728][6] ), .B(\registers[729][6] ), .C(
        \registers[730][6] ), .D(\registers[731][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3441) );
  MX4X1 U5807 ( .A(\registers[732][6] ), .B(\registers[733][6] ), .C(
        \registers[734][6] ), .D(\registers[735][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3440) );
  MX4X1 U5808 ( .A(\registers[720][6] ), .B(\registers[721][6] ), .C(
        \registers[722][6] ), .D(\registers[723][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3443) );
  MX4X1 U5809 ( .A(n3464), .B(n3462), .C(n3463), .D(n3461), .S0(n4617), .S1(
        n4555), .Y(n3465) );
  MX4X1 U5810 ( .A(\registers[664][6] ), .B(\registers[665][6] ), .C(
        \registers[666][6] ), .D(\registers[667][6] ), .S0(n4239), .S1(n4471), 
        .Y(n3462) );
  MX4X1 U5811 ( .A(\registers[668][6] ), .B(\registers[669][6] ), .C(
        \registers[670][6] ), .D(\registers[671][6] ), .S0(n4239), .S1(n4471), 
        .Y(n3461) );
  MX4X1 U5812 ( .A(\registers[656][6] ), .B(\registers[657][6] ), .C(
        \registers[658][6] ), .D(\registers[659][6] ), .S0(n4239), .S1(n4471), 
        .Y(n3464) );
  MX4X1 U5813 ( .A(n3910), .B(n3908), .C(n3909), .D(n3907), .S0(n4624), .S1(
        n4558), .Y(n3911) );
  MX4X1 U5814 ( .A(\registers[344][7] ), .B(\registers[345][7] ), .C(
        \registers[346][7] ), .D(\registers[347][7] ), .S0(n4267), .S1(n4492), 
        .Y(n3908) );
  MX4X1 U5815 ( .A(\registers[348][7] ), .B(\registers[349][7] ), .C(
        \registers[350][7] ), .D(\registers[351][7] ), .S0(n4267), .S1(n4479), 
        .Y(n3907) );
  MX4X1 U5816 ( .A(\registers[336][7] ), .B(\registers[337][7] ), .C(
        \registers[338][7] ), .D(\registers[339][7] ), .S0(n4267), .S1(n4478), 
        .Y(n3910) );
  MX4X1 U5817 ( .A(n3931), .B(n3929), .C(n3930), .D(n3928), .S0(n4624), .S1(
        n4558), .Y(n3932) );
  MX4X1 U5818 ( .A(\registers[280][7] ), .B(\registers[281][7] ), .C(
        \registers[282][7] ), .D(\registers[283][7] ), .S0(n4269), .S1(n4497), 
        .Y(n3929) );
  MX4X1 U5819 ( .A(\registers[284][7] ), .B(\registers[285][7] ), .C(
        \registers[286][7] ), .D(\registers[287][7] ), .S0(n4269), .S1(n4497), 
        .Y(n3928) );
  MX4X1 U5820 ( .A(\registers[272][7] ), .B(\registers[273][7] ), .C(
        \registers[274][7] ), .D(\registers[275][7] ), .S0(n4269), .S1(n4497), 
        .Y(n3931) );
  MX4X1 U5821 ( .A(n3868), .B(n3866), .C(n3867), .D(n3865), .S0(n4623), .S1(
        n4530), .Y(n3869) );
  MX4X1 U5822 ( .A(\registers[472][7] ), .B(\registers[473][7] ), .C(
        \registers[474][7] ), .D(\registers[475][7] ), .S0(n4265), .S1(n4494), 
        .Y(n3866) );
  MX4X1 U5823 ( .A(\registers[476][7] ), .B(\registers[477][7] ), .C(
        \registers[478][7] ), .D(\registers[479][7] ), .S0(n4265), .S1(n4494), 
        .Y(n3865) );
  MX4X1 U5824 ( .A(\registers[464][7] ), .B(\registers[465][7] ), .C(
        \registers[466][7] ), .D(\registers[467][7] ), .S0(n4265), .S1(n4495), 
        .Y(n3868) );
  MX4X1 U5825 ( .A(n3889), .B(n3887), .C(n3888), .D(n3886), .S0(n4623), .S1(
        n4558), .Y(n3890) );
  MX4X1 U5826 ( .A(\registers[408][7] ), .B(\registers[409][7] ), .C(
        \registers[410][7] ), .D(\registers[411][7] ), .S0(n4266), .S1(n4496), 
        .Y(n3887) );
  MX4X1 U5827 ( .A(\registers[412][7] ), .B(\registers[413][7] ), .C(
        \registers[414][7] ), .D(\registers[415][7] ), .S0(n4266), .S1(n4496), 
        .Y(n3886) );
  MX4X1 U5828 ( .A(\registers[400][7] ), .B(\registers[401][7] ), .C(
        \registers[402][7] ), .D(\registers[403][7] ), .S0(n4266), .S1(n4496), 
        .Y(n3889) );
  MX4X1 U5829 ( .A(n3995), .B(n3993), .C(n3994), .D(n3992), .S0(n4619), .S1(
        n4559), .Y(n3996) );
  MX4X1 U5830 ( .A(\registers[88][7] ), .B(\registers[89][7] ), .C(
        \registers[90][7] ), .D(\registers[91][7] ), .S0(n4273), .S1(n4463), 
        .Y(n3993) );
  MX4X1 U5831 ( .A(\registers[92][7] ), .B(\registers[93][7] ), .C(
        \registers[94][7] ), .D(\registers[95][7] ), .S0(n4273), .S1(n4462), 
        .Y(n3992) );
  MX4X1 U5832 ( .A(\registers[80][7] ), .B(\registers[81][7] ), .C(
        \registers[82][7] ), .D(\registers[83][7] ), .S0(n4273), .S1(n4466), 
        .Y(n3995) );
  MX4X1 U5833 ( .A(n4016), .B(n4014), .C(n4015), .D(n4013), .S0(N71), .S1(
        n4559), .Y(n4017) );
  MX4X1 U5834 ( .A(\registers[24][7] ), .B(\registers[25][7] ), .C(
        \registers[26][7] ), .D(\registers[27][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4014) );
  MX4X1 U5835 ( .A(\registers[28][7] ), .B(\registers[29][7] ), .C(
        \registers[30][7] ), .D(\registers[31][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4013) );
  MX4X1 U5836 ( .A(\registers[16][7] ), .B(\registers[17][7] ), .C(
        \registers[18][7] ), .D(\registers[19][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4016) );
  MX4X1 U5837 ( .A(n3953), .B(n3951), .C(n3952), .D(n3950), .S0(n4624), .S1(
        n4558), .Y(n3954) );
  MX4X1 U5838 ( .A(\registers[216][7] ), .B(\registers[217][7] ), .C(
        \registers[218][7] ), .D(\registers[219][7] ), .S0(n4270), .S1(n4498), 
        .Y(n3951) );
  MX4X1 U5839 ( .A(\registers[220][7] ), .B(\registers[221][7] ), .C(
        \registers[222][7] ), .D(\registers[223][7] ), .S0(n4270), .S1(n4498), 
        .Y(n3950) );
  MX4X1 U5840 ( .A(\registers[208][7] ), .B(\registers[209][7] ), .C(
        \registers[210][7] ), .D(\registers[211][7] ), .S0(n4270), .S1(n4498), 
        .Y(n3953) );
  MX4X1 U5841 ( .A(n3974), .B(n3972), .C(n3973), .D(n3971), .S0(N71), .S1(
        n4559), .Y(n3975) );
  MX4X1 U5842 ( .A(\registers[152][7] ), .B(\registers[153][7] ), .C(
        \registers[154][7] ), .D(\registers[155][7] ), .S0(n4271), .S1(n4500), 
        .Y(n3972) );
  MX4X1 U5843 ( .A(\registers[156][7] ), .B(\registers[157][7] ), .C(
        \registers[158][7] ), .D(\registers[159][7] ), .S0(n4271), .S1(n4499), 
        .Y(n3971) );
  MX4X1 U5844 ( .A(\registers[144][7] ), .B(\registers[145][7] ), .C(
        \registers[146][7] ), .D(\registers[147][7] ), .S0(n4271), .S1(n4500), 
        .Y(n3974) );
  MX4X1 U5845 ( .A(n3740), .B(n3738), .C(n3739), .D(n3737), .S0(n4621), .S1(
        n4540), .Y(n3741) );
  MX4X1 U5846 ( .A(\registers[856][7] ), .B(\registers[857][7] ), .C(
        \registers[858][7] ), .D(\registers[859][7] ), .S0(n4257), .S1(n4487), 
        .Y(n3738) );
  MX4X1 U5847 ( .A(\registers[860][7] ), .B(\registers[861][7] ), .C(
        \registers[862][7] ), .D(\registers[863][7] ), .S0(n4257), .S1(n4487), 
        .Y(n3737) );
  MX4X1 U5848 ( .A(\registers[848][7] ), .B(\registers[849][7] ), .C(
        \registers[850][7] ), .D(\registers[851][7] ), .S0(n4257), .S1(n4487), 
        .Y(n3740) );
  MX4X1 U5849 ( .A(n3761), .B(n3759), .C(n3760), .D(n3758), .S0(n4621), .S1(
        n4528), .Y(n3762) );
  MX4X1 U5850 ( .A(\registers[792][7] ), .B(\registers[793][7] ), .C(
        \registers[794][7] ), .D(\registers[795][7] ), .S0(n4258), .S1(n4488), 
        .Y(n3759) );
  MX4X1 U5851 ( .A(\registers[796][7] ), .B(\registers[797][7] ), .C(
        \registers[798][7] ), .D(\registers[799][7] ), .S0(n4258), .S1(n4488), 
        .Y(n3758) );
  MX4X1 U5852 ( .A(\registers[784][7] ), .B(\registers[785][7] ), .C(
        \registers[786][7] ), .D(\registers[787][7] ), .S0(n4258), .S1(n4488), 
        .Y(n3761) );
  MX4X1 U5853 ( .A(n3698), .B(n3696), .C(n3697), .D(n3695), .S0(n4620), .S1(
        n4544), .Y(n3699) );
  MX4X1 U5854 ( .A(\registers[984][7] ), .B(\registers[985][7] ), .C(
        \registers[986][7] ), .D(\registers[987][7] ), .S0(n4254), .S1(n4485), 
        .Y(n3696) );
  MX4X1 U5855 ( .A(\registers[988][7] ), .B(\registers[989][7] ), .C(
        \registers[990][7] ), .D(\registers[991][7] ), .S0(n4254), .S1(n4484), 
        .Y(n3695) );
  MX4X1 U5856 ( .A(\registers[976][7] ), .B(\registers[977][7] ), .C(
        \registers[978][7] ), .D(\registers[979][7] ), .S0(n4254), .S1(n4485), 
        .Y(n3698) );
  MX4X1 U5857 ( .A(n3719), .B(n3717), .C(n3718), .D(n3716), .S0(n4621), .S1(
        n4538), .Y(n3720) );
  MX4X1 U5858 ( .A(\registers[920][7] ), .B(\registers[921][7] ), .C(
        \registers[922][7] ), .D(\registers[923][7] ), .S0(n4255), .S1(n4486), 
        .Y(n3717) );
  MX4X1 U5859 ( .A(\registers[924][7] ), .B(\registers[925][7] ), .C(
        \registers[926][7] ), .D(\registers[927][7] ), .S0(n4255), .S1(n4486), 
        .Y(n3716) );
  MX4X1 U5860 ( .A(\registers[912][7] ), .B(\registers[913][7] ), .C(
        \registers[914][7] ), .D(\registers[915][7] ), .S0(n4255), .S1(n4486), 
        .Y(n3719) );
  MX4X1 U5861 ( .A(n3825), .B(n3823), .C(n3824), .D(n3822), .S0(n4622), .S1(
        n4536), .Y(n3826) );
  MX4X1 U5862 ( .A(\registers[600][7] ), .B(\registers[601][7] ), .C(
        \registers[602][7] ), .D(\registers[603][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3823) );
  MX4X1 U5863 ( .A(\registers[604][7] ), .B(\registers[605][7] ), .C(
        \registers[606][7] ), .D(\registers[607][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3822) );
  MX4X1 U5864 ( .A(\registers[592][7] ), .B(\registers[593][7] ), .C(
        \registers[594][7] ), .D(\registers[595][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3825) );
  MX4X1 U5865 ( .A(n3846), .B(n3844), .C(n3845), .D(n3843), .S0(n4623), .S1(
        n4543), .Y(n3847) );
  MX4X1 U5866 ( .A(\registers[536][7] ), .B(\registers[537][7] ), .C(
        \registers[538][7] ), .D(\registers[539][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3844) );
  MX4X1 U5867 ( .A(\registers[540][7] ), .B(\registers[541][7] ), .C(
        \registers[542][7] ), .D(\registers[543][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3843) );
  MX4X1 U5868 ( .A(\registers[528][7] ), .B(\registers[529][7] ), .C(
        \registers[530][7] ), .D(\registers[531][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3846) );
  MX4X1 U5869 ( .A(n3783), .B(n3781), .C(n3782), .D(n3780), .S0(n4622), .S1(
        n4537), .Y(n3784) );
  MX4X1 U5870 ( .A(\registers[728][7] ), .B(\registers[729][7] ), .C(
        \registers[730][7] ), .D(\registers[731][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3781) );
  MX4X1 U5871 ( .A(\registers[732][7] ), .B(\registers[733][7] ), .C(
        \registers[734][7] ), .D(\registers[735][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3780) );
  MX4X1 U5872 ( .A(\registers[720][7] ), .B(\registers[721][7] ), .C(
        \registers[722][7] ), .D(\registers[723][7] ), .S0(n4259), .S1(n4490), 
        .Y(n3783) );
  MX4X1 U5873 ( .A(n3804), .B(n3802), .C(n3803), .D(n3801), .S0(n4622), .S1(
        n4539), .Y(n3805) );
  MX4X1 U5874 ( .A(\registers[664][7] ), .B(\registers[665][7] ), .C(
        \registers[666][7] ), .D(\registers[667][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3802) );
  MX4X1 U5875 ( .A(\registers[668][7] ), .B(\registers[669][7] ), .C(
        \registers[670][7] ), .D(\registers[671][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3801) );
  MX4X1 U5876 ( .A(\registers[656][7] ), .B(\registers[657][7] ), .C(
        \registers[658][7] ), .D(\registers[659][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3804) );
  MX4X1 U5877 ( .A(n4875), .B(n4873), .C(n4874), .D(n4872), .S0(n7958), .S1(
        n7869), .Y(n4876) );
  MX4X1 U5878 ( .A(\registers[344][0] ), .B(\registers[345][0] ), .C(
        \registers[346][0] ), .D(\registers[347][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4873) );
  MX4X1 U5879 ( .A(\registers[348][0] ), .B(\registers[349][0] ), .C(
        \registers[350][0] ), .D(\registers[351][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4872) );
  MX4X1 U5880 ( .A(\registers[336][0] ), .B(\registers[337][0] ), .C(
        \registers[338][0] ), .D(\registers[339][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4875) );
  MX4X1 U5881 ( .A(n4896), .B(n4894), .C(n4895), .D(n4893), .S0(n7930), .S1(
        n7870), .Y(n4897) );
  MX4X1 U5882 ( .A(\registers[280][0] ), .B(\registers[281][0] ), .C(
        \registers[282][0] ), .D(\registers[283][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4894) );
  MX4X1 U5883 ( .A(\registers[284][0] ), .B(\registers[285][0] ), .C(
        \registers[286][0] ), .D(\registers[287][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4893) );
  MX4X1 U5884 ( .A(\registers[272][0] ), .B(\registers[273][0] ), .C(
        \registers[274][0] ), .D(\registers[275][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4896) );
  MX4X1 U5885 ( .A(n4833), .B(n4831), .C(n4832), .D(n4830), .S0(n7947), .S1(
        n7869), .Y(n4834) );
  MX4X1 U5886 ( .A(\registers[472][0] ), .B(\registers[473][0] ), .C(
        \registers[474][0] ), .D(\registers[475][0] ), .S0(n7458), .S1(n7701), 
        .Y(n4831) );
  MX4X1 U5887 ( .A(\registers[476][0] ), .B(\registers[477][0] ), .C(
        \registers[478][0] ), .D(\registers[479][0] ), .S0(n7458), .S1(n7700), 
        .Y(n4830) );
  MX4X1 U5888 ( .A(\registers[464][0] ), .B(\registers[465][0] ), .C(
        \registers[466][0] ), .D(\registers[467][0] ), .S0(n7458), .S1(n7701), 
        .Y(n4833) );
  MX4X1 U5889 ( .A(n4854), .B(n4852), .C(n4853), .D(n4851), .S0(n7950), .S1(
        n7869), .Y(n4855) );
  MX4X1 U5890 ( .A(\registers[408][0] ), .B(\registers[409][0] ), .C(
        \registers[410][0] ), .D(\registers[411][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4852) );
  MX4X1 U5891 ( .A(\registers[412][0] ), .B(\registers[413][0] ), .C(
        \registers[414][0] ), .D(\registers[415][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4851) );
  MX4X1 U5892 ( .A(\registers[400][0] ), .B(\registers[401][0] ), .C(
        \registers[402][0] ), .D(\registers[403][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4854) );
  MX4X1 U5893 ( .A(n4960), .B(n4958), .C(n4959), .D(n4957), .S0(n7931), .S1(
        n7871), .Y(n4961) );
  MX4X1 U5894 ( .A(\registers[88][0] ), .B(\registers[89][0] ), .C(
        \registers[90][0] ), .D(\registers[91][0] ), .S0(n7466), .S1(n7708), 
        .Y(n4958) );
  MX4X1 U5895 ( .A(\registers[92][0] ), .B(\registers[93][0] ), .C(
        \registers[94][0] ), .D(\registers[95][0] ), .S0(n7466), .S1(n7708), 
        .Y(n4957) );
  MX4X1 U5896 ( .A(\registers[80][0] ), .B(\registers[81][0] ), .C(
        \registers[82][0] ), .D(\registers[83][0] ), .S0(n7466), .S1(n7708), 
        .Y(n4960) );
  MX4X1 U5897 ( .A(n4981), .B(n4979), .C(n4980), .D(n4978), .S0(n7931), .S1(
        n7871), .Y(n4982) );
  MX4X1 U5898 ( .A(\registers[24][0] ), .B(\registers[25][0] ), .C(
        \registers[26][0] ), .D(\registers[27][0] ), .S0(n7468), .S1(n7709), 
        .Y(n4979) );
  MX4X1 U5899 ( .A(\registers[28][0] ), .B(\registers[29][0] ), .C(
        \registers[30][0] ), .D(\registers[31][0] ), .S0(n7468), .S1(n7709), 
        .Y(n4978) );
  MX4X1 U5900 ( .A(\registers[16][0] ), .B(\registers[17][0] ), .C(
        \registers[18][0] ), .D(\registers[19][0] ), .S0(n7468), .S1(n7709), 
        .Y(n4981) );
  MX4X1 U5901 ( .A(n4918), .B(n4916), .C(n4917), .D(n4915), .S0(n7930), .S1(
        n7870), .Y(n4919) );
  MX4X1 U5902 ( .A(\registers[216][0] ), .B(\registers[217][0] ), .C(
        \registers[218][0] ), .D(\registers[219][0] ), .S0(n7464), .S1(n7705), 
        .Y(n4916) );
  MX4X1 U5903 ( .A(\registers[220][0] ), .B(\registers[221][0] ), .C(
        \registers[222][0] ), .D(\registers[223][0] ), .S0(n7464), .S1(n7705), 
        .Y(n4915) );
  MX4X1 U5904 ( .A(\registers[208][0] ), .B(\registers[209][0] ), .C(
        \registers[210][0] ), .D(\registers[211][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4918) );
  MX4X1 U5905 ( .A(n4939), .B(n4937), .C(n4938), .D(n4936), .S0(n7930), .S1(
        n7870), .Y(n4940) );
  MX4X1 U5906 ( .A(\registers[152][0] ), .B(\registers[153][0] ), .C(
        \registers[154][0] ), .D(\registers[155][0] ), .S0(n7465), .S1(n7707), 
        .Y(n4937) );
  MX4X1 U5907 ( .A(\registers[156][0] ), .B(\registers[157][0] ), .C(
        \registers[158][0] ), .D(\registers[159][0] ), .S0(n7465), .S1(n7707), 
        .Y(n4936) );
  MX4X1 U5908 ( .A(\registers[144][0] ), .B(\registers[145][0] ), .C(
        \registers[146][0] ), .D(\registers[147][0] ), .S0(n7465), .S1(n7707), 
        .Y(n4939) );
  MX4X1 U5909 ( .A(n4705), .B(n4703), .C(n4704), .D(n4702), .S0(n7933), .S1(
        n7867), .Y(n4706) );
  MX4X1 U5910 ( .A(\registers[856][0] ), .B(\registers[857][0] ), .C(
        \registers[858][0] ), .D(\registers[859][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4703) );
  MX4X1 U5911 ( .A(\registers[860][0] ), .B(\registers[861][0] ), .C(
        \registers[862][0] ), .D(\registers[863][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4702) );
  MX4X1 U5912 ( .A(\registers[848][0] ), .B(\registers[849][0] ), .C(
        \registers[850][0] ), .D(\registers[851][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4705) );
  MX4X1 U5913 ( .A(n4726), .B(n4724), .C(n4725), .D(n4723), .S0(n7934), .S1(
        n7867), .Y(n4727) );
  MX4X1 U5914 ( .A(\registers[792][0] ), .B(\registers[793][0] ), .C(
        \registers[794][0] ), .D(\registers[795][0] ), .S0(n7452), .S1(n7694), 
        .Y(n4724) );
  MX4X1 U5915 ( .A(\registers[796][0] ), .B(\registers[797][0] ), .C(
        \registers[798][0] ), .D(\registers[799][0] ), .S0(n7452), .S1(n7694), 
        .Y(n4723) );
  MX4X1 U5916 ( .A(\registers[784][0] ), .B(\registers[785][0] ), .C(
        \registers[786][0] ), .D(\registers[787][0] ), .S0(n7452), .S1(n7695), 
        .Y(n4726) );
  MX4X1 U5917 ( .A(n4790), .B(n4788), .C(n4789), .D(n4787), .S0(n7948), .S1(
        n7868), .Y(n4791) );
  MX4X1 U5918 ( .A(\registers[600][0] ), .B(\registers[601][0] ), .C(
        \registers[602][0] ), .D(\registers[603][0] ), .S0(n7456), .S1(n7698), 
        .Y(n4788) );
  MX4X1 U5919 ( .A(\registers[604][0] ), .B(\registers[605][0] ), .C(
        \registers[606][0] ), .D(\registers[607][0] ), .S0(n7456), .S1(n7698), 
        .Y(n4787) );
  MX4X1 U5920 ( .A(\registers[592][0] ), .B(\registers[593][0] ), .C(
        \registers[594][0] ), .D(\registers[595][0] ), .S0(n7456), .S1(n7698), 
        .Y(n4790) );
  MX4X1 U5921 ( .A(n4811), .B(n4809), .C(n4810), .D(n4808), .S0(n7949), .S1(
        n7868), .Y(n4812) );
  MX4X1 U5922 ( .A(\registers[536][0] ), .B(\registers[537][0] ), .C(
        \registers[538][0] ), .D(\registers[539][0] ), .S0(n7457), .S1(n7699), 
        .Y(n4809) );
  MX4X1 U5923 ( .A(\registers[540][0] ), .B(\registers[541][0] ), .C(
        \registers[542][0] ), .D(\registers[543][0] ), .S0(n7457), .S1(n7699), 
        .Y(n4808) );
  MX4X1 U5924 ( .A(\registers[528][0] ), .B(\registers[529][0] ), .C(
        \registers[530][0] ), .D(\registers[531][0] ), .S0(n7457), .S1(n7699), 
        .Y(n4811) );
  MX4X1 U5925 ( .A(n4748), .B(n4746), .C(n4747), .D(n4745), .S0(n7931), .S1(
        n7868), .Y(n4749) );
  MX4X1 U5926 ( .A(\registers[728][0] ), .B(\registers[729][0] ), .C(
        \registers[730][0] ), .D(\registers[731][0] ), .S0(n7453), .S1(n7696), 
        .Y(n4746) );
  MX4X1 U5927 ( .A(\registers[732][0] ), .B(\registers[733][0] ), .C(
        \registers[734][0] ), .D(\registers[735][0] ), .S0(n7453), .S1(n7696), 
        .Y(n4745) );
  MX4X1 U5928 ( .A(\registers[720][0] ), .B(\registers[721][0] ), .C(
        \registers[722][0] ), .D(\registers[723][0] ), .S0(n7453), .S1(n7696), 
        .Y(n4748) );
  MX4X1 U5929 ( .A(n4769), .B(n4767), .C(n4768), .D(n4766), .S0(n7954), .S1(
        n7868), .Y(n4770) );
  MX4X1 U5930 ( .A(\registers[664][0] ), .B(\registers[665][0] ), .C(
        \registers[666][0] ), .D(\registers[667][0] ), .S0(n7454), .S1(n7697), 
        .Y(n4767) );
  MX4X1 U5931 ( .A(\registers[668][0] ), .B(\registers[669][0] ), .C(
        \registers[670][0] ), .D(\registers[671][0] ), .S0(n7454), .S1(n7697), 
        .Y(n4766) );
  MX4X1 U5932 ( .A(\registers[656][0] ), .B(\registers[657][0] ), .C(
        \registers[658][0] ), .D(\registers[659][0] ), .S0(n7454), .S1(n7697), 
        .Y(n4769) );
  MX4X1 U5933 ( .A(n5215), .B(n5213), .C(n5214), .D(n5212), .S0(n7935), .S1(
        n7874), .Y(n5216) );
  MX4X1 U5934 ( .A(\registers[344][1] ), .B(\registers[345][1] ), .C(
        \registers[346][1] ), .D(\registers[347][1] ), .S0(n7482), .S1(n7723), 
        .Y(n5213) );
  MX4X1 U5935 ( .A(\registers[348][1] ), .B(\registers[349][1] ), .C(
        \registers[350][1] ), .D(\registers[351][1] ), .S0(n7482), .S1(n7723), 
        .Y(n5212) );
  MX4X1 U5936 ( .A(\registers[336][1] ), .B(\registers[337][1] ), .C(
        \registers[338][1] ), .D(\registers[339][1] ), .S0(n7482), .S1(n7723), 
        .Y(n5215) );
  MX4X1 U5937 ( .A(n5236), .B(n5234), .C(n5235), .D(n5233), .S0(n7935), .S1(
        n7875), .Y(n5237) );
  MX4X1 U5938 ( .A(\registers[280][1] ), .B(\registers[281][1] ), .C(
        \registers[282][1] ), .D(\registers[283][1] ), .S0(n7484), .S1(n7724), 
        .Y(n5234) );
  MX4X1 U5939 ( .A(\registers[284][1] ), .B(\registers[285][1] ), .C(
        \registers[286][1] ), .D(\registers[287][1] ), .S0(n7484), .S1(n7724), 
        .Y(n5233) );
  MX4X1 U5940 ( .A(\registers[272][1] ), .B(\registers[273][1] ), .C(
        \registers[274][1] ), .D(\registers[275][1] ), .S0(n7484), .S1(n7724), 
        .Y(n5236) );
  MX4X1 U5941 ( .A(n5173), .B(n5171), .C(n5172), .D(n5170), .S0(n7934), .S1(
        n7874), .Y(n5174) );
  MX4X1 U5942 ( .A(\registers[472][1] ), .B(\registers[473][1] ), .C(
        \registers[474][1] ), .D(\registers[475][1] ), .S0(n7480), .S1(n7720), 
        .Y(n5171) );
  MX4X1 U5943 ( .A(\registers[476][1] ), .B(\registers[477][1] ), .C(
        \registers[478][1] ), .D(\registers[479][1] ), .S0(n7480), .S1(n7720), 
        .Y(n5170) );
  MX4X1 U5944 ( .A(\registers[464][1] ), .B(\registers[465][1] ), .C(
        \registers[466][1] ), .D(\registers[467][1] ), .S0(n7480), .S1(n7720), 
        .Y(n5173) );
  MX4X1 U5945 ( .A(n5194), .B(n5192), .C(n5193), .D(n5191), .S0(n7934), .S1(
        n7874), .Y(n5195) );
  MX4X1 U5946 ( .A(\registers[408][1] ), .B(\registers[409][1] ), .C(
        \registers[410][1] ), .D(\registers[411][1] ), .S0(n7481), .S1(n7721), 
        .Y(n5192) );
  MX4X1 U5947 ( .A(\registers[412][1] ), .B(\registers[413][1] ), .C(
        \registers[414][1] ), .D(\registers[415][1] ), .S0(n7481), .S1(n7721), 
        .Y(n5191) );
  MX4X1 U5948 ( .A(\registers[400][1] ), .B(\registers[401][1] ), .C(
        \registers[402][1] ), .D(\registers[403][1] ), .S0(n7481), .S1(n7722), 
        .Y(n5194) );
  MX4X1 U5949 ( .A(n5300), .B(n5298), .C(n5299), .D(n5297), .S0(n7936), .S1(
        n7876), .Y(n5301) );
  MX4X1 U5950 ( .A(\registers[88][1] ), .B(\registers[89][1] ), .C(
        \registers[90][1] ), .D(\registers[91][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5298) );
  MX4X1 U5951 ( .A(\registers[92][1] ), .B(\registers[93][1] ), .C(
        \registers[94][1] ), .D(\registers[95][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5297) );
  MX4X1 U5952 ( .A(\registers[80][1] ), .B(\registers[81][1] ), .C(
        \registers[82][1] ), .D(\registers[83][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5300) );
  MX4X1 U5953 ( .A(n5321), .B(n5319), .C(n5320), .D(n5318), .S0(n7936), .S1(
        n7876), .Y(n5322) );
  MX4X1 U5954 ( .A(\registers[24][1] ), .B(\registers[25][1] ), .C(
        \registers[26][1] ), .D(\registers[27][1] ), .S0(n7489), .S1(n7729), 
        .Y(n5319) );
  MX4X1 U5955 ( .A(\registers[28][1] ), .B(\registers[29][1] ), .C(
        \registers[30][1] ), .D(\registers[31][1] ), .S0(n7489), .S1(n7729), 
        .Y(n5318) );
  MX4X1 U5956 ( .A(\registers[16][1] ), .B(\registers[17][1] ), .C(
        \registers[18][1] ), .D(\registers[19][1] ), .S0(n7489), .S1(n7729), 
        .Y(n5321) );
  MX4X1 U5957 ( .A(n5258), .B(n5256), .C(n5257), .D(n5255), .S0(n7935), .S1(
        n7875), .Y(n5259) );
  MX4X1 U5958 ( .A(\registers[216][1] ), .B(\registers[217][1] ), .C(
        \registers[218][1] ), .D(\registers[219][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5256) );
  MX4X1 U5959 ( .A(\registers[220][1] ), .B(\registers[221][1] ), .C(
        \registers[222][1] ), .D(\registers[223][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5255) );
  MX4X1 U5960 ( .A(\registers[208][1] ), .B(\registers[209][1] ), .C(
        \registers[210][1] ), .D(\registers[211][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5258) );
  MX4X1 U5961 ( .A(n5279), .B(n5277), .C(n5278), .D(n5276), .S0(n7936), .S1(
        n7875), .Y(n5280) );
  MX4X1 U5962 ( .A(\registers[152][1] ), .B(\registers[153][1] ), .C(
        \registers[154][1] ), .D(\registers[155][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5277) );
  MX4X1 U5963 ( .A(\registers[156][1] ), .B(\registers[157][1] ), .C(
        \registers[158][1] ), .D(\registers[159][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5276) );
  MX4X1 U5964 ( .A(\registers[144][1] ), .B(\registers[145][1] ), .C(
        \registers[146][1] ), .D(\registers[147][1] ), .S0(n7486), .S1(n7727), 
        .Y(n5279) );
  MX4X1 U5965 ( .A(n5045), .B(n5043), .C(n5044), .D(n5042), .S0(n7932), .S1(
        n7872), .Y(n5046) );
  MX4X1 U5966 ( .A(\registers[856][1] ), .B(\registers[857][1] ), .C(
        \registers[858][1] ), .D(\registers[859][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5043) );
  MX4X1 U5967 ( .A(\registers[860][1] ), .B(\registers[861][1] ), .C(
        \registers[862][1] ), .D(\registers[863][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5042) );
  MX4X1 U5968 ( .A(\registers[848][1] ), .B(\registers[849][1] ), .C(
        \registers[850][1] ), .D(\registers[851][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5045) );
  MX4X1 U5969 ( .A(n5066), .B(n5064), .C(n5065), .D(n5063), .S0(n7932), .S1(
        n7872), .Y(n5067) );
  MX4X1 U5970 ( .A(\registers[792][1] ), .B(\registers[793][1] ), .C(
        \registers[794][1] ), .D(\registers[795][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5064) );
  MX4X1 U5971 ( .A(\registers[796][1] ), .B(\registers[797][1] ), .C(
        \registers[798][1] ), .D(\registers[799][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5063) );
  MX4X1 U5972 ( .A(\registers[784][1] ), .B(\registers[785][1] ), .C(
        \registers[786][1] ), .D(\registers[787][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5066) );
  MX4X1 U5973 ( .A(n5003), .B(n5001), .C(n5002), .D(n5000), .S0(n7931), .S1(
        n7871), .Y(n5004) );
  MX4X1 U5974 ( .A(\registers[984][1] ), .B(\registers[985][1] ), .C(
        \registers[986][1] ), .D(\registers[987][1] ), .S0(n7469), .S1(n7710), 
        .Y(n5001) );
  MX4X1 U5975 ( .A(\registers[988][1] ), .B(\registers[989][1] ), .C(
        \registers[990][1] ), .D(\registers[991][1] ), .S0(n7469), .S1(n7710), 
        .Y(n5000) );
  MX4X1 U5976 ( .A(\registers[976][1] ), .B(\registers[977][1] ), .C(
        \registers[978][1] ), .D(\registers[979][1] ), .S0(n7469), .S1(n7711), 
        .Y(n5003) );
  MX4X1 U5977 ( .A(n5024), .B(n5022), .C(n5023), .D(n5021), .S0(n7932), .S1(
        n7872), .Y(n5025) );
  MX4X1 U5978 ( .A(\registers[920][1] ), .B(\registers[921][1] ), .C(
        \registers[922][1] ), .D(\registers[923][1] ), .S0(n7470), .S1(n7712), 
        .Y(n5022) );
  MX4X1 U5979 ( .A(\registers[924][1] ), .B(\registers[925][1] ), .C(
        \registers[926][1] ), .D(\registers[927][1] ), .S0(n7470), .S1(n7712), 
        .Y(n5021) );
  MX4X1 U5980 ( .A(\registers[912][1] ), .B(\registers[913][1] ), .C(
        \registers[914][1] ), .D(\registers[915][1] ), .S0(n7470), .S1(n7712), 
        .Y(n5024) );
  MX4X1 U5981 ( .A(n5130), .B(n5128), .C(n5129), .D(n5127), .S0(n7933), .S1(
        n7873), .Y(n5131) );
  MX4X1 U5982 ( .A(\registers[600][1] ), .B(\registers[601][1] ), .C(
        \registers[602][1] ), .D(\registers[603][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5128) );
  MX4X1 U5983 ( .A(\registers[604][1] ), .B(\registers[605][1] ), .C(
        \registers[606][1] ), .D(\registers[607][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5127) );
  MX4X1 U5984 ( .A(\registers[592][1] ), .B(\registers[593][1] ), .C(
        \registers[594][1] ), .D(\registers[595][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5130) );
  MX4X1 U5985 ( .A(n5151), .B(n5149), .C(n5150), .D(n5148), .S0(n7934), .S1(
        n7873), .Y(n5152) );
  MX4X1 U5986 ( .A(\registers[536][1] ), .B(\registers[537][1] ), .C(
        \registers[538][1] ), .D(\registers[539][1] ), .S0(n7478), .S1(n7719), 
        .Y(n5149) );
  MX4X1 U5987 ( .A(\registers[540][1] ), .B(\registers[541][1] ), .C(
        \registers[542][1] ), .D(\registers[543][1] ), .S0(n7478), .S1(n7719), 
        .Y(n5148) );
  MX4X1 U5988 ( .A(\registers[528][1] ), .B(\registers[529][1] ), .C(
        \registers[530][1] ), .D(\registers[531][1] ), .S0(n7478), .S1(n7719), 
        .Y(n5151) );
  MX4X1 U5989 ( .A(n5088), .B(n5086), .C(n5087), .D(n5085), .S0(n7933), .S1(
        n7872), .Y(n5089) );
  MX4X1 U5990 ( .A(\registers[728][1] ), .B(\registers[729][1] ), .C(
        \registers[730][1] ), .D(\registers[731][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5086) );
  MX4X1 U5991 ( .A(\registers[732][1] ), .B(\registers[733][1] ), .C(
        \registers[734][1] ), .D(\registers[735][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5085) );
  MX4X1 U5992 ( .A(\registers[720][1] ), .B(\registers[721][1] ), .C(
        \registers[722][1] ), .D(\registers[723][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5088) );
  MX4X1 U5993 ( .A(n5109), .B(n5107), .C(n5108), .D(n5106), .S0(n7933), .S1(
        n7873), .Y(n5110) );
  MX4X1 U5994 ( .A(\registers[664][1] ), .B(\registers[665][1] ), .C(
        \registers[666][1] ), .D(\registers[667][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5107) );
  MX4X1 U5995 ( .A(\registers[668][1] ), .B(\registers[669][1] ), .C(
        \registers[670][1] ), .D(\registers[671][1] ), .S0(n7476), .S1(n7716), 
        .Y(n5106) );
  MX4X1 U5996 ( .A(\registers[656][1] ), .B(\registers[657][1] ), .C(
        \registers[658][1] ), .D(\registers[659][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5109) );
  MX4X1 U5997 ( .A(n5555), .B(n5553), .C(n5554), .D(n5552), .S0(n7940), .S1(
        n7879), .Y(n5556) );
  MX4X1 U5998 ( .A(\registers[344][2] ), .B(\registers[345][2] ), .C(
        \registers[346][2] ), .D(\registers[347][2] ), .S0(n7504), .S1(n7742), 
        .Y(n5553) );
  MX4X1 U5999 ( .A(\registers[348][2] ), .B(\registers[349][2] ), .C(
        \registers[350][2] ), .D(\registers[351][2] ), .S0(n7504), .S1(n7742), 
        .Y(n5552) );
  MX4X1 U6000 ( .A(\registers[336][2] ), .B(\registers[337][2] ), .C(
        \registers[338][2] ), .D(\registers[339][2] ), .S0(n7504), .S1(n7743), 
        .Y(n5555) );
  MX4X1 U6001 ( .A(n5576), .B(n5574), .C(n5575), .D(n5573), .S0(n7940), .S1(
        n7880), .Y(n5577) );
  MX4X1 U6002 ( .A(\registers[280][2] ), .B(\registers[281][2] ), .C(
        \registers[282][2] ), .D(\registers[283][2] ), .S0(n7505), .S1(n7744), 
        .Y(n5574) );
  MX4X1 U6003 ( .A(\registers[284][2] ), .B(\registers[285][2] ), .C(
        \registers[286][2] ), .D(\registers[287][2] ), .S0(n7505), .S1(n7744), 
        .Y(n5573) );
  MX4X1 U6004 ( .A(\registers[272][2] ), .B(\registers[273][2] ), .C(
        \registers[274][2] ), .D(\registers[275][2] ), .S0(n7505), .S1(n7744), 
        .Y(n5576) );
  MX4X1 U6005 ( .A(n5513), .B(n5511), .C(n5512), .D(n5510), .S0(n7939), .S1(
        n7879), .Y(n5514) );
  MX4X1 U6006 ( .A(\registers[472][2] ), .B(\registers[473][2] ), .C(
        \registers[474][2] ), .D(\registers[475][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5511) );
  MX4X1 U6007 ( .A(\registers[476][2] ), .B(\registers[477][2] ), .C(
        \registers[478][2] ), .D(\registers[479][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5510) );
  MX4X1 U6008 ( .A(\registers[464][2] ), .B(\registers[465][2] ), .C(
        \registers[466][2] ), .D(\registers[467][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5513) );
  MX4X1 U6009 ( .A(n5534), .B(n5532), .C(n5533), .D(n5531), .S0(n7940), .S1(
        n7879), .Y(n5535) );
  MX4X1 U6010 ( .A(\registers[408][2] ), .B(\registers[409][2] ), .C(
        \registers[410][2] ), .D(\registers[411][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5532) );
  MX4X1 U6011 ( .A(\registers[412][2] ), .B(\registers[413][2] ), .C(
        \registers[414][2] ), .D(\registers[415][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5531) );
  MX4X1 U6012 ( .A(\registers[400][2] ), .B(\registers[401][2] ), .C(
        \registers[402][2] ), .D(\registers[403][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5534) );
  MX4X1 U6013 ( .A(n5640), .B(n5638), .C(n5639), .D(n5637), .S0(n7941), .S1(
        n7880), .Y(n5641) );
  MX4X1 U6014 ( .A(\registers[88][2] ), .B(\registers[89][2] ), .C(
        \registers[90][2] ), .D(\registers[91][2] ), .S0(n7509), .S1(n7747), 
        .Y(n5638) );
  MX4X1 U6015 ( .A(\registers[92][2] ), .B(\registers[93][2] ), .C(
        \registers[94][2] ), .D(\registers[95][2] ), .S0(n7509), .S1(n7747), 
        .Y(n5637) );
  MX4X1 U6016 ( .A(\registers[80][2] ), .B(\registers[81][2] ), .C(
        \registers[82][2] ), .D(\registers[83][2] ), .S0(n7509), .S1(n7747), 
        .Y(n5640) );
  MX4X1 U6017 ( .A(n5661), .B(n5659), .C(n5660), .D(n5658), .S0(n7942), .S1(
        n7881), .Y(n5662) );
  MX4X1 U6018 ( .A(\registers[24][2] ), .B(\registers[25][2] ), .C(
        \registers[26][2] ), .D(\registers[27][2] ), .S0(n7510), .S1(n7749), 
        .Y(n5659) );
  MX4X1 U6019 ( .A(\registers[28][2] ), .B(\registers[29][2] ), .C(
        \registers[30][2] ), .D(\registers[31][2] ), .S0(n7510), .S1(n7748), 
        .Y(n5658) );
  MX4X1 U6020 ( .A(\registers[16][2] ), .B(\registers[17][2] ), .C(
        \registers[18][2] ), .D(\registers[19][2] ), .S0(n7510), .S1(n7749), 
        .Y(n5661) );
  MX4X1 U6021 ( .A(n5598), .B(n5596), .C(n5597), .D(n5595), .S0(n7941), .S1(
        n7880), .Y(n5599) );
  MX4X1 U6022 ( .A(\registers[216][2] ), .B(\registers[217][2] ), .C(
        \registers[218][2] ), .D(\registers[219][2] ), .S0(n7506), .S1(n7745), 
        .Y(n5596) );
  MX4X1 U6023 ( .A(\registers[220][2] ), .B(\registers[221][2] ), .C(
        \registers[222][2] ), .D(\registers[223][2] ), .S0(n7506), .S1(n7745), 
        .Y(n5595) );
  MX4X1 U6024 ( .A(\registers[208][2] ), .B(\registers[209][2] ), .C(
        \registers[210][2] ), .D(\registers[211][2] ), .S0(n7506), .S1(n7745), 
        .Y(n5598) );
  MX4X1 U6025 ( .A(n5619), .B(n5617), .C(n5618), .D(n5616), .S0(n7941), .S1(
        n7880), .Y(n5620) );
  MX4X1 U6026 ( .A(\registers[152][2] ), .B(\registers[153][2] ), .C(
        \registers[154][2] ), .D(\registers[155][2] ), .S0(n7508), .S1(n7746), 
        .Y(n5617) );
  MX4X1 U6027 ( .A(\registers[156][2] ), .B(\registers[157][2] ), .C(
        \registers[158][2] ), .D(\registers[159][2] ), .S0(n7508), .S1(n7746), 
        .Y(n5616) );
  MX4X1 U6028 ( .A(\registers[144][2] ), .B(\registers[145][2] ), .C(
        \registers[146][2] ), .D(\registers[147][2] ), .S0(n7508), .S1(n7746), 
        .Y(n5619) );
  MX4X1 U6029 ( .A(n5385), .B(n5383), .C(n5384), .D(n5382), .S0(n7937), .S1(
        n7877), .Y(n5386) );
  MX4X1 U6030 ( .A(\registers[856][2] ), .B(\registers[857][2] ), .C(
        \registers[858][2] ), .D(\registers[859][2] ), .S0(n7493), .S1(n7733), 
        .Y(n5383) );
  MX4X1 U6031 ( .A(\registers[860][2] ), .B(\registers[861][2] ), .C(
        \registers[862][2] ), .D(\registers[863][2] ), .S0(n7493), .S1(n7732), 
        .Y(n5382) );
  MX4X1 U6032 ( .A(\registers[848][2] ), .B(\registers[849][2] ), .C(
        \registers[850][2] ), .D(\registers[851][2] ), .S0(n7493), .S1(n7733), 
        .Y(n5385) );
  MX4X1 U6033 ( .A(n5406), .B(n5404), .C(n5405), .D(n5403), .S0(n7938), .S1(
        n7877), .Y(n5407) );
  MX4X1 U6034 ( .A(\registers[792][2] ), .B(\registers[793][2] ), .C(
        \registers[794][2] ), .D(\registers[795][2] ), .S0(n7494), .S1(n7734), 
        .Y(n5404) );
  MX4X1 U6035 ( .A(\registers[796][2] ), .B(\registers[797][2] ), .C(
        \registers[798][2] ), .D(\registers[799][2] ), .S0(n7494), .S1(n7734), 
        .Y(n5403) );
  MX4X1 U6036 ( .A(\registers[784][2] ), .B(\registers[785][2] ), .C(
        \registers[786][2] ), .D(\registers[787][2] ), .S0(n7494), .S1(n7734), 
        .Y(n5406) );
  MX4X1 U6037 ( .A(n5343), .B(n5341), .C(n5342), .D(n5340), .S0(n7937), .S1(
        n7876), .Y(n5344) );
  MX4X1 U6038 ( .A(\registers[984][2] ), .B(\registers[985][2] ), .C(
        \registers[986][2] ), .D(\registers[987][2] ), .S0(n7490), .S1(n7730), 
        .Y(n5341) );
  MX4X1 U6039 ( .A(\registers[988][2] ), .B(\registers[989][2] ), .C(
        \registers[990][2] ), .D(\registers[991][2] ), .S0(n7490), .S1(n7730), 
        .Y(n5340) );
  MX4X1 U6040 ( .A(\registers[976][2] ), .B(\registers[977][2] ), .C(
        \registers[978][2] ), .D(\registers[979][2] ), .S0(n7490), .S1(n7730), 
        .Y(n5343) );
  MX4X1 U6041 ( .A(n5364), .B(n5362), .C(n5363), .D(n5361), .S0(n7937), .S1(
        n7876), .Y(n5365) );
  MX4X1 U6042 ( .A(\registers[920][2] ), .B(\registers[921][2] ), .C(
        \registers[922][2] ), .D(\registers[923][2] ), .S0(n7492), .S1(n7731), 
        .Y(n5362) );
  MX4X1 U6043 ( .A(\registers[924][2] ), .B(\registers[925][2] ), .C(
        \registers[926][2] ), .D(\registers[927][2] ), .S0(n7492), .S1(n7731), 
        .Y(n5361) );
  MX4X1 U6044 ( .A(\registers[912][2] ), .B(\registers[913][2] ), .C(
        \registers[914][2] ), .D(\registers[915][2] ), .S0(n7492), .S1(n7731), 
        .Y(n5364) );
  MX4X1 U6045 ( .A(n5470), .B(n5468), .C(n5469), .D(n5467), .S0(n7939), .S1(
        n7878), .Y(n5471) );
  MX4X1 U6046 ( .A(\registers[600][2] ), .B(\registers[601][2] ), .C(
        \registers[602][2] ), .D(\registers[603][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5468) );
  MX4X1 U6047 ( .A(\registers[604][2] ), .B(\registers[605][2] ), .C(
        \registers[606][2] ), .D(\registers[607][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5467) );
  MX4X1 U6048 ( .A(\registers[592][2] ), .B(\registers[593][2] ), .C(
        \registers[594][2] ), .D(\registers[595][2] ), .S0(n7498), .S1(n7738), 
        .Y(n5470) );
  MX4X1 U6049 ( .A(n5491), .B(n5489), .C(n5490), .D(n5488), .S0(n7939), .S1(
        n7878), .Y(n5492) );
  MX4X1 U6050 ( .A(\registers[536][2] ), .B(\registers[537][2] ), .C(
        \registers[538][2] ), .D(\registers[539][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5489) );
  MX4X1 U6051 ( .A(\registers[540][2] ), .B(\registers[541][2] ), .C(
        \registers[542][2] ), .D(\registers[543][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5488) );
  MX4X1 U6052 ( .A(\registers[528][2] ), .B(\registers[529][2] ), .C(
        \registers[530][2] ), .D(\registers[531][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5491) );
  MX4X1 U6053 ( .A(n5428), .B(n5426), .C(n5427), .D(n5425), .S0(n7938), .S1(
        n7877), .Y(n5429) );
  MX4X1 U6054 ( .A(\registers[728][2] ), .B(\registers[729][2] ), .C(
        \registers[730][2] ), .D(\registers[731][2] ), .S0(n7496), .S1(n7735), 
        .Y(n5426) );
  MX4X1 U6055 ( .A(\registers[732][2] ), .B(\registers[733][2] ), .C(
        \registers[734][2] ), .D(\registers[735][2] ), .S0(n7496), .S1(n7735), 
        .Y(n5425) );
  MX4X1 U6056 ( .A(\registers[720][2] ), .B(\registers[721][2] ), .C(
        \registers[722][2] ), .D(\registers[723][2] ), .S0(n7496), .S1(n7735), 
        .Y(n5428) );
  MX4X1 U6057 ( .A(n5449), .B(n5447), .C(n5448), .D(n5446), .S0(n7938), .S1(
        n7878), .Y(n5450) );
  MX4X1 U6058 ( .A(\registers[664][2] ), .B(\registers[665][2] ), .C(
        \registers[666][2] ), .D(\registers[667][2] ), .S0(n7497), .S1(n7736), 
        .Y(n5447) );
  MX4X1 U6059 ( .A(\registers[668][2] ), .B(\registers[669][2] ), .C(
        \registers[670][2] ), .D(\registers[671][2] ), .S0(n7497), .S1(n7736), 
        .Y(n5446) );
  MX4X1 U6060 ( .A(\registers[656][2] ), .B(\registers[657][2] ), .C(
        \registers[658][2] ), .D(\registers[659][2] ), .S0(n7497), .S1(n7736), 
        .Y(n5449) );
  MX4X1 U6061 ( .A(n5895), .B(n5893), .C(n5894), .D(n5892), .S0(n7945), .S1(
        n7884), .Y(n5896) );
  MX4X1 U6062 ( .A(\registers[344][3] ), .B(\registers[345][3] ), .C(
        \registers[346][3] ), .D(\registers[347][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5893) );
  MX4X1 U6063 ( .A(\registers[348][3] ), .B(\registers[349][3] ), .C(
        \registers[350][3] ), .D(\registers[351][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5892) );
  MX4X1 U6064 ( .A(\registers[336][3] ), .B(\registers[337][3] ), .C(
        \registers[338][3] ), .D(\registers[339][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5895) );
  MX4X1 U6065 ( .A(n5916), .B(n5914), .C(n5915), .D(n5913), .S0(n7946), .S1(
        n7884), .Y(n5917) );
  MX4X1 U6066 ( .A(\registers[280][3] ), .B(\registers[281][3] ), .C(
        \registers[282][3] ), .D(\registers[283][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5914) );
  MX4X1 U6067 ( .A(\registers[284][3] ), .B(\registers[285][3] ), .C(
        \registers[286][3] ), .D(\registers[287][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5913) );
  MX4X1 U6068 ( .A(\registers[272][3] ), .B(\registers[273][3] ), .C(
        \registers[274][3] ), .D(\registers[275][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5916) );
  MX4X1 U6069 ( .A(n5853), .B(n5851), .C(n5852), .D(n5850), .S0(n7945), .S1(
        n7884), .Y(n5854) );
  MX4X1 U6070 ( .A(\registers[472][3] ), .B(\registers[473][3] ), .C(
        \registers[474][3] ), .D(\registers[475][3] ), .S0(n7522), .S1(n7760), 
        .Y(n5851) );
  MX4X1 U6071 ( .A(\registers[476][3] ), .B(\registers[477][3] ), .C(
        \registers[478][3] ), .D(\registers[479][3] ), .S0(n7522), .S1(n7760), 
        .Y(n5850) );
  MX4X1 U6072 ( .A(\registers[464][3] ), .B(\registers[465][3] ), .C(
        \registers[466][3] ), .D(\registers[467][3] ), .S0(n7522), .S1(n7760), 
        .Y(n5853) );
  MX4X1 U6073 ( .A(n5874), .B(n5872), .C(n5873), .D(n5871), .S0(n7945), .S1(
        n7884), .Y(n5875) );
  MX4X1 U6074 ( .A(\registers[408][3] ), .B(\registers[409][3] ), .C(
        \registers[410][3] ), .D(\registers[411][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5872) );
  MX4X1 U6075 ( .A(\registers[412][3] ), .B(\registers[413][3] ), .C(
        \registers[414][3] ), .D(\registers[415][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5871) );
  MX4X1 U6076 ( .A(\registers[400][3] ), .B(\registers[401][3] ), .C(
        \registers[402][3] ), .D(\registers[403][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5874) );
  MX4X1 U6077 ( .A(n5980), .B(n5978), .C(n5979), .D(n5977), .S0(n7947), .S1(
        n7885), .Y(n5981) );
  MX4X1 U6078 ( .A(\registers[88][3] ), .B(\registers[89][3] ), .C(
        \registers[90][3] ), .D(\registers[91][3] ), .S0(n7530), .S1(n7767), 
        .Y(n5978) );
  MX4X1 U6079 ( .A(\registers[92][3] ), .B(\registers[93][3] ), .C(
        \registers[94][3] ), .D(\registers[95][3] ), .S0(n7530), .S1(n7767), 
        .Y(n5977) );
  MX4X1 U6080 ( .A(\registers[80][3] ), .B(\registers[81][3] ), .C(
        \registers[82][3] ), .D(\registers[83][3] ), .S0(n7530), .S1(n7767), 
        .Y(n5980) );
  MX4X1 U6081 ( .A(n6001), .B(n5999), .C(n6000), .D(n5998), .S0(n7947), .S1(
        n7886), .Y(n6002) );
  MX4X1 U6082 ( .A(\registers[24][3] ), .B(\registers[25][3] ), .C(
        \registers[26][3] ), .D(\registers[27][3] ), .S0(n7532), .S1(n7768), 
        .Y(n5999) );
  MX4X1 U6083 ( .A(\registers[28][3] ), .B(\registers[29][3] ), .C(
        \registers[30][3] ), .D(\registers[31][3] ), .S0(n7532), .S1(n7768), 
        .Y(n5998) );
  MX4X1 U6084 ( .A(\registers[16][3] ), .B(\registers[17][3] ), .C(
        \registers[18][3] ), .D(\registers[19][3] ), .S0(n7532), .S1(n7768), 
        .Y(n6001) );
  MX4X1 U6085 ( .A(n5938), .B(n5936), .C(n5937), .D(n5935), .S0(n7946), .S1(
        n7885), .Y(n5939) );
  MX4X1 U6086 ( .A(\registers[216][3] ), .B(\registers[217][3] ), .C(
        \registers[218][3] ), .D(\registers[219][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5936) );
  MX4X1 U6087 ( .A(\registers[220][3] ), .B(\registers[221][3] ), .C(
        \registers[222][3] ), .D(\registers[223][3] ), .S0(n7528), .S1(n7764), 
        .Y(n5935) );
  MX4X1 U6088 ( .A(\registers[208][3] ), .B(\registers[209][3] ), .C(
        \registers[210][3] ), .D(\registers[211][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5938) );
  MX4X1 U6089 ( .A(n5959), .B(n5957), .C(n5958), .D(n5956), .S0(n7946), .S1(
        n7885), .Y(n5960) );
  MX4X1 U6090 ( .A(\registers[152][3] ), .B(\registers[153][3] ), .C(
        \registers[154][3] ), .D(\registers[155][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5957) );
  MX4X1 U6091 ( .A(\registers[156][3] ), .B(\registers[157][3] ), .C(
        \registers[158][3] ), .D(\registers[159][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5956) );
  MX4X1 U6092 ( .A(\registers[144][3] ), .B(\registers[145][3] ), .C(
        \registers[146][3] ), .D(\registers[147][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5959) );
  MX4X1 U6093 ( .A(n5725), .B(n5723), .C(n5724), .D(n5722), .S0(n7943), .S1(
        n7882), .Y(n5726) );
  MX4X1 U6094 ( .A(\registers[856][3] ), .B(\registers[857][3] ), .C(
        \registers[858][3] ), .D(\registers[859][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5723) );
  MX4X1 U6095 ( .A(\registers[860][3] ), .B(\registers[861][3] ), .C(
        \registers[862][3] ), .D(\registers[863][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5722) );
  MX4X1 U6096 ( .A(\registers[848][3] ), .B(\registers[849][3] ), .C(
        \registers[850][3] ), .D(\registers[851][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5725) );
  MX4X1 U6097 ( .A(n5746), .B(n5744), .C(n5745), .D(n5743), .S0(n7943), .S1(
        n7882), .Y(n5747) );
  MX4X1 U6098 ( .A(\registers[792][3] ), .B(\registers[793][3] ), .C(
        \registers[794][3] ), .D(\registers[795][3] ), .S0(n7516), .S1(n7753), 
        .Y(n5744) );
  MX4X1 U6099 ( .A(\registers[796][3] ), .B(\registers[797][3] ), .C(
        \registers[798][3] ), .D(\registers[799][3] ), .S0(n7516), .S1(n7753), 
        .Y(n5743) );
  MX4X1 U6100 ( .A(\registers[784][3] ), .B(\registers[785][3] ), .C(
        \registers[786][3] ), .D(\registers[787][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5746) );
  MX4X1 U6101 ( .A(n5683), .B(n5681), .C(n5682), .D(n5680), .S0(n7942), .S1(
        n7881), .Y(n5684) );
  MX4X1 U6102 ( .A(\registers[984][3] ), .B(\registers[985][3] ), .C(
        \registers[986][3] ), .D(\registers[987][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5681) );
  MX4X1 U6103 ( .A(\registers[988][3] ), .B(\registers[989][3] ), .C(
        \registers[990][3] ), .D(\registers[991][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5680) );
  MX4X1 U6104 ( .A(\registers[976][3] ), .B(\registers[977][3] ), .C(
        \registers[978][3] ), .D(\registers[979][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5683) );
  MX4X1 U6105 ( .A(n5704), .B(n5702), .C(n5703), .D(n5701), .S0(n7942), .S1(
        n7881), .Y(n5705) );
  MX4X1 U6106 ( .A(\registers[920][3] ), .B(\registers[921][3] ), .C(
        \registers[922][3] ), .D(\registers[923][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5702) );
  MX4X1 U6107 ( .A(\registers[924][3] ), .B(\registers[925][3] ), .C(
        \registers[926][3] ), .D(\registers[927][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5701) );
  MX4X1 U6108 ( .A(\registers[912][3] ), .B(\registers[913][3] ), .C(
        \registers[914][3] ), .D(\registers[915][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5704) );
  MX4X1 U6109 ( .A(n5810), .B(n5808), .C(n5809), .D(n5807), .S0(n7944), .S1(
        n7883), .Y(n5811) );
  MX4X1 U6110 ( .A(\registers[600][3] ), .B(\registers[601][3] ), .C(
        \registers[602][3] ), .D(\registers[603][3] ), .S0(n7520), .S1(n7757), 
        .Y(n5808) );
  MX4X1 U6111 ( .A(\registers[604][3] ), .B(\registers[605][3] ), .C(
        \registers[606][3] ), .D(\registers[607][3] ), .S0(n7520), .S1(n7757), 
        .Y(n5807) );
  MX4X1 U6112 ( .A(\registers[592][3] ), .B(\registers[593][3] ), .C(
        \registers[594][3] ), .D(\registers[595][3] ), .S0(n7520), .S1(n7757), 
        .Y(n5810) );
  MX4X1 U6113 ( .A(n5831), .B(n5829), .C(n5830), .D(n5828), .S0(n7944), .S1(
        n7883), .Y(n5832) );
  MX4X1 U6114 ( .A(\registers[536][3] ), .B(\registers[537][3] ), .C(
        \registers[538][3] ), .D(\registers[539][3] ), .S0(n7521), .S1(n7758), 
        .Y(n5829) );
  MX4X1 U6115 ( .A(\registers[540][3] ), .B(\registers[541][3] ), .C(
        \registers[542][3] ), .D(\registers[543][3] ), .S0(n7521), .S1(n7758), 
        .Y(n5828) );
  MX4X1 U6116 ( .A(\registers[528][3] ), .B(\registers[529][3] ), .C(
        \registers[530][3] ), .D(\registers[531][3] ), .S0(n7521), .S1(n7759), 
        .Y(n5831) );
  MX4X1 U6117 ( .A(n5768), .B(n5766), .C(n5767), .D(n5765), .S0(n7943), .S1(
        n7882), .Y(n5769) );
  MX4X1 U6118 ( .A(\registers[728][3] ), .B(\registers[729][3] ), .C(
        \registers[730][3] ), .D(\registers[731][3] ), .S0(n7517), .S1(n7755), 
        .Y(n5766) );
  MX4X1 U6119 ( .A(\registers[732][3] ), .B(\registers[733][3] ), .C(
        \registers[734][3] ), .D(\registers[735][3] ), .S0(n7517), .S1(n7755), 
        .Y(n5765) );
  MX4X1 U6120 ( .A(\registers[720][3] ), .B(\registers[721][3] ), .C(
        \registers[722][3] ), .D(\registers[723][3] ), .S0(n7517), .S1(n7755), 
        .Y(n5768) );
  MX4X1 U6121 ( .A(n5789), .B(n5787), .C(n5788), .D(n5786), .S0(n7944), .S1(
        n7883), .Y(n5790) );
  MX4X1 U6122 ( .A(\registers[664][3] ), .B(\registers[665][3] ), .C(
        \registers[666][3] ), .D(\registers[667][3] ), .S0(n7518), .S1(n7756), 
        .Y(n5787) );
  MX4X1 U6123 ( .A(\registers[668][3] ), .B(\registers[669][3] ), .C(
        \registers[670][3] ), .D(\registers[671][3] ), .S0(n7518), .S1(n7756), 
        .Y(n5786) );
  MX4X1 U6124 ( .A(\registers[656][3] ), .B(\registers[657][3] ), .C(
        \registers[658][3] ), .D(\registers[659][3] ), .S0(n7518), .S1(n7756), 
        .Y(n5789) );
  MX4X1 U6125 ( .A(n6235), .B(n6233), .C(n6234), .D(n6232), .S0(n7951), .S1(
        n7889), .Y(n6236) );
  MX4X1 U6126 ( .A(\registers[344][4] ), .B(\registers[345][4] ), .C(
        \registers[346][4] ), .D(\registers[347][4] ), .S0(n7546), .S1(n7782), 
        .Y(n6233) );
  MX4X1 U6127 ( .A(\registers[348][4] ), .B(\registers[349][4] ), .C(
        \registers[350][4] ), .D(\registers[351][4] ), .S0(n7546), .S1(n7782), 
        .Y(n6232) );
  MX4X1 U6128 ( .A(\registers[336][4] ), .B(\registers[337][4] ), .C(
        \registers[338][4] ), .D(\registers[339][4] ), .S0(n7546), .S1(n7782), 
        .Y(n6235) );
  MX4X1 U6129 ( .A(n6256), .B(n6254), .C(n6255), .D(n6253), .S0(n7951), .S1(
        n7889), .Y(n6257) );
  MX4X1 U6130 ( .A(\registers[280][4] ), .B(\registers[281][4] ), .C(
        \registers[282][4] ), .D(\registers[283][4] ), .S0(n7548), .S1(n7783), 
        .Y(n6254) );
  MX4X1 U6131 ( .A(\registers[284][4] ), .B(\registers[285][4] ), .C(
        \registers[286][4] ), .D(\registers[287][4] ), .S0(n7548), .S1(n7783), 
        .Y(n6253) );
  MX4X1 U6132 ( .A(\registers[272][4] ), .B(\registers[273][4] ), .C(
        \registers[274][4] ), .D(\registers[275][4] ), .S0(n7548), .S1(n7783), 
        .Y(n6256) );
  MX4X1 U6133 ( .A(n6193), .B(n6191), .C(n6192), .D(n6190), .S0(n7950), .S1(
        n7888), .Y(n6194) );
  MX4X1 U6134 ( .A(\registers[472][4] ), .B(\registers[473][4] ), .C(
        \registers[474][4] ), .D(\registers[475][4] ), .S0(n7544), .S1(n7779), 
        .Y(n6191) );
  MX4X1 U6135 ( .A(\registers[476][4] ), .B(\registers[477][4] ), .C(
        \registers[478][4] ), .D(\registers[479][4] ), .S0(n7544), .S1(n7779), 
        .Y(n6190) );
  MX4X1 U6136 ( .A(\registers[464][4] ), .B(\registers[465][4] ), .C(
        \registers[466][4] ), .D(\registers[467][4] ), .S0(n7544), .S1(n7779), 
        .Y(n6193) );
  MX4X1 U6137 ( .A(n6214), .B(n6212), .C(n6213), .D(n6211), .S0(n7950), .S1(
        n7889), .Y(n6215) );
  MX4X1 U6138 ( .A(\registers[408][4] ), .B(\registers[409][4] ), .C(
        \registers[410][4] ), .D(\registers[411][4] ), .S0(n7545), .S1(n7781), 
        .Y(n6212) );
  MX4X1 U6139 ( .A(\registers[412][4] ), .B(\registers[413][4] ), .C(
        \registers[414][4] ), .D(\registers[415][4] ), .S0(n7545), .S1(n7780), 
        .Y(n6211) );
  MX4X1 U6140 ( .A(\registers[400][4] ), .B(\registers[401][4] ), .C(
        \registers[402][4] ), .D(\registers[403][4] ), .S0(n7545), .S1(n7781), 
        .Y(n6214) );
  MX4X1 U6141 ( .A(n6320), .B(n6318), .C(n6319), .D(n6317), .S0(n7952), .S1(
        n7890), .Y(n6321) );
  MX4X1 U6142 ( .A(\registers[88][4] ), .B(\registers[89][4] ), .C(
        \registers[90][4] ), .D(\registers[91][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6318) );
  MX4X1 U6143 ( .A(\registers[92][4] ), .B(\registers[93][4] ), .C(
        \registers[94][4] ), .D(\registers[95][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6317) );
  MX4X1 U6144 ( .A(\registers[80][4] ), .B(\registers[81][4] ), .C(
        \registers[82][4] ), .D(\registers[83][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6320) );
  MX4X1 U6145 ( .A(n6341), .B(n6339), .C(n6340), .D(n6338), .S0(n7952), .S1(
        n7891), .Y(n6342) );
  MX4X1 U6146 ( .A(\registers[24][4] ), .B(\registers[25][4] ), .C(
        \registers[26][4] ), .D(\registers[27][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6339) );
  MX4X1 U6147 ( .A(\registers[28][4] ), .B(\registers[29][4] ), .C(
        \registers[30][4] ), .D(\registers[31][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6338) );
  MX4X1 U6148 ( .A(\registers[16][4] ), .B(\registers[17][4] ), .C(
        \registers[18][4] ), .D(\registers[19][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6341) );
  MX4X1 U6149 ( .A(n6278), .B(n6276), .C(n6277), .D(n6275), .S0(n7951), .S1(
        n7890), .Y(n6279) );
  MX4X1 U6150 ( .A(\registers[216][4] ), .B(\registers[217][4] ), .C(
        \registers[218][4] ), .D(\registers[219][4] ), .S0(n7549), .S1(n7784), 
        .Y(n6276) );
  MX4X1 U6151 ( .A(\registers[220][4] ), .B(\registers[221][4] ), .C(
        \registers[222][4] ), .D(\registers[223][4] ), .S0(n7549), .S1(n7784), 
        .Y(n6275) );
  MX4X1 U6152 ( .A(\registers[208][4] ), .B(\registers[209][4] ), .C(
        \registers[210][4] ), .D(\registers[211][4] ), .S0(n7549), .S1(n7784), 
        .Y(n6278) );
  MX4X1 U6153 ( .A(n6299), .B(n6297), .C(n6298), .D(n6296), .S0(n7952), .S1(
        n7890), .Y(n6300) );
  MX4X1 U6154 ( .A(\registers[152][4] ), .B(\registers[153][4] ), .C(
        \registers[154][4] ), .D(\registers[155][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6297) );
  MX4X1 U6155 ( .A(\registers[156][4] ), .B(\registers[157][4] ), .C(
        \registers[158][4] ), .D(\registers[159][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6296) );
  MX4X1 U6156 ( .A(\registers[144][4] ), .B(\registers[145][4] ), .C(
        \registers[146][4] ), .D(\registers[147][4] ), .S0(n7550), .S1(n7786), 
        .Y(n6299) );
  MX4X1 U6157 ( .A(n6065), .B(n6063), .C(n6064), .D(n6062), .S0(n7948), .S1(
        n7887), .Y(n6066) );
  MX4X1 U6158 ( .A(\registers[856][4] ), .B(\registers[857][4] ), .C(
        \registers[858][4] ), .D(\registers[859][4] ), .S0(n7536), .S1(n7772), 
        .Y(n6063) );
  MX4X1 U6159 ( .A(\registers[860][4] ), .B(\registers[861][4] ), .C(
        \registers[862][4] ), .D(\registers[863][4] ), .S0(n7536), .S1(n7772), 
        .Y(n6062) );
  MX4X1 U6160 ( .A(\registers[848][4] ), .B(\registers[849][4] ), .C(
        \registers[850][4] ), .D(\registers[851][4] ), .S0(n7536), .S1(n7772), 
        .Y(n6065) );
  MX4X1 U6161 ( .A(n6086), .B(n6084), .C(n6085), .D(n6083), .S0(n7948), .S1(
        n7887), .Y(n6087) );
  MX4X1 U6162 ( .A(\registers[792][4] ), .B(\registers[793][4] ), .C(
        \registers[794][4] ), .D(\registers[795][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6084) );
  MX4X1 U6163 ( .A(\registers[796][4] ), .B(\registers[797][4] ), .C(
        \registers[798][4] ), .D(\registers[799][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6083) );
  MX4X1 U6164 ( .A(\registers[784][4] ), .B(\registers[785][4] ), .C(
        \registers[786][4] ), .D(\registers[787][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6086) );
  MX4X1 U6165 ( .A(n6023), .B(n6021), .C(n6022), .D(n6020), .S0(n7947), .S1(
        n7886), .Y(n6024) );
  MX4X1 U6166 ( .A(\registers[984][4] ), .B(\registers[985][4] ), .C(
        \registers[986][4] ), .D(\registers[987][4] ), .S0(n7533), .S1(n7769), 
        .Y(n6021) );
  MX4X1 U6167 ( .A(\registers[988][4] ), .B(\registers[989][4] ), .C(
        \registers[990][4] ), .D(\registers[991][4] ), .S0(n7533), .S1(n7769), 
        .Y(n6020) );
  MX4X1 U6168 ( .A(\registers[976][4] ), .B(\registers[977][4] ), .C(
        \registers[978][4] ), .D(\registers[979][4] ), .S0(n7533), .S1(n7770), 
        .Y(n6023) );
  MX4X1 U6169 ( .A(n6044), .B(n6042), .C(n6043), .D(n6041), .S0(n7948), .S1(
        n7886), .Y(n6045) );
  MX4X1 U6170 ( .A(\registers[920][4] ), .B(\registers[921][4] ), .C(
        \registers[922][4] ), .D(\registers[923][4] ), .S0(n7534), .S1(n7771), 
        .Y(n6042) );
  MX4X1 U6171 ( .A(\registers[924][4] ), .B(\registers[925][4] ), .C(
        \registers[926][4] ), .D(\registers[927][4] ), .S0(n7534), .S1(n7771), 
        .Y(n6041) );
  MX4X1 U6172 ( .A(\registers[912][4] ), .B(\registers[913][4] ), .C(
        \registers[914][4] ), .D(\registers[915][4] ), .S0(n7534), .S1(n7771), 
        .Y(n6044) );
  MX4X1 U6173 ( .A(n6150), .B(n6148), .C(n6149), .D(n6147), .S0(n7949), .S1(
        n7888), .Y(n6151) );
  MX4X1 U6174 ( .A(\registers[600][4] ), .B(\registers[601][4] ), .C(
        \registers[602][4] ), .D(\registers[603][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6148) );
  MX4X1 U6175 ( .A(\registers[604][4] ), .B(\registers[605][4] ), .C(
        \registers[606][4] ), .D(\registers[607][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6147) );
  MX4X1 U6176 ( .A(\registers[592][4] ), .B(\registers[593][4] ), .C(
        \registers[594][4] ), .D(\registers[595][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6150) );
  MX4X1 U6177 ( .A(n6171), .B(n6169), .C(n6170), .D(n6168), .S0(n7950), .S1(
        n7888), .Y(n6172) );
  MX4X1 U6178 ( .A(\registers[536][4] ), .B(\registers[537][4] ), .C(
        \registers[538][4] ), .D(\registers[539][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6169) );
  MX4X1 U6179 ( .A(\registers[540][4] ), .B(\registers[541][4] ), .C(
        \registers[542][4] ), .D(\registers[543][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6168) );
  MX4X1 U6180 ( .A(\registers[528][4] ), .B(\registers[529][4] ), .C(
        \registers[530][4] ), .D(\registers[531][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6171) );
  MX4X1 U6181 ( .A(n6108), .B(n6106), .C(n6107), .D(n6105), .S0(n7949), .S1(
        n7887), .Y(n6109) );
  MX4X1 U6182 ( .A(\registers[728][4] ), .B(\registers[729][4] ), .C(
        \registers[730][4] ), .D(\registers[731][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6106) );
  MX4X1 U6183 ( .A(\registers[732][4] ), .B(\registers[733][4] ), .C(
        \registers[734][4] ), .D(\registers[735][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6105) );
  MX4X1 U6184 ( .A(\registers[720][4] ), .B(\registers[721][4] ), .C(
        \registers[722][4] ), .D(\registers[723][4] ), .S0(n7538), .S1(n7775), 
        .Y(n6108) );
  MX4X1 U6185 ( .A(n6129), .B(n6127), .C(n6128), .D(n6126), .S0(n7949), .S1(
        n7888), .Y(n6130) );
  MX4X1 U6186 ( .A(\registers[664][4] ), .B(\registers[665][4] ), .C(
        \registers[666][4] ), .D(\registers[667][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6127) );
  MX4X1 U6187 ( .A(\registers[668][4] ), .B(\registers[669][4] ), .C(
        \registers[670][4] ), .D(\registers[671][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6126) );
  MX4X1 U6188 ( .A(\registers[656][4] ), .B(\registers[657][4] ), .C(
        \registers[658][4] ), .D(\registers[659][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6129) );
  MX4X1 U6189 ( .A(n6575), .B(n6573), .C(n6574), .D(n6572), .S0(n7956), .S1(
        n7894), .Y(n6576) );
  MX4X1 U6190 ( .A(\registers[344][5] ), .B(\registers[345][5] ), .C(
        \registers[346][5] ), .D(\registers[347][5] ), .S0(n7568), .S1(n7801), 
        .Y(n6573) );
  MX4X1 U6191 ( .A(\registers[348][5] ), .B(\registers[349][5] ), .C(
        \registers[350][5] ), .D(\registers[351][5] ), .S0(n7568), .S1(n7801), 
        .Y(n6572) );
  MX4X1 U6192 ( .A(\registers[336][5] ), .B(\registers[337][5] ), .C(
        \registers[338][5] ), .D(\registers[339][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6575) );
  MX4X1 U6193 ( .A(n6596), .B(n6594), .C(n6595), .D(n6593), .S0(n7956), .S1(
        n7894), .Y(n6597) );
  MX4X1 U6194 ( .A(\registers[280][5] ), .B(\registers[281][5] ), .C(
        \registers[282][5] ), .D(\registers[283][5] ), .S0(n7569), .S1(n7803), 
        .Y(n6594) );
  MX4X1 U6195 ( .A(\registers[284][5] ), .B(\registers[285][5] ), .C(
        \registers[286][5] ), .D(\registers[287][5] ), .S0(n7569), .S1(n7803), 
        .Y(n6593) );
  MX4X1 U6196 ( .A(\registers[272][5] ), .B(\registers[273][5] ), .C(
        \registers[274][5] ), .D(\registers[275][5] ), .S0(n7569), .S1(n7803), 
        .Y(n6596) );
  MX4X1 U6197 ( .A(n6533), .B(n6531), .C(n6532), .D(n6530), .S0(n7955), .S1(
        n7893), .Y(n6534) );
  MX4X1 U6198 ( .A(\registers[472][5] ), .B(\registers[473][5] ), .C(
        \registers[474][5] ), .D(\registers[475][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6531) );
  MX4X1 U6199 ( .A(\registers[476][5] ), .B(\registers[477][5] ), .C(
        \registers[478][5] ), .D(\registers[479][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6530) );
  MX4X1 U6200 ( .A(\registers[464][5] ), .B(\registers[465][5] ), .C(
        \registers[466][5] ), .D(\registers[467][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6533) );
  MX4X1 U6201 ( .A(n6554), .B(n6552), .C(n6553), .D(n6551), .S0(n7956), .S1(
        n7894), .Y(n6555) );
  MX4X1 U6202 ( .A(\registers[408][5] ), .B(\registers[409][5] ), .C(
        \registers[410][5] ), .D(\registers[411][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6552) );
  MX4X1 U6203 ( .A(\registers[412][5] ), .B(\registers[413][5] ), .C(
        \registers[414][5] ), .D(\registers[415][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6551) );
  MX4X1 U6204 ( .A(\registers[400][5] ), .B(\registers[401][5] ), .C(
        \registers[402][5] ), .D(\registers[403][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6554) );
  MX4X1 U6205 ( .A(n6660), .B(n6658), .C(n6659), .D(n6657), .S0(n7957), .S1(
        n7895), .Y(n6661) );
  MX4X1 U6206 ( .A(\registers[88][5] ), .B(\registers[89][5] ), .C(
        \registers[90][5] ), .D(\registers[91][5] ), .S0(n7573), .S1(n7805), 
        .Y(n6658) );
  MX4X1 U6207 ( .A(\registers[92][5] ), .B(\registers[93][5] ), .C(
        \registers[94][5] ), .D(\registers[95][5] ), .S0(n7573), .S1(n7805), 
        .Y(n6657) );
  MX4X1 U6208 ( .A(\registers[80][5] ), .B(\registers[81][5] ), .C(
        \registers[82][5] ), .D(\registers[83][5] ), .S0(n7573), .S1(n7806), 
        .Y(n6660) );
  MX4X1 U6209 ( .A(n6681), .B(n6679), .C(n6680), .D(n6678), .S0(n7958), .S1(
        n7896), .Y(n6682) );
  MX4X1 U6210 ( .A(\registers[24][5] ), .B(\registers[25][5] ), .C(
        \registers[26][5] ), .D(\registers[27][5] ), .S0(n7574), .S1(n7807), 
        .Y(n6679) );
  MX4X1 U6211 ( .A(\registers[28][5] ), .B(\registers[29][5] ), .C(
        \registers[30][5] ), .D(\registers[31][5] ), .S0(n7574), .S1(n7807), 
        .Y(n6678) );
  MX4X1 U6212 ( .A(\registers[16][5] ), .B(\registers[17][5] ), .C(
        \registers[18][5] ), .D(\registers[19][5] ), .S0(n7574), .S1(n7807), 
        .Y(n6681) );
  MX4X1 U6213 ( .A(n6618), .B(n6616), .C(n6617), .D(n6615), .S0(n7957), .S1(
        n7895), .Y(n6619) );
  MX4X1 U6214 ( .A(\registers[216][5] ), .B(\registers[217][5] ), .C(
        \registers[218][5] ), .D(\registers[219][5] ), .S0(n7570), .S1(n7818), 
        .Y(n6616) );
  MX4X1 U6215 ( .A(\registers[220][5] ), .B(\registers[221][5] ), .C(
        \registers[222][5] ), .D(\registers[223][5] ), .S0(n7570), .S1(n7702), 
        .Y(n6615) );
  MX4X1 U6216 ( .A(\registers[208][5] ), .B(\registers[209][5] ), .C(
        \registers[210][5] ), .D(\registers[211][5] ), .S0(n7570), .S1(n7697), 
        .Y(n6618) );
  MX4X1 U6217 ( .A(n6639), .B(n6637), .C(n6638), .D(n6636), .S0(n7957), .S1(
        n7895), .Y(n6640) );
  MX4X1 U6218 ( .A(\registers[152][5] ), .B(\registers[153][5] ), .C(
        \registers[154][5] ), .D(\registers[155][5] ), .S0(n7572), .S1(n7804), 
        .Y(n6637) );
  MX4X1 U6219 ( .A(\registers[156][5] ), .B(\registers[157][5] ), .C(
        \registers[158][5] ), .D(\registers[159][5] ), .S0(n7572), .S1(n7804), 
        .Y(n6636) );
  MX4X1 U6220 ( .A(\registers[144][5] ), .B(\registers[145][5] ), .C(
        \registers[146][5] ), .D(\registers[147][5] ), .S0(n7572), .S1(n7804), 
        .Y(n6639) );
  MX4X1 U6221 ( .A(n6405), .B(n6403), .C(n6404), .D(n6402), .S0(n7953), .S1(
        n7892), .Y(n6406) );
  MX4X1 U6222 ( .A(\registers[856][5] ), .B(\registers[857][5] ), .C(
        \registers[858][5] ), .D(\registers[859][5] ), .S0(n7557), .S1(n7792), 
        .Y(n6403) );
  MX4X1 U6223 ( .A(\registers[860][5] ), .B(\registers[861][5] ), .C(
        \registers[862][5] ), .D(\registers[863][5] ), .S0(n7557), .S1(n7792), 
        .Y(n6402) );
  MX4X1 U6224 ( .A(\registers[848][5] ), .B(\registers[849][5] ), .C(
        \registers[850][5] ), .D(\registers[851][5] ), .S0(n7557), .S1(n7792), 
        .Y(n6405) );
  MX4X1 U6225 ( .A(n6426), .B(n6424), .C(n6425), .D(n6423), .S0(n7954), .S1(
        n7892), .Y(n6427) );
  MX4X1 U6226 ( .A(\registers[792][5] ), .B(\registers[793][5] ), .C(
        \registers[794][5] ), .D(\registers[795][5] ), .S0(n7558), .S1(n7793), 
        .Y(n6424) );
  MX4X1 U6227 ( .A(\registers[796][5] ), .B(\registers[797][5] ), .C(
        \registers[798][5] ), .D(\registers[799][5] ), .S0(n7558), .S1(n7793), 
        .Y(n6423) );
  MX4X1 U6228 ( .A(\registers[784][5] ), .B(\registers[785][5] ), .C(
        \registers[786][5] ), .D(\registers[787][5] ), .S0(n7558), .S1(n7793), 
        .Y(n6426) );
  MX4X1 U6229 ( .A(n6363), .B(n6361), .C(n6362), .D(n6360), .S0(n7953), .S1(
        n7891), .Y(n6364) );
  MX4X1 U6230 ( .A(\registers[984][5] ), .B(\registers[985][5] ), .C(
        \registers[986][5] ), .D(\registers[987][5] ), .S0(n7554), .S1(n7789), 
        .Y(n6361) );
  MX4X1 U6231 ( .A(\registers[988][5] ), .B(\registers[989][5] ), .C(
        \registers[990][5] ), .D(\registers[991][5] ), .S0(n7554), .S1(n7789), 
        .Y(n6360) );
  MX4X1 U6232 ( .A(\registers[976][5] ), .B(\registers[977][5] ), .C(
        \registers[978][5] ), .D(\registers[979][5] ), .S0(n7554), .S1(n7789), 
        .Y(n6363) );
  MX4X1 U6233 ( .A(n6384), .B(n6382), .C(n6383), .D(n6381), .S0(n7953), .S1(
        n7891), .Y(n6385) );
  MX4X1 U6234 ( .A(\registers[920][5] ), .B(\registers[921][5] ), .C(
        \registers[922][5] ), .D(\registers[923][5] ), .S0(n7556), .S1(n7790), 
        .Y(n6382) );
  MX4X1 U6235 ( .A(\registers[924][5] ), .B(\registers[925][5] ), .C(
        \registers[926][5] ), .D(\registers[927][5] ), .S0(n7556), .S1(n7790), 
        .Y(n6381) );
  MX4X1 U6236 ( .A(\registers[912][5] ), .B(\registers[913][5] ), .C(
        \registers[914][5] ), .D(\registers[915][5] ), .S0(n7556), .S1(n7791), 
        .Y(n6384) );
  MX4X1 U6237 ( .A(n6490), .B(n6488), .C(n6489), .D(n6487), .S0(n7955), .S1(
        n7893), .Y(n6491) );
  MX4X1 U6238 ( .A(\registers[600][5] ), .B(\registers[601][5] ), .C(
        \registers[602][5] ), .D(\registers[603][5] ), .S0(n7562), .S1(n7797), 
        .Y(n6488) );
  MX4X1 U6239 ( .A(\registers[604][5] ), .B(\registers[605][5] ), .C(
        \registers[606][5] ), .D(\registers[607][5] ), .S0(n7562), .S1(n7796), 
        .Y(n6487) );
  MX4X1 U6240 ( .A(\registers[592][5] ), .B(\registers[593][5] ), .C(
        \registers[594][5] ), .D(\registers[595][5] ), .S0(n7562), .S1(n7797), 
        .Y(n6490) );
  MX4X1 U6241 ( .A(n6511), .B(n6509), .C(n6510), .D(n6508), .S0(n7955), .S1(
        n7893), .Y(n6512) );
  MX4X1 U6242 ( .A(\registers[536][5] ), .B(\registers[537][5] ), .C(
        \registers[538][5] ), .D(\registers[539][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6509) );
  MX4X1 U6243 ( .A(\registers[540][5] ), .B(\registers[541][5] ), .C(
        \registers[542][5] ), .D(\registers[543][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6508) );
  MX4X1 U6244 ( .A(\registers[528][5] ), .B(\registers[529][5] ), .C(
        \registers[530][5] ), .D(\registers[531][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6511) );
  MX4X1 U6245 ( .A(n6448), .B(n6446), .C(n6447), .D(n6445), .S0(n7954), .S1(
        n7892), .Y(n6449) );
  MX4X1 U6246 ( .A(\registers[728][5] ), .B(\registers[729][5] ), .C(
        \registers[730][5] ), .D(\registers[731][5] ), .S0(n7560), .S1(n7794), 
        .Y(n6446) );
  MX4X1 U6247 ( .A(\registers[732][5] ), .B(\registers[733][5] ), .C(
        \registers[734][5] ), .D(\registers[735][5] ), .S0(n7560), .S1(n7794), 
        .Y(n6445) );
  MX4X1 U6248 ( .A(\registers[720][5] ), .B(\registers[721][5] ), .C(
        \registers[722][5] ), .D(\registers[723][5] ), .S0(n7560), .S1(n7794), 
        .Y(n6448) );
  MX4X1 U6249 ( .A(n6469), .B(n6467), .C(n6468), .D(n6466), .S0(n7954), .S1(
        n7892), .Y(n6470) );
  MX4X1 U6250 ( .A(\registers[664][5] ), .B(\registers[665][5] ), .C(
        \registers[666][5] ), .D(\registers[667][5] ), .S0(n7561), .S1(n7795), 
        .Y(n6467) );
  MX4X1 U6251 ( .A(\registers[668][5] ), .B(\registers[669][5] ), .C(
        \registers[670][5] ), .D(\registers[671][5] ), .S0(n7561), .S1(n7795), 
        .Y(n6466) );
  MX4X1 U6252 ( .A(\registers[656][5] ), .B(\registers[657][5] ), .C(
        \registers[658][5] ), .D(\registers[659][5] ), .S0(n7561), .S1(n7795), 
        .Y(n6469) );
  MX4X1 U6253 ( .A(n6915), .B(n6913), .C(n6914), .D(n6912), .S0(n7961), .S1(
        n7897), .Y(n6916) );
  MX4X1 U6254 ( .A(\registers[344][6] ), .B(\registers[345][6] ), .C(
        \registers[346][6] ), .D(\registers[347][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6913) );
  MX4X1 U6255 ( .A(\registers[348][6] ), .B(\registers[349][6] ), .C(
        \registers[350][6] ), .D(\registers[351][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6912) );
  MX4X1 U6256 ( .A(\registers[336][6] ), .B(\registers[337][6] ), .C(
        \registers[338][6] ), .D(\registers[339][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6915) );
  MX4X1 U6257 ( .A(n6936), .B(n6934), .C(n6935), .D(n6933), .S0(n7962), .S1(
        n7897), .Y(n6937) );
  MX4X1 U6258 ( .A(\registers[280][6] ), .B(\registers[281][6] ), .C(
        \registers[282][6] ), .D(\registers[283][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6934) );
  MX4X1 U6259 ( .A(\registers[284][6] ), .B(\registers[285][6] ), .C(
        \registers[286][6] ), .D(\registers[287][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6933) );
  MX4X1 U6260 ( .A(\registers[272][6] ), .B(\registers[273][6] ), .C(
        \registers[274][6] ), .D(\registers[275][6] ), .S0(n7590), .S1(n7822), 
        .Y(n6936) );
  MX4X1 U6261 ( .A(n6873), .B(n6871), .C(n6872), .D(n6870), .S0(n7961), .S1(
        n7899), .Y(n6874) );
  MX4X1 U6262 ( .A(\registers[472][6] ), .B(\registers[473][6] ), .C(
        \registers[474][6] ), .D(\registers[475][6] ), .S0(n7586), .S1(n7818), 
        .Y(n6871) );
  MX4X1 U6263 ( .A(\registers[476][6] ), .B(\registers[477][6] ), .C(
        \registers[478][6] ), .D(\registers[479][6] ), .S0(n7586), .S1(n7818), 
        .Y(n6870) );
  MX4X1 U6264 ( .A(\registers[464][6] ), .B(\registers[465][6] ), .C(
        \registers[466][6] ), .D(\registers[467][6] ), .S0(n7586), .S1(n7818), 
        .Y(n6873) );
  MX4X1 U6265 ( .A(n6894), .B(n6892), .C(n6893), .D(n6891), .S0(n7961), .S1(
        n7897), .Y(n6895) );
  MX4X1 U6266 ( .A(\registers[408][6] ), .B(\registers[409][6] ), .C(
        \registers[410][6] ), .D(\registers[411][6] ), .S0(n7588), .S1(n7819), 
        .Y(n6892) );
  MX4X1 U6267 ( .A(\registers[412][6] ), .B(\registers[413][6] ), .C(
        \registers[414][6] ), .D(\registers[415][6] ), .S0(n7588), .S1(n7819), 
        .Y(n6891) );
  MX4X1 U6268 ( .A(\registers[400][6] ), .B(\registers[401][6] ), .C(
        \registers[402][6] ), .D(\registers[403][6] ), .S0(n7588), .S1(n7819), 
        .Y(n6894) );
  MX4X1 U6269 ( .A(n7000), .B(n6998), .C(n6999), .D(n6997), .S0(n7963), .S1(
        n7898), .Y(n7001) );
  MX4X1 U6270 ( .A(\registers[88][6] ), .B(\registers[89][6] ), .C(
        \registers[90][6] ), .D(\registers[91][6] ), .S0(n7594), .S1(n7825), 
        .Y(n6998) );
  MX4X1 U6271 ( .A(\registers[92][6] ), .B(\registers[93][6] ), .C(
        \registers[94][6] ), .D(\registers[95][6] ), .S0(n7594), .S1(n7825), 
        .Y(n6997) );
  MX4X1 U6272 ( .A(\registers[80][6] ), .B(\registers[81][6] ), .C(
        \registers[82][6] ), .D(\registers[83][6] ), .S0(n7594), .S1(n7825), 
        .Y(n7000) );
  MX4X1 U6273 ( .A(n7021), .B(n7019), .C(n7020), .D(n7018), .S0(n7963), .S1(
        n7898), .Y(n7022) );
  MX4X1 U6274 ( .A(\registers[24][6] ), .B(\registers[25][6] ), .C(
        \registers[26][6] ), .D(\registers[27][6] ), .S0(n7596), .S1(n7826), 
        .Y(n7019) );
  MX4X1 U6275 ( .A(\registers[28][6] ), .B(\registers[29][6] ), .C(
        \registers[30][6] ), .D(\registers[31][6] ), .S0(n7596), .S1(n7826), 
        .Y(n7018) );
  MX4X1 U6276 ( .A(\registers[16][6] ), .B(\registers[17][6] ), .C(
        \registers[18][6] ), .D(\registers[19][6] ), .S0(n7596), .S1(n7826), 
        .Y(n7021) );
  MX4X1 U6277 ( .A(n6958), .B(n6956), .C(n6957), .D(n6955), .S0(n7962), .S1(
        n7898), .Y(n6959) );
  MX4X1 U6278 ( .A(\registers[216][6] ), .B(\registers[217][6] ), .C(
        \registers[218][6] ), .D(\registers[219][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6956) );
  MX4X1 U6279 ( .A(\registers[220][6] ), .B(\registers[221][6] ), .C(
        \registers[222][6] ), .D(\registers[223][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6955) );
  MX4X1 U6280 ( .A(\registers[208][6] ), .B(\registers[209][6] ), .C(
        \registers[210][6] ), .D(\registers[211][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6958) );
  MX4X1 U6281 ( .A(n6979), .B(n6977), .C(n6978), .D(n6976), .S0(n7962), .S1(
        n7898), .Y(n6980) );
  MX4X1 U6282 ( .A(\registers[152][6] ), .B(\registers[153][6] ), .C(
        \registers[154][6] ), .D(\registers[155][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6977) );
  MX4X1 U6283 ( .A(\registers[156][6] ), .B(\registers[157][6] ), .C(
        \registers[158][6] ), .D(\registers[159][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6976) );
  MX4X1 U6284 ( .A(\registers[144][6] ), .B(\registers[145][6] ), .C(
        \registers[146][6] ), .D(\registers[147][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6979) );
  MX4X1 U6285 ( .A(n6745), .B(n6743), .C(n6744), .D(n6742), .S0(n7959), .S1(
        n7896), .Y(n6746) );
  MX4X1 U6286 ( .A(\registers[856][6] ), .B(\registers[857][6] ), .C(
        \registers[858][6] ), .D(\registers[859][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6743) );
  MX4X1 U6287 ( .A(\registers[860][6] ), .B(\registers[861][6] ), .C(
        \registers[862][6] ), .D(\registers[863][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6742) );
  MX4X1 U6288 ( .A(\registers[848][6] ), .B(\registers[849][6] ), .C(
        \registers[850][6] ), .D(\registers[851][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6745) );
  MX4X1 U6289 ( .A(n6766), .B(n6764), .C(n6765), .D(n6763), .S0(n7959), .S1(
        n7901), .Y(n6767) );
  MX4X1 U6290 ( .A(\registers[792][6] ), .B(\registers[793][6] ), .C(
        \registers[794][6] ), .D(\registers[795][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6764) );
  MX4X1 U6291 ( .A(\registers[796][6] ), .B(\registers[797][6] ), .C(
        \registers[798][6] ), .D(\registers[799][6] ), .S0(n7580), .S1(n7811), 
        .Y(n6763) );
  MX4X1 U6292 ( .A(\registers[784][6] ), .B(\registers[785][6] ), .C(
        \registers[786][6] ), .D(\registers[787][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6766) );
  MX4X1 U6293 ( .A(n6703), .B(n6701), .C(n6702), .D(n6700), .S0(n7958), .S1(
        n7896), .Y(n6704) );
  MX4X1 U6294 ( .A(\registers[984][6] ), .B(\registers[985][6] ), .C(
        \registers[986][6] ), .D(\registers[987][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6701) );
  MX4X1 U6295 ( .A(\registers[988][6] ), .B(\registers[989][6] ), .C(
        \registers[990][6] ), .D(\registers[991][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6700) );
  MX4X1 U6296 ( .A(\registers[976][6] ), .B(\registers[977][6] ), .C(
        \registers[978][6] ), .D(\registers[979][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6703) );
  MX4X1 U6297 ( .A(n6724), .B(n6722), .C(n6723), .D(n6721), .S0(n7958), .S1(
        n7896), .Y(n6725) );
  MX4X1 U6298 ( .A(\registers[920][6] ), .B(\registers[921][6] ), .C(
        \registers[922][6] ), .D(\registers[923][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6722) );
  MX4X1 U6299 ( .A(\registers[924][6] ), .B(\registers[925][6] ), .C(
        \registers[926][6] ), .D(\registers[927][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6721) );
  MX4X1 U6300 ( .A(\registers[912][6] ), .B(\registers[913][6] ), .C(
        \registers[914][6] ), .D(\registers[915][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6724) );
  MX4X1 U6301 ( .A(n6830), .B(n6828), .C(n6829), .D(n6827), .S0(n7960), .S1(
        n7888), .Y(n6831) );
  MX4X1 U6302 ( .A(\registers[600][6] ), .B(\registers[601][6] ), .C(
        \registers[602][6] ), .D(\registers[603][6] ), .S0(n7584), .S1(n7815), 
        .Y(n6828) );
  MX4X1 U6303 ( .A(\registers[604][6] ), .B(\registers[605][6] ), .C(
        \registers[606][6] ), .D(\registers[607][6] ), .S0(n7584), .S1(n7815), 
        .Y(n6827) );
  MX4X1 U6304 ( .A(\registers[592][6] ), .B(\registers[593][6] ), .C(
        \registers[594][6] ), .D(\registers[595][6] ), .S0(n7584), .S1(n7815), 
        .Y(n6830) );
  MX4X1 U6305 ( .A(n6851), .B(n6849), .C(n6850), .D(n6848), .S0(n7960), .S1(
        n7902), .Y(n6852) );
  MX4X1 U6306 ( .A(\registers[536][6] ), .B(\registers[537][6] ), .C(
        \registers[538][6] ), .D(\registers[539][6] ), .S0(n7585), .S1(n7816), 
        .Y(n6849) );
  MX4X1 U6307 ( .A(\registers[540][6] ), .B(\registers[541][6] ), .C(
        \registers[542][6] ), .D(\registers[543][6] ), .S0(n7585), .S1(n7816), 
        .Y(n6848) );
  MX4X1 U6308 ( .A(\registers[528][6] ), .B(\registers[529][6] ), .C(
        \registers[530][6] ), .D(\registers[531][6] ), .S0(n7585), .S1(n7817), 
        .Y(n6851) );
  MX4X1 U6309 ( .A(n6788), .B(n6786), .C(n6787), .D(n6785), .S0(n7959), .S1(
        n7892), .Y(n6789) );
  MX4X1 U6310 ( .A(\registers[728][6] ), .B(\registers[729][6] ), .C(
        \registers[730][6] ), .D(\registers[731][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6786) );
  MX4X1 U6311 ( .A(\registers[732][6] ), .B(\registers[733][6] ), .C(
        \registers[734][6] ), .D(\registers[735][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6785) );
  MX4X1 U6312 ( .A(\registers[720][6] ), .B(\registers[721][6] ), .C(
        \registers[722][6] ), .D(\registers[723][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6788) );
  MX4X1 U6313 ( .A(n6809), .B(n6807), .C(n6808), .D(n6806), .S0(n7960), .S1(
        n7867), .Y(n6810) );
  MX4X1 U6314 ( .A(\registers[664][6] ), .B(\registers[665][6] ), .C(
        \registers[666][6] ), .D(\registers[667][6] ), .S0(n7582), .S1(n7814), 
        .Y(n6807) );
  MX4X1 U6315 ( .A(\registers[668][6] ), .B(\registers[669][6] ), .C(
        \registers[670][6] ), .D(\registers[671][6] ), .S0(n7582), .S1(n7814), 
        .Y(n6806) );
  MX4X1 U6316 ( .A(\registers[656][6] ), .B(\registers[657][6] ), .C(
        \registers[658][6] ), .D(\registers[659][6] ), .S0(n7582), .S1(n7814), 
        .Y(n6809) );
  MX4X1 U6317 ( .A(n7255), .B(n7253), .C(n7254), .D(n7252), .S0(n7967), .S1(
        n7896), .Y(n7256) );
  MX4X1 U6318 ( .A(\registers[344][7] ), .B(\registers[345][7] ), .C(
        \registers[346][7] ), .D(\registers[347][7] ), .S0(n7610), .S1(n7840), 
        .Y(n7253) );
  MX4X1 U6319 ( .A(\registers[348][7] ), .B(\registers[349][7] ), .C(
        \registers[350][7] ), .D(\registers[351][7] ), .S0(n7610), .S1(n7840), 
        .Y(n7252) );
  MX4X1 U6320 ( .A(\registers[336][7] ), .B(\registers[337][7] ), .C(
        \registers[338][7] ), .D(\registers[339][7] ), .S0(n7610), .S1(n7840), 
        .Y(n7255) );
  MX4X1 U6321 ( .A(n7213), .B(n7211), .C(n7212), .D(n7210), .S0(n7966), .S1(
        n7901), .Y(n7214) );
  MX4X1 U6322 ( .A(\registers[472][7] ), .B(\registers[473][7] ), .C(
        \registers[474][7] ), .D(\registers[475][7] ), .S0(n7608), .S1(n7837), 
        .Y(n7211) );
  MX4X1 U6323 ( .A(\registers[476][7] ), .B(\registers[477][7] ), .C(
        \registers[478][7] ), .D(\registers[479][7] ), .S0(n7608), .S1(n7837), 
        .Y(n7210) );
  MX4X1 U6324 ( .A(\registers[464][7] ), .B(\registers[465][7] ), .C(
        \registers[466][7] ), .D(\registers[467][7] ), .S0(n7608), .S1(n7838), 
        .Y(n7213) );
  MX4X1 U6325 ( .A(n7234), .B(n7232), .C(n7233), .D(n7231), .S0(n7966), .S1(
        n7896), .Y(n7235) );
  MX4X1 U6326 ( .A(\registers[408][7] ), .B(\registers[409][7] ), .C(
        \registers[410][7] ), .D(\registers[411][7] ), .S0(n7609), .S1(n7839), 
        .Y(n7232) );
  MX4X1 U6327 ( .A(\registers[412][7] ), .B(\registers[413][7] ), .C(
        \registers[414][7] ), .D(\registers[415][7] ), .S0(n7609), .S1(n7839), 
        .Y(n7231) );
  MX4X1 U6328 ( .A(\registers[400][7] ), .B(\registers[401][7] ), .C(
        \registers[402][7] ), .D(\registers[403][7] ), .S0(n7609), .S1(n7839), 
        .Y(n7234) );
  MX4X1 U6329 ( .A(n7276), .B(n7274), .C(n7275), .D(n7273), .S0(n7967), .S1(
        n7897), .Y(n7277) );
  MX4X1 U6330 ( .A(\registers[280][7] ), .B(\registers[281][7] ), .C(
        \registers[282][7] ), .D(\registers[283][7] ), .S0(n7612), .S1(n7841), 
        .Y(n7274) );
  MX4X1 U6331 ( .A(\registers[284][7] ), .B(\registers[285][7] ), .C(
        \registers[286][7] ), .D(\registers[287][7] ), .S0(n7612), .S1(n7841), 
        .Y(n7273) );
  MX4X1 U6332 ( .A(\registers[272][7] ), .B(\registers[273][7] ), .C(
        \registers[274][7] ), .D(\registers[275][7] ), .S0(n7612), .S1(n7841), 
        .Y(n7276) );
  MX4X1 U6333 ( .A(n7298), .B(n7296), .C(n7297), .D(n7295), .S0(n7967), .S1(
        n7869), .Y(n7299) );
  MX4X1 U6334 ( .A(\registers[216][7] ), .B(\registers[217][7] ), .C(
        \registers[218][7] ), .D(\registers[219][7] ), .S0(n7613), .S1(n7842), 
        .Y(n7296) );
  MX4X1 U6335 ( .A(\registers[220][7] ), .B(\registers[221][7] ), .C(
        \registers[222][7] ), .D(\registers[223][7] ), .S0(n7613), .S1(n7842), 
        .Y(n7295) );
  MX4X1 U6336 ( .A(\registers[208][7] ), .B(\registers[209][7] ), .C(
        \registers[210][7] ), .D(\registers[211][7] ), .S0(n7613), .S1(n7842), 
        .Y(n7298) );
  MX4X1 U6337 ( .A(n7340), .B(n7338), .C(n7339), .D(n7337), .S0(n7962), .S1(
        n7902), .Y(n7341) );
  MX4X1 U6338 ( .A(\registers[88][7] ), .B(\registers[89][7] ), .C(
        \registers[90][7] ), .D(\registers[91][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7338) );
  MX4X1 U6339 ( .A(\registers[92][7] ), .B(\registers[93][7] ), .C(
        \registers[94][7] ), .D(\registers[95][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7337) );
  MX4X1 U6340 ( .A(\registers[80][7] ), .B(\registers[81][7] ), .C(
        \registers[82][7] ), .D(\registers[83][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7340) );
  MX4X1 U6341 ( .A(n7361), .B(n7359), .C(n7360), .D(n7358), .S0(N81), .S1(
        n7902), .Y(n7362) );
  MX4X1 U6342 ( .A(\registers[24][7] ), .B(\registers[25][7] ), .C(
        \registers[26][7] ), .D(\registers[27][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7359) );
  MX4X1 U6343 ( .A(\registers[28][7] ), .B(\registers[29][7] ), .C(
        \registers[30][7] ), .D(\registers[31][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7358) );
  MX4X1 U6344 ( .A(\registers[16][7] ), .B(\registers[17][7] ), .C(
        \registers[18][7] ), .D(\registers[19][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7361) );
  MX4X1 U6345 ( .A(n7319), .B(n7317), .C(n7318), .D(n7316), .S0(N81), .S1(
        n7902), .Y(n7320) );
  MX4X1 U6346 ( .A(\registers[152][7] ), .B(\registers[153][7] ), .C(
        \registers[154][7] ), .D(\registers[155][7] ), .S0(n7614), .S1(n7844), 
        .Y(n7317) );
  MX4X1 U6347 ( .A(\registers[156][7] ), .B(\registers[157][7] ), .C(
        \registers[158][7] ), .D(\registers[159][7] ), .S0(n7614), .S1(n7843), 
        .Y(n7316) );
  MX4X1 U6348 ( .A(\registers[144][7] ), .B(\registers[145][7] ), .C(
        \registers[146][7] ), .D(\registers[147][7] ), .S0(n7614), .S1(n7844), 
        .Y(n7319) );
  MX4X1 U6349 ( .A(n7085), .B(n7083), .C(n7084), .D(n7082), .S0(n7964), .S1(
        n7899), .Y(n7086) );
  MX4X1 U6350 ( .A(\registers[856][7] ), .B(\registers[857][7] ), .C(
        \registers[858][7] ), .D(\registers[859][7] ), .S0(n7600), .S1(n7830), 
        .Y(n7083) );
  MX4X1 U6351 ( .A(\registers[860][7] ), .B(\registers[861][7] ), .C(
        \registers[862][7] ), .D(\registers[863][7] ), .S0(n7600), .S1(n7830), 
        .Y(n7082) );
  MX4X1 U6352 ( .A(\registers[848][7] ), .B(\registers[849][7] ), .C(
        \registers[850][7] ), .D(\registers[851][7] ), .S0(n7600), .S1(n7830), 
        .Y(n7085) );
  MX4X1 U6353 ( .A(n7106), .B(n7104), .C(n7105), .D(n7103), .S0(n7964), .S1(
        n7900), .Y(n7107) );
  MX4X1 U6354 ( .A(\registers[792][7] ), .B(\registers[793][7] ), .C(
        \registers[794][7] ), .D(\registers[795][7] ), .S0(n7601), .S1(n7831), 
        .Y(n7104) );
  MX4X1 U6355 ( .A(\registers[796][7] ), .B(\registers[797][7] ), .C(
        \registers[798][7] ), .D(\registers[799][7] ), .S0(n7601), .S1(n7831), 
        .Y(n7103) );
  MX4X1 U6356 ( .A(\registers[784][7] ), .B(\registers[785][7] ), .C(
        \registers[786][7] ), .D(\registers[787][7] ), .S0(n7601), .S1(n7831), 
        .Y(n7106) );
  MX4X1 U6357 ( .A(n7043), .B(n7041), .C(n7042), .D(n7040), .S0(n7963), .S1(
        n7899), .Y(n7044) );
  MX4X1 U6358 ( .A(\registers[984][7] ), .B(\registers[985][7] ), .C(
        \registers[986][7] ), .D(\registers[987][7] ), .S0(n7597), .S1(n7828), 
        .Y(n7041) );
  MX4X1 U6359 ( .A(\registers[988][7] ), .B(\registers[989][7] ), .C(
        \registers[990][7] ), .D(\registers[991][7] ), .S0(n7597), .S1(n7827), 
        .Y(n7040) );
  MX4X1 U6360 ( .A(\registers[976][7] ), .B(\registers[977][7] ), .C(
        \registers[978][7] ), .D(\registers[979][7] ), .S0(n7597), .S1(n7828), 
        .Y(n7043) );
  MX4X1 U6361 ( .A(n7064), .B(n7062), .C(n7063), .D(n7061), .S0(n7964), .S1(
        n7899), .Y(n7065) );
  MX4X1 U6362 ( .A(\registers[920][7] ), .B(\registers[921][7] ), .C(
        \registers[922][7] ), .D(\registers[923][7] ), .S0(n7598), .S1(n7829), 
        .Y(n7062) );
  MX4X1 U6363 ( .A(\registers[924][7] ), .B(\registers[925][7] ), .C(
        \registers[926][7] ), .D(\registers[927][7] ), .S0(n7598), .S1(n7829), 
        .Y(n7061) );
  MX4X1 U6364 ( .A(\registers[912][7] ), .B(\registers[913][7] ), .C(
        \registers[914][7] ), .D(\registers[915][7] ), .S0(n7598), .S1(n7829), 
        .Y(n7064) );
  MX4X1 U6365 ( .A(n7170), .B(n7168), .C(n7169), .D(n7167), .S0(n7965), .S1(
        n7901), .Y(n7171) );
  MX4X1 U6366 ( .A(\registers[600][7] ), .B(\registers[601][7] ), .C(
        \registers[602][7] ), .D(\registers[603][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7168) );
  MX4X1 U6367 ( .A(\registers[604][7] ), .B(\registers[605][7] ), .C(
        \registers[606][7] ), .D(\registers[607][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7167) );
  MX4X1 U6368 ( .A(\registers[592][7] ), .B(\registers[593][7] ), .C(
        \registers[594][7] ), .D(\registers[595][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7170) );
  MX4X1 U6369 ( .A(n7191), .B(n7189), .C(n7190), .D(n7188), .S0(n7966), .S1(
        n7901), .Y(n7192) );
  MX4X1 U6370 ( .A(\registers[536][7] ), .B(\registers[537][7] ), .C(
        \registers[538][7] ), .D(\registers[539][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7189) );
  MX4X1 U6371 ( .A(\registers[540][7] ), .B(\registers[541][7] ), .C(
        \registers[542][7] ), .D(\registers[543][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7188) );
  MX4X1 U6372 ( .A(\registers[528][7] ), .B(\registers[529][7] ), .C(
        \registers[530][7] ), .D(\registers[531][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7191) );
  MX4X1 U6373 ( .A(n7128), .B(n7126), .C(n7127), .D(n7125), .S0(n7965), .S1(
        n7900), .Y(n7129) );
  MX4X1 U6374 ( .A(\registers[728][7] ), .B(\registers[729][7] ), .C(
        \registers[730][7] ), .D(\registers[731][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7126) );
  MX4X1 U6375 ( .A(\registers[732][7] ), .B(\registers[733][7] ), .C(
        \registers[734][7] ), .D(\registers[735][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7125) );
  MX4X1 U6376 ( .A(\registers[720][7] ), .B(\registers[721][7] ), .C(
        \registers[722][7] ), .D(\registers[723][7] ), .S0(n7602), .S1(n7833), 
        .Y(n7128) );
  MX4X1 U6377 ( .A(n7149), .B(n7147), .C(n7148), .D(n7146), .S0(n7965), .S1(
        n7900), .Y(n7150) );
  MX4X1 U6378 ( .A(\registers[664][7] ), .B(\registers[665][7] ), .C(
        \registers[666][7] ), .D(\registers[667][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7147) );
  MX4X1 U6379 ( .A(\registers[668][7] ), .B(\registers[669][7] ), .C(
        \registers[670][7] ), .D(\registers[671][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7146) );
  MX4X1 U6380 ( .A(\registers[656][7] ), .B(\registers[657][7] ), .C(
        \registers[658][7] ), .D(\registers[659][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7149) );
  MX4X1 U6381 ( .A(\registers[1008][0] ), .B(\registers[1009][0] ), .C(
        \registers[1010][0] ), .D(\registers[1011][0] ), .S0(n4242), .S1(n4460), .Y(n1048) );
  MX4X1 U6382 ( .A(\registers[992][0] ), .B(\registers[993][0] ), .C(
        \registers[994][0] ), .D(\registers[995][0] ), .S0(n4270), .S1(n4349), 
        .Y(n1053) );
  MX4X1 U6383 ( .A(\registers[1008][0] ), .B(\registers[1009][0] ), .C(
        \registers[1010][0] ), .D(\registers[1011][0] ), .S0(n7564), .S1(n7810), .Y(n4653) );
  MX4X1 U6384 ( .A(\registers[992][0] ), .B(\registers[993][0] ), .C(
        \registers[994][0] ), .D(\registers[995][0] ), .S0(n7565), .S1(n7691), 
        .Y(n4658) );
  MX4X1 U6385 ( .A(\registers[320][0] ), .B(\registers[321][0] ), .C(
        \registers[322][0] ), .D(\registers[323][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1431) );
  MX4X1 U6386 ( .A(\registers[368][0] ), .B(\registers[369][0] ), .C(
        \registers[370][0] ), .D(\registers[371][0] ), .S0(n4117), .S1(n4359), 
        .Y(n1416) );
  MX4X1 U6387 ( .A(\registers[352][0] ), .B(\registers[353][0] ), .C(
        \registers[354][0] ), .D(\registers[355][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1421) );
  MX4X1 U6388 ( .A(\registers[64][0] ), .B(\registers[65][0] ), .C(
        \registers[66][0] ), .D(\registers[67][0] ), .S0(n4124), .S1(n4364), 
        .Y(n1522) );
  MX4X1 U6389 ( .A(\registers[112][0] ), .B(\registers[113][0] ), .C(
        \registers[114][0] ), .D(\registers[115][0] ), .S0(n4123), .S1(n4363), 
        .Y(n1507) );
  MX4X1 U6390 ( .A(\registers[96][0] ), .B(\registers[97][0] ), .C(
        \registers[98][0] ), .D(\registers[99][0] ), .S0(n4123), .S1(n4364), 
        .Y(n1512) );
  MX4X1 U6391 ( .A(\registers[0][0] ), .B(\registers[1][0] ), .C(
        \registers[2][0] ), .D(\registers[3][0] ), .S0(n4125), .S1(n4366), .Y(
        n1545) );
  MX4X1 U6392 ( .A(\registers[48][0] ), .B(\registers[49][0] ), .C(
        \registers[50][0] ), .D(\registers[51][0] ), .S0(n4124), .S1(n4365), 
        .Y(n1528) );
  MX4X1 U6393 ( .A(\registers[32][0] ), .B(\registers[33][0] ), .C(
        \registers[34][0] ), .D(\registers[35][0] ), .S0(n4124), .S1(n4365), 
        .Y(n1533) );
  MX4X1 U6394 ( .A(\registers[192][0] ), .B(\registers[193][0] ), .C(
        \registers[194][0] ), .D(\registers[195][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1478) );
  MX4X1 U6395 ( .A(\registers[240][0] ), .B(\registers[241][0] ), .C(
        \registers[242][0] ), .D(\registers[243][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1461) );
  MX4X1 U6396 ( .A(\registers[224][0] ), .B(\registers[225][0] ), .C(
        \registers[226][0] ), .D(\registers[227][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1466) );
  MX4X1 U6397 ( .A(\registers[128][0] ), .B(\registers[129][0] ), .C(
        \registers[130][0] ), .D(\registers[131][0] ), .S0(n4122), .S1(n4363), 
        .Y(n1499) );
  MX4X1 U6398 ( .A(\registers[176][0] ), .B(\registers[177][0] ), .C(
        \registers[178][0] ), .D(\registers[179][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1484) );
  MX4X1 U6399 ( .A(\registers[160][0] ), .B(\registers[161][0] ), .C(
        \registers[162][0] ), .D(\registers[163][0] ), .S0(n4122), .S1(n4363), 
        .Y(n1489) );
  MX4X1 U6400 ( .A(\registers[832][0] ), .B(\registers[833][0] ), .C(
        \registers[834][0] ), .D(\registers[835][0] ), .S0(n4108), .S1(n4405), 
        .Y(n1105) );
  MX4X1 U6401 ( .A(\registers[880][0] ), .B(\registers[881][0] ), .C(
        \registers[882][0] ), .D(\registers[883][0] ), .S0(n4107), .S1(n4486), 
        .Y(n1090) );
  MX4X1 U6402 ( .A(\registers[864][0] ), .B(\registers[865][0] ), .C(
        \registers[866][0] ), .D(\registers[867][0] ), .S0(n4107), .S1(n4455), 
        .Y(n1095) );
  MX4X1 U6403 ( .A(\registers[768][0] ), .B(\registers[769][0] ), .C(
        \registers[770][0] ), .D(\registers[771][0] ), .S0(n4109), .S1(n4351), 
        .Y(n1168) );
  MX4X1 U6404 ( .A(\registers[816][0] ), .B(\registers[817][0] ), .C(
        \registers[818][0] ), .D(\registers[819][0] ), .S0(n4108), .S1(n4425), 
        .Y(n1153) );
  MX4X1 U6405 ( .A(\registers[800][0] ), .B(\registers[801][0] ), .C(
        \registers[802][0] ), .D(\registers[803][0] ), .S0(n4108), .S1(n4376), 
        .Y(n1158) );
  MX4X1 U6406 ( .A(\registers[960][0] ), .B(\registers[961][0] ), .C(
        \registers[962][0] ), .D(\registers[963][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1063) );
  MX4X1 U6407 ( .A(\registers[896][0] ), .B(\registers[897][0] ), .C(
        \registers[898][0] ), .D(\registers[899][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1084) );
  MX4X1 U6408 ( .A(\registers[944][0] ), .B(\registers[945][0] ), .C(
        \registers[946][0] ), .D(\registers[947][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1069) );
  MX4X1 U6409 ( .A(\registers[928][0] ), .B(\registers[929][0] ), .C(
        \registers[930][0] ), .D(\registers[931][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1074) );
  MX4X1 U6410 ( .A(\registers[576][0] ), .B(\registers[577][0] ), .C(
        \registers[578][0] ), .D(\registers[579][0] ), .S0(n4113), .S1(n4355), 
        .Y(n1341) );
  MX4X1 U6411 ( .A(\registers[624][0] ), .B(\registers[625][0] ), .C(
        \registers[626][0] ), .D(\registers[627][0] ), .S0(n4112), .S1(n4354), 
        .Y(n1317) );
  MX4X1 U6412 ( .A(\registers[608][0] ), .B(\registers[609][0] ), .C(
        \registers[610][0] ), .D(\registers[611][0] ), .S0(n4112), .S1(n4354), 
        .Y(n1327) );
  MX4X1 U6413 ( .A(\registers[512][0] ), .B(\registers[513][0] ), .C(
        \registers[514][0] ), .D(\registers[515][0] ), .S0(n4114), .S1(n4356), 
        .Y(n1362) );
  MX4X1 U6414 ( .A(\registers[560][0] ), .B(\registers[561][0] ), .C(
        \registers[562][0] ), .D(\registers[563][0] ), .S0(n4113), .S1(n4355), 
        .Y(n1347) );
  MX4X1 U6415 ( .A(\registers[544][0] ), .B(\registers[545][0] ), .C(
        \registers[546][0] ), .D(\registers[547][0] ), .S0(n4114), .S1(n4355), 
        .Y(n1352) );
  MX4X1 U6416 ( .A(\registers[704][0] ), .B(\registers[705][0] ), .C(
        \registers[706][0] ), .D(\registers[707][0] ), .S0(n4110), .S1(n4352), 
        .Y(n1205) );
  MX4X1 U6417 ( .A(\registers[752][0] ), .B(\registers[753][0] ), .C(
        \registers[754][0] ), .D(\registers[755][0] ), .S0(n4109), .S1(n4351), 
        .Y(n1175) );
  MX4X1 U6418 ( .A(\registers[736][0] ), .B(\registers[737][0] ), .C(
        \registers[738][0] ), .D(\registers[739][0] ), .S0(n4110), .S1(n4351), 
        .Y(n1180) );
  MX4X1 U6419 ( .A(\registers[640][0] ), .B(\registers[641][0] ), .C(
        \registers[642][0] ), .D(\registers[643][0] ), .S0(n4112), .S1(n4353), 
        .Y(n1305) );
  MX4X1 U6420 ( .A(\registers[688][0] ), .B(\registers[689][0] ), .C(
        \registers[690][0] ), .D(\registers[691][0] ), .S0(n4111), .S1(n4352), 
        .Y(n1275) );
  MX4X1 U6421 ( .A(\registers[672][0] ), .B(\registers[673][0] ), .C(
        \registers[674][0] ), .D(\registers[675][0] ), .S0(n4111), .S1(n4353), 
        .Y(n1285) );
  MX4X1 U6422 ( .A(\registers[320][1] ), .B(\registers[321][1] ), .C(
        \registers[322][1] ), .D(\registers[323][1] ), .S0(n4140), .S1(n4379), 
        .Y(n1789) );
  MX4X1 U6423 ( .A(\registers[368][1] ), .B(\registers[369][1] ), .C(
        \registers[370][1] ), .D(\registers[371][1] ), .S0(n4139), .S1(n4378), 
        .Y(n1774) );
  MX4X1 U6424 ( .A(\registers[352][1] ), .B(\registers[353][1] ), .C(
        \registers[354][1] ), .D(\registers[355][1] ), .S0(n4139), .S1(n4379), 
        .Y(n1779) );
  MX4X1 U6425 ( .A(\registers[64][1] ), .B(\registers[65][1] ), .C(
        \registers[66][1] ), .D(\registers[67][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1878) );
  MX4X1 U6426 ( .A(\registers[112][1] ), .B(\registers[113][1] ), .C(
        \registers[114][1] ), .D(\registers[115][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1861) );
  MX4X1 U6427 ( .A(\registers[96][1] ), .B(\registers[97][1] ), .C(
        \registers[98][1] ), .D(\registers[99][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1866) );
  MX4X1 U6428 ( .A(\registers[0][1] ), .B(\registers[1][1] ), .C(
        \registers[2][1] ), .D(\registers[3][1] ), .S0(n4146), .S1(n4385), .Y(
        n1899) );
  MX4X1 U6429 ( .A(\registers[48][1] ), .B(\registers[49][1] ), .C(
        \registers[50][1] ), .D(\registers[51][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1884) );
  MX4X1 U6430 ( .A(\registers[32][1] ), .B(\registers[33][1] ), .C(
        \registers[34][1] ), .D(\registers[35][1] ), .S0(n4146), .S1(n4385), 
        .Y(n1889) );
  MX4X1 U6431 ( .A(\registers[192][1] ), .B(\registers[193][1] ), .C(
        \registers[194][1] ), .D(\registers[195][1] ), .S0(n4142), .S1(n4382), 
        .Y(n1833) );
  MX4X1 U6432 ( .A(\registers[240][1] ), .B(\registers[241][1] ), .C(
        \registers[242][1] ), .D(\registers[243][1] ), .S0(n4141), .S1(n4381), 
        .Y(n1818) );
  MX4X1 U6433 ( .A(\registers[224][1] ), .B(\registers[225][1] ), .C(
        \registers[226][1] ), .D(\registers[227][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1823) );
  MX4X1 U6434 ( .A(\registers[128][1] ), .B(\registers[129][1] ), .C(
        \registers[130][1] ), .D(\registers[131][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1855) );
  MX4X1 U6435 ( .A(\registers[176][1] ), .B(\registers[177][1] ), .C(
        \registers[178][1] ), .D(\registers[179][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1840) );
  MX4X1 U6436 ( .A(\registers[160][1] ), .B(\registers[161][1] ), .C(
        \registers[162][1] ), .D(\registers[163][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1845) );
  MX4X1 U6437 ( .A(\registers[832][1] ), .B(\registers[833][1] ), .C(
        \registers[834][1] ), .D(\registers[835][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1614) );
  MX4X1 U6438 ( .A(\registers[880][1] ), .B(\registers[881][1] ), .C(
        \registers[882][1] ), .D(\registers[883][1] ), .S0(n4128), .S1(n4368), 
        .Y(n1596) );
  MX4X1 U6439 ( .A(\registers[864][1] ), .B(\registers[865][1] ), .C(
        \registers[866][1] ), .D(\registers[867][1] ), .S0(n4128), .S1(n4369), 
        .Y(n1601) );
  MX4X1 U6440 ( .A(\registers[768][1] ), .B(\registers[769][1] ), .C(
        \registers[770][1] ), .D(\registers[771][1] ), .S0(n4130), .S1(n4371), 
        .Y(n1635) );
  MX4X1 U6441 ( .A(\registers[816][1] ), .B(\registers[817][1] ), .C(
        \registers[818][1] ), .D(\registers[819][1] ), .S0(n4129), .S1(n4370), 
        .Y(n1620) );
  MX4X1 U6442 ( .A(\registers[800][1] ), .B(\registers[801][1] ), .C(
        \registers[802][1] ), .D(\registers[803][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1625) );
  MX4X1 U6443 ( .A(\registers[960][1] ), .B(\registers[961][1] ), .C(
        \registers[962][1] ), .D(\registers[963][1] ), .S0(n4126), .S1(n4367), 
        .Y(n1567) );
  MX4X1 U6444 ( .A(\registers[1008][1] ), .B(\registers[1009][1] ), .C(
        \registers[1010][1] ), .D(\registers[1011][1] ), .S0(n4125), .S1(n4366), .Y(n1552) );
  MX4X1 U6445 ( .A(\registers[992][1] ), .B(\registers[993][1] ), .C(
        \registers[994][1] ), .D(\registers[995][1] ), .S0(n4126), .S1(n4366), 
        .Y(n1557) );
  MX4X1 U6446 ( .A(\registers[896][1] ), .B(\registers[897][1] ), .C(
        \registers[898][1] ), .D(\registers[899][1] ), .S0(n4128), .S1(n4368), 
        .Y(n1590) );
  MX4X1 U6447 ( .A(\registers[944][1] ), .B(\registers[945][1] ), .C(
        \registers[946][1] ), .D(\registers[947][1] ), .S0(n4127), .S1(n4367), 
        .Y(n1575) );
  MX4X1 U6448 ( .A(\registers[928][1] ), .B(\registers[929][1] ), .C(
        \registers[930][1] ), .D(\registers[931][1] ), .S0(n4127), .S1(n4367), 
        .Y(n1580) );
  MX4X1 U6449 ( .A(\registers[576][1] ), .B(\registers[577][1] ), .C(
        \registers[578][1] ), .D(\registers[579][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1701) );
  MX4X1 U6450 ( .A(\registers[624][1] ), .B(\registers[625][1] ), .C(
        \registers[626][1] ), .D(\registers[627][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1686) );
  MX4X1 U6451 ( .A(\registers[608][1] ), .B(\registers[609][1] ), .C(
        \registers[610][1] ), .D(\registers[611][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1691) );
  MX4X1 U6452 ( .A(\registers[512][1] ), .B(\registers[513][1] ), .C(
        \registers[514][1] ), .D(\registers[515][1] ), .S0(n4136), .S1(n4375), 
        .Y(n1723) );
  MX4X1 U6453 ( .A(\registers[560][1] ), .B(\registers[561][1] ), .C(
        \registers[562][1] ), .D(\registers[563][1] ), .S0(n4135), .S1(n4375), 
        .Y(n1708) );
  MX4X1 U6454 ( .A(\registers[544][1] ), .B(\registers[545][1] ), .C(
        \registers[546][1] ), .D(\registers[547][1] ), .S0(n4135), .S1(n4375), 
        .Y(n1713) );
  MX4X1 U6455 ( .A(\registers[704][1] ), .B(\registers[705][1] ), .C(
        \registers[706][1] ), .D(\registers[707][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1658) );
  MX4X1 U6456 ( .A(\registers[752][1] ), .B(\registers[753][1] ), .C(
        \registers[754][1] ), .D(\registers[755][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1643) );
  MX4X1 U6457 ( .A(\registers[736][1] ), .B(\registers[737][1] ), .C(
        \registers[738][1] ), .D(\registers[739][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1648) );
  MX4X1 U6458 ( .A(\registers[640][1] ), .B(\registers[641][1] ), .C(
        \registers[642][1] ), .D(\registers[643][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1680) );
  MX4X1 U6459 ( .A(\registers[688][1] ), .B(\registers[689][1] ), .C(
        \registers[690][1] ), .D(\registers[691][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1664) );
  MX4X1 U6460 ( .A(\registers[672][1] ), .B(\registers[673][1] ), .C(
        \registers[674][1] ), .D(\registers[675][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1669) );
  MX4X1 U6461 ( .A(\registers[320][2] ), .B(\registers[321][2] ), .C(
        \registers[322][2] ), .D(\registers[323][2] ), .S0(n4161), .S1(n4399), 
        .Y(n2142) );
  MX4X1 U6462 ( .A(\registers[368][2] ), .B(\registers[369][2] ), .C(
        \registers[370][2] ), .D(\registers[371][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2125) );
  MX4X1 U6463 ( .A(\registers[352][2] ), .B(\registers[353][2] ), .C(
        \registers[354][2] ), .D(\registers[355][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2130) );
  MX4X1 U6464 ( .A(\registers[64][2] ), .B(\registers[65][2] ), .C(
        \registers[66][2] ), .D(\registers[67][2] ), .S0(n4166), .S1(n4404), 
        .Y(n2229) );
  MX4X1 U6465 ( .A(\registers[112][2] ), .B(\registers[113][2] ), .C(
        \registers[114][2] ), .D(\registers[115][2] ), .S0(n4165), .S1(n4403), 
        .Y(n2214) );
  MX4X1 U6466 ( .A(\registers[96][2] ), .B(\registers[97][2] ), .C(
        \registers[98][2] ), .D(\registers[99][2] ), .S0(n4166), .S1(n4403), 
        .Y(n2219) );
  MX4X1 U6467 ( .A(\registers[0][2] ), .B(\registers[1][2] ), .C(
        \registers[2][2] ), .D(\registers[3][2] ), .S0(n4168), .S1(n4405), .Y(
        n2251) );
  MX4X1 U6468 ( .A(\registers[48][2] ), .B(\registers[49][2] ), .C(
        \registers[50][2] ), .D(\registers[51][2] ), .S0(n4167), .S1(n4404), 
        .Y(n2235) );
  MX4X1 U6469 ( .A(\registers[32][2] ), .B(\registers[33][2] ), .C(
        \registers[34][2] ), .D(\registers[35][2] ), .S0(n4167), .S1(n4404), 
        .Y(n2241) );
  MX4X1 U6470 ( .A(\registers[192][2] ), .B(\registers[193][2] ), .C(
        \registers[194][2] ), .D(\registers[195][2] ), .S0(n4164), .S1(n4401), 
        .Y(n2186) );
  MX4X1 U6471 ( .A(\registers[240][2] ), .B(\registers[241][2] ), .C(
        \registers[242][2] ), .D(\registers[243][2] ), .S0(n4163), .S1(n4400), 
        .Y(n2170) );
  MX4X1 U6472 ( .A(\registers[224][2] ), .B(\registers[225][2] ), .C(
        \registers[226][2] ), .D(\registers[227][2] ), .S0(n4163), .S1(n4401), 
        .Y(n2176) );
  MX4X1 U6473 ( .A(\registers[128][2] ), .B(\registers[129][2] ), .C(
        \registers[130][2] ), .D(\registers[131][2] ), .S0(n4165), .S1(n4403), 
        .Y(n2208) );
  MX4X1 U6474 ( .A(\registers[176][2] ), .B(\registers[177][2] ), .C(
        \registers[178][2] ), .D(\registers[179][2] ), .S0(n4164), .S1(n4402), 
        .Y(n2192) );
  MX4X1 U6475 ( .A(\registers[160][2] ), .B(\registers[161][2] ), .C(
        \registers[162][2] ), .D(\registers[163][2] ), .S0(n4164), .S1(n4402), 
        .Y(n2197) );
  MX4X1 U6476 ( .A(\registers[832][2] ), .B(\registers[833][2] ), .C(
        \registers[834][2] ), .D(\registers[835][2] ), .S0(n4150), .S1(n4389), 
        .Y(n1965) );
  MX4X1 U6477 ( .A(\registers[880][2] ), .B(\registers[881][2] ), .C(
        \registers[882][2] ), .D(\registers[883][2] ), .S0(n4149), .S1(n4388), 
        .Y(n1950) );
  MX4X1 U6478 ( .A(\registers[864][2] ), .B(\registers[865][2] ), .C(
        \registers[866][2] ), .D(\registers[867][2] ), .S0(n4150), .S1(n4388), 
        .Y(n1955) );
  MX4X1 U6479 ( .A(\registers[768][2] ), .B(\registers[769][2] ), .C(
        \registers[770][2] ), .D(\registers[771][2] ), .S0(n4152), .S1(n4390), 
        .Y(n1987) );
  MX4X1 U6480 ( .A(\registers[816][2] ), .B(\registers[817][2] ), .C(
        \registers[818][2] ), .D(\registers[819][2] ), .S0(n4151), .S1(n4389), 
        .Y(n1971) );
  MX4X1 U6481 ( .A(\registers[800][2] ), .B(\registers[801][2] ), .C(
        \registers[802][2] ), .D(\registers[803][2] ), .S0(n4151), .S1(n4390), 
        .Y(n1977) );
  MX4X1 U6482 ( .A(\registers[960][2] ), .B(\registers[961][2] ), .C(
        \registers[962][2] ), .D(\registers[963][2] ), .S0(n4148), .S1(n4387), 
        .Y(n1922) );
  MX4X1 U6483 ( .A(\registers[1008][2] ), .B(\registers[1009][2] ), .C(
        \registers[1010][2] ), .D(\registers[1011][2] ), .S0(n4147), .S1(n4386), .Y(n1907) );
  MX4X1 U6484 ( .A(\registers[992][2] ), .B(\registers[993][2] ), .C(
        \registers[994][2] ), .D(\registers[995][2] ), .S0(n4147), .S1(n4386), 
        .Y(n1912) );
  MX4X1 U6485 ( .A(\registers[896][2] ), .B(\registers[897][2] ), .C(
        \registers[898][2] ), .D(\registers[899][2] ), .S0(n4149), .S1(n4388), 
        .Y(n1944) );
  MX4X1 U6486 ( .A(\registers[944][2] ), .B(\registers[945][2] ), .C(
        \registers[946][2] ), .D(\registers[947][2] ), .S0(n4148), .S1(n4387), 
        .Y(n1928) );
  MX4X1 U6487 ( .A(\registers[928][2] ), .B(\registers[929][2] ), .C(
        \registers[930][2] ), .D(\registers[931][2] ), .S0(n4148), .S1(n4387), 
        .Y(n1933) );
  MX4X1 U6488 ( .A(\registers[576][2] ), .B(\registers[577][2] ), .C(
        \registers[578][2] ), .D(\registers[579][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2053) );
  MX4X1 U6489 ( .A(\registers[624][2] ), .B(\registers[625][2] ), .C(
        \registers[626][2] ), .D(\registers[627][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2037) );
  MX4X1 U6490 ( .A(\registers[608][2] ), .B(\registers[609][2] ), .C(
        \registers[610][2] ), .D(\registers[611][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2043) );
  MX4X1 U6491 ( .A(\registers[512][2] ), .B(\registers[513][2] ), .C(
        \registers[514][2] ), .D(\registers[515][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2075) );
  MX4X1 U6492 ( .A(\registers[560][2] ), .B(\registers[561][2] ), .C(
        \registers[562][2] ), .D(\registers[563][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2059) );
  MX4X1 U6493 ( .A(\registers[544][2] ), .B(\registers[545][2] ), .C(
        \registers[546][2] ), .D(\registers[547][2] ), .S0(n4156), .S1(n4395), 
        .Y(n2064) );
  MX4X1 U6494 ( .A(\registers[704][2] ), .B(\registers[705][2] ), .C(
        \registers[706][2] ), .D(\registers[707][2] ), .S0(n4153), .S1(n4391), 
        .Y(n2010) );
  MX4X1 U6495 ( .A(\registers[752][2] ), .B(\registers[753][2] ), .C(
        \registers[754][2] ), .D(\registers[755][2] ), .S0(n4152), .S1(n4391), 
        .Y(n1994) );
  MX4X1 U6496 ( .A(\registers[736][2] ), .B(\registers[737][2] ), .C(
        \registers[738][2] ), .D(\registers[739][2] ), .S0(n4152), .S1(n4391), 
        .Y(n1999) );
  MX4X1 U6497 ( .A(\registers[640][2] ), .B(\registers[641][2] ), .C(
        \registers[642][2] ), .D(\registers[643][2] ), .S0(n4154), .S1(n4393), 
        .Y(n2031) );
  MX4X1 U6498 ( .A(\registers[688][2] ), .B(\registers[689][2] ), .C(
        \registers[690][2] ), .D(\registers[691][2] ), .S0(n4153), .S1(n4392), 
        .Y(n2016) );
  MX4X1 U6499 ( .A(\registers[672][2] ), .B(\registers[673][2] ), .C(
        \registers[674][2] ), .D(\registers[675][2] ), .S0(n4154), .S1(n4392), 
        .Y(n2021) );
  MX4X1 U6500 ( .A(\registers[320][3] ), .B(\registers[321][3] ), .C(
        \registers[322][3] ), .D(\registers[323][3] ), .S0(n4182), .S1(n4419), 
        .Y(n2555) );
  MX4X1 U6501 ( .A(\registers[368][3] ), .B(\registers[369][3] ), .C(
        \registers[370][3] ), .D(\registers[371][3] ), .S0(n4181), .S1(n4418), 
        .Y(n2540) );
  MX4X1 U6502 ( .A(\registers[352][3] ), .B(\registers[353][3] ), .C(
        \registers[354][3] ), .D(\registers[355][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2545) );
  MX4X1 U6503 ( .A(\registers[64][3] ), .B(\registers[65][3] ), .C(
        \registers[66][3] ), .D(\registers[67][3] ), .S0(n4188), .S1(n4423), 
        .Y(n2640) );
  MX4X1 U6504 ( .A(\registers[112][3] ), .B(\registers[113][3] ), .C(
        \registers[114][3] ), .D(\registers[115][3] ), .S0(n4187), .S1(n4423), 
        .Y(n2625) );
  MX4X1 U6505 ( .A(\registers[96][3] ), .B(\registers[97][3] ), .C(
        \registers[98][3] ), .D(\registers[99][3] ), .S0(n4187), .S1(n4423), 
        .Y(n2630) );
  MX4X1 U6506 ( .A(\registers[0][3] ), .B(\registers[1][3] ), .C(
        \registers[2][3] ), .D(\registers[3][3] ), .S0(n4189), .S1(n4425), .Y(
        n2661) );
  MX4X1 U6507 ( .A(\registers[48][3] ), .B(\registers[49][3] ), .C(
        \registers[50][3] ), .D(\registers[51][3] ), .S0(n4188), .S1(n4424), 
        .Y(n2646) );
  MX4X1 U6508 ( .A(\registers[32][3] ), .B(\registers[33][3] ), .C(
        \registers[34][3] ), .D(\registers[35][3] ), .S0(n4188), .S1(n4424), 
        .Y(n2651) );
  MX4X1 U6509 ( .A(\registers[192][3] ), .B(\registers[193][3] ), .C(
        \registers[194][3] ), .D(\registers[195][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2598) );
  MX4X1 U6510 ( .A(\registers[240][3] ), .B(\registers[241][3] ), .C(
        \registers[242][3] ), .D(\registers[243][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2583) );
  MX4X1 U6511 ( .A(\registers[224][3] ), .B(\registers[225][3] ), .C(
        \registers[226][3] ), .D(\registers[227][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2588) );
  MX4X1 U6512 ( .A(\registers[128][3] ), .B(\registers[129][3] ), .C(
        \registers[130][3] ), .D(\registers[131][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2619) );
  MX4X1 U6513 ( .A(\registers[176][3] ), .B(\registers[177][3] ), .C(
        \registers[178][3] ), .D(\registers[179][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2604) );
  MX4X1 U6514 ( .A(\registers[160][3] ), .B(\registers[161][3] ), .C(
        \registers[162][3] ), .D(\registers[163][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2609) );
  MX4X1 U6515 ( .A(\registers[832][3] ), .B(\registers[833][3] ), .C(
        \registers[834][3] ), .D(\registers[835][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2317) );
  MX4X1 U6516 ( .A(\registers[880][3] ), .B(\registers[881][3] ), .C(
        \registers[882][3] ), .D(\registers[883][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2301) );
  MX4X1 U6517 ( .A(\registers[864][3] ), .B(\registers[865][3] ), .C(
        \registers[866][3] ), .D(\registers[867][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2307) );
  MX4X1 U6518 ( .A(\registers[768][3] ), .B(\registers[769][3] ), .C(
        \registers[770][3] ), .D(\registers[771][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2343) );
  MX4X1 U6519 ( .A(\registers[816][3] ), .B(\registers[817][3] ), .C(
        \registers[818][3] ), .D(\registers[819][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2323) );
  MX4X1 U6520 ( .A(\registers[800][3] ), .B(\registers[801][3] ), .C(
        \registers[802][3] ), .D(\registers[803][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2328) );
  MX4X1 U6521 ( .A(\registers[960][3] ), .B(\registers[961][3] ), .C(
        \registers[962][3] ), .D(\registers[963][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2274) );
  MX4X1 U6522 ( .A(\registers[1008][3] ), .B(\registers[1009][3] ), .C(
        \registers[1010][3] ), .D(\registers[1011][3] ), .S0(n4168), .S1(n4405), .Y(n2258) );
  MX4X1 U6523 ( .A(\registers[992][3] ), .B(\registers[993][3] ), .C(
        \registers[994][3] ), .D(\registers[995][3] ), .S0(n4168), .S1(n4406), 
        .Y(n2263) );
  MX4X1 U6524 ( .A(\registers[896][3] ), .B(\registers[897][3] ), .C(
        \registers[898][3] ), .D(\registers[899][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2295) );
  MX4X1 U6525 ( .A(\registers[944][3] ), .B(\registers[945][3] ), .C(
        \registers[946][3] ), .D(\registers[947][3] ), .S0(n4169), .S1(n4407), 
        .Y(n2280) );
  MX4X1 U6526 ( .A(\registers[928][3] ), .B(\registers[929][3] ), .C(
        \registers[930][3] ), .D(\registers[931][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2285) );
  MX4X1 U6527 ( .A(\registers[576][3] ), .B(\registers[577][3] ), .C(
        \registers[578][3] ), .D(\registers[579][3] ), .S0(n4177), .S1(n4414), 
        .Y(n2470) );
  MX4X1 U6528 ( .A(\registers[624][3] ), .B(\registers[625][3] ), .C(
        \registers[626][3] ), .D(\registers[627][3] ), .S0(n4176), .S1(n4413), 
        .Y(n2455) );
  MX4X1 U6529 ( .A(\registers[608][3] ), .B(\registers[609][3] ), .C(
        \registers[610][3] ), .D(\registers[611][3] ), .S0(n4176), .S1(n4413), 
        .Y(n2460) );
  MX4X1 U6530 ( .A(\registers[512][3] ), .B(\registers[513][3] ), .C(
        \registers[514][3] ), .D(\registers[515][3] ), .S0(n4178), .S1(n4415), 
        .Y(n2491) );
  MX4X1 U6531 ( .A(\registers[560][3] ), .B(\registers[561][3] ), .C(
        \registers[562][3] ), .D(\registers[563][3] ), .S0(n4177), .S1(n4414), 
        .Y(n2476) );
  MX4X1 U6532 ( .A(\registers[544][3] ), .B(\registers[545][3] ), .C(
        \registers[546][3] ), .D(\registers[547][3] ), .S0(n4178), .S1(n4414), 
        .Y(n2481) );
  MX4X1 U6533 ( .A(\registers[704][3] ), .B(\registers[705][3] ), .C(
        \registers[706][3] ), .D(\registers[707][3] ), .S0(n4174), .S1(n4411), 
        .Y(n2373) );
  MX4X1 U6534 ( .A(\registers[752][3] ), .B(\registers[753][3] ), .C(
        \registers[754][3] ), .D(\registers[755][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2356) );
  MX4X1 U6535 ( .A(\registers[736][3] ), .B(\registers[737][3] ), .C(
        \registers[738][3] ), .D(\registers[739][3] ), .S0(n4174), .S1(n4411), 
        .Y(n2361) );
  MX4X1 U6536 ( .A(\registers[640][3] ), .B(\registers[641][3] ), .C(
        \registers[642][3] ), .D(\registers[643][3] ), .S0(n4176), .S1(n4412), 
        .Y(n2449) );
  MX4X1 U6537 ( .A(\registers[688][3] ), .B(\registers[689][3] ), .C(
        \registers[690][3] ), .D(\registers[691][3] ), .S0(n4175), .S1(n4411), 
        .Y(n2379) );
  MX4X1 U6538 ( .A(\registers[672][3] ), .B(\registers[673][3] ), .C(
        \registers[674][3] ), .D(\registers[675][3] ), .S0(n4175), .S1(n4412), 
        .Y(n2439) );
  MX4X1 U6539 ( .A(\registers[320][4] ), .B(\registers[321][4] ), .C(
        \registers[322][4] ), .D(\registers[323][4] ), .S0(n4204), .S1(n4438), 
        .Y(n2895) );
  MX4X1 U6540 ( .A(\registers[368][4] ), .B(\registers[369][4] ), .C(
        \registers[370][4] ), .D(\registers[371][4] ), .S0(n4203), .S1(n4437), 
        .Y(n2880) );
  MX4X1 U6541 ( .A(\registers[352][4] ), .B(\registers[353][4] ), .C(
        \registers[354][4] ), .D(\registers[355][4] ), .S0(n4203), .S1(n4438), 
        .Y(n2885) );
  MX4X1 U6542 ( .A(\registers[64][4] ), .B(\registers[65][4] ), .C(
        \registers[66][4] ), .D(\registers[67][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2980) );
  MX4X1 U6543 ( .A(\registers[112][4] ), .B(\registers[113][4] ), .C(
        \registers[114][4] ), .D(\registers[115][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2965) );
  MX4X1 U6544 ( .A(\registers[96][4] ), .B(\registers[97][4] ), .C(
        \registers[98][4] ), .D(\registers[99][4] ), .S0(n4208), .S1(n4443), 
        .Y(n2970) );
  MX4X1 U6545 ( .A(\registers[0][4] ), .B(\registers[1][4] ), .C(
        \registers[2][4] ), .D(\registers[3][4] ), .S0(n4210), .S1(n4444), .Y(
        n3001) );
  MX4X1 U6546 ( .A(\registers[48][4] ), .B(\registers[49][4] ), .C(
        \registers[50][4] ), .D(\registers[51][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2986) );
  MX4X1 U6547 ( .A(\registers[32][4] ), .B(\registers[33][4] ), .C(
        \registers[34][4] ), .D(\registers[35][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2991) );
  MX4X1 U6548 ( .A(\registers[192][4] ), .B(\registers[193][4] ), .C(
        \registers[194][4] ), .D(\registers[195][4] ), .S0(n4206), .S1(n4441), 
        .Y(n2938) );
  MX4X1 U6549 ( .A(\registers[240][4] ), .B(\registers[241][4] ), .C(
        \registers[242][4] ), .D(\registers[243][4] ), .S0(n4205), .S1(n4440), 
        .Y(n2923) );
  MX4X1 U6550 ( .A(\registers[224][4] ), .B(\registers[225][4] ), .C(
        \registers[226][4] ), .D(\registers[227][4] ), .S0(n4206), .S1(n4440), 
        .Y(n2928) );
  MX4X1 U6551 ( .A(\registers[128][4] ), .B(\registers[129][4] ), .C(
        \registers[130][4] ), .D(\registers[131][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2959) );
  MX4X1 U6552 ( .A(\registers[176][4] ), .B(\registers[177][4] ), .C(
        \registers[178][4] ), .D(\registers[179][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2944) );
  MX4X1 U6553 ( .A(\registers[160][4] ), .B(\registers[161][4] ), .C(
        \registers[162][4] ), .D(\registers[163][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2949) );
  MX4X1 U6554 ( .A(\registers[832][4] ), .B(\registers[833][4] ), .C(
        \registers[834][4] ), .D(\registers[835][4] ), .S0(n4193), .S1(n4428), 
        .Y(n2725) );
  MX4X1 U6555 ( .A(\registers[880][4] ), .B(\registers[881][4] ), .C(
        \registers[882][4] ), .D(\registers[883][4] ), .S0(n4192), .S1(n4427), 
        .Y(n2710) );
  MX4X1 U6556 ( .A(\registers[864][4] ), .B(\registers[865][4] ), .C(
        \registers[866][4] ), .D(\registers[867][4] ), .S0(n4192), .S1(n4428), 
        .Y(n2715) );
  MX4X1 U6557 ( .A(\registers[768][4] ), .B(\registers[769][4] ), .C(
        \registers[770][4] ), .D(\registers[771][4] ), .S0(n4194), .S1(n4430), 
        .Y(n2746) );
  MX4X1 U6558 ( .A(\registers[816][4] ), .B(\registers[817][4] ), .C(
        \registers[818][4] ), .D(\registers[819][4] ), .S0(n4193), .S1(n4429), 
        .Y(n2731) );
  MX4X1 U6559 ( .A(\registers[800][4] ), .B(\registers[801][4] ), .C(
        \registers[802][4] ), .D(\registers[803][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2736) );
  MX4X1 U6560 ( .A(\registers[960][4] ), .B(\registers[961][4] ), .C(
        \registers[962][4] ), .D(\registers[963][4] ), .S0(n4190), .S1(n4426), 
        .Y(n2683) );
  MX4X1 U6561 ( .A(\registers[1008][4] ), .B(\registers[1009][4] ), .C(
        \registers[1010][4] ), .D(\registers[1011][4] ), .S0(n4189), .S1(n4425), .Y(n2668) );
  MX4X1 U6562 ( .A(\registers[992][4] ), .B(\registers[993][4] ), .C(
        \registers[994][4] ), .D(\registers[995][4] ), .S0(n4190), .S1(n4425), 
        .Y(n2673) );
  MX4X1 U6563 ( .A(\registers[896][4] ), .B(\registers[897][4] ), .C(
        \registers[898][4] ), .D(\registers[899][4] ), .S0(n4192), .S1(n4427), 
        .Y(n2704) );
  MX4X1 U6564 ( .A(\registers[944][4] ), .B(\registers[945][4] ), .C(
        \registers[946][4] ), .D(\registers[947][4] ), .S0(n4191), .S1(n4426), 
        .Y(n2689) );
  MX4X1 U6565 ( .A(\registers[928][4] ), .B(\registers[929][4] ), .C(
        \registers[930][4] ), .D(\registers[931][4] ), .S0(n4191), .S1(n4427), 
        .Y(n2694) );
  MX4X1 U6566 ( .A(\registers[576][4] ), .B(\registers[577][4] ), .C(
        \registers[578][4] ), .D(\registers[579][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2810) );
  MX4X1 U6567 ( .A(\registers[624][4] ), .B(\registers[625][4] ), .C(
        \registers[626][4] ), .D(\registers[627][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2795) );
  MX4X1 U6568 ( .A(\registers[608][4] ), .B(\registers[609][4] ), .C(
        \registers[610][4] ), .D(\registers[611][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2800) );
  MX4X1 U6569 ( .A(\registers[512][4] ), .B(\registers[513][4] ), .C(
        \registers[514][4] ), .D(\registers[515][4] ), .S0(n4200), .S1(n4435), 
        .Y(n2831) );
  MX4X1 U6570 ( .A(\registers[560][4] ), .B(\registers[561][4] ), .C(
        \registers[562][4] ), .D(\registers[563][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2816) );
  MX4X1 U6571 ( .A(\registers[544][4] ), .B(\registers[545][4] ), .C(
        \registers[546][4] ), .D(\registers[547][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2821) );
  MX4X1 U6572 ( .A(\registers[704][4] ), .B(\registers[705][4] ), .C(
        \registers[706][4] ), .D(\registers[707][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2768) );
  MX4X1 U6573 ( .A(\registers[752][4] ), .B(\registers[753][4] ), .C(
        \registers[754][4] ), .D(\registers[755][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2753) );
  MX4X1 U6574 ( .A(\registers[736][4] ), .B(\registers[737][4] ), .C(
        \registers[738][4] ), .D(\registers[739][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2758) );
  MX4X1 U6575 ( .A(\registers[640][4] ), .B(\registers[641][4] ), .C(
        \registers[642][4] ), .D(\registers[643][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2789) );
  MX4X1 U6576 ( .A(\registers[688][4] ), .B(\registers[689][4] ), .C(
        \registers[690][4] ), .D(\registers[691][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2774) );
  MX4X1 U6577 ( .A(\registers[672][4] ), .B(\registers[673][4] ), .C(
        \registers[674][4] ), .D(\registers[675][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2779) );
  MX4X1 U6578 ( .A(\registers[320][5] ), .B(\registers[321][5] ), .C(
        \registers[322][5] ), .D(\registers[323][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3235) );
  MX4X1 U6579 ( .A(\registers[368][5] ), .B(\registers[369][5] ), .C(
        \registers[370][5] ), .D(\registers[371][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3220) );
  MX4X1 U6580 ( .A(\registers[352][5] ), .B(\registers[353][5] ), .C(
        \registers[354][5] ), .D(\registers[355][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3225) );
  MX4X1 U6581 ( .A(\registers[64][5] ), .B(\registers[65][5] ), .C(
        \registers[66][5] ), .D(\registers[67][5] ), .S0(n4230), .S1(n4463), 
        .Y(n3320) );
  MX4X1 U6582 ( .A(\registers[112][5] ), .B(\registers[113][5] ), .C(
        \registers[114][5] ), .D(\registers[115][5] ), .S0(n4229), .S1(n4462), 
        .Y(n3305) );
  MX4X1 U6583 ( .A(\registers[96][5] ), .B(\registers[97][5] ), .C(
        \registers[98][5] ), .D(\registers[99][5] ), .S0(n4230), .S1(n4462), 
        .Y(n3310) );
  MX4X1 U6584 ( .A(\registers[0][5] ), .B(\registers[1][5] ), .C(
        \registers[2][5] ), .D(\registers[3][5] ), .S0(n4232), .S1(n4464), .Y(
        n3341) );
  MX4X1 U6585 ( .A(\registers[48][5] ), .B(\registers[49][5] ), .C(
        \registers[50][5] ), .D(\registers[51][5] ), .S0(n4231), .S1(n4463), 
        .Y(n3326) );
  MX4X1 U6586 ( .A(\registers[32][5] ), .B(\registers[33][5] ), .C(
        \registers[34][5] ), .D(\registers[35][5] ), .S0(n4231), .S1(n4463), 
        .Y(n3331) );
  MX4X1 U6587 ( .A(\registers[192][5] ), .B(\registers[193][5] ), .C(
        \registers[194][5] ), .D(\registers[195][5] ), .S0(n4228), .S1(n4460), 
        .Y(n3278) );
  MX4X1 U6588 ( .A(\registers[240][5] ), .B(\registers[241][5] ), .C(
        \registers[242][5] ), .D(\registers[243][5] ), .S0(n4227), .S1(n4459), 
        .Y(n3263) );
  MX4X1 U6589 ( .A(\registers[224][5] ), .B(\registers[225][5] ), .C(
        \registers[226][5] ), .D(\registers[227][5] ), .S0(n4227), .S1(n4460), 
        .Y(n3268) );
  MX4X1 U6590 ( .A(\registers[128][5] ), .B(\registers[129][5] ), .C(
        \registers[130][5] ), .D(\registers[131][5] ), .S0(n4229), .S1(n4462), 
        .Y(n3299) );
  MX4X1 U6591 ( .A(\registers[176][5] ), .B(\registers[177][5] ), .C(
        \registers[178][5] ), .D(\registers[179][5] ), .S0(n4228), .S1(n4461), 
        .Y(n3284) );
  MX4X1 U6592 ( .A(\registers[160][5] ), .B(\registers[161][5] ), .C(
        \registers[162][5] ), .D(\registers[163][5] ), .S0(n4228), .S1(n4461), 
        .Y(n3289) );
  MX4X1 U6593 ( .A(\registers[832][5] ), .B(\registers[833][5] ), .C(
        \registers[834][5] ), .D(\registers[835][5] ), .S0(n4214), .S1(n4448), 
        .Y(n3065) );
  MX4X1 U6594 ( .A(\registers[880][5] ), .B(\registers[881][5] ), .C(
        \registers[882][5] ), .D(\registers[883][5] ), .S0(n4213), .S1(n4447), 
        .Y(n3050) );
  MX4X1 U6595 ( .A(\registers[864][5] ), .B(\registers[865][5] ), .C(
        \registers[866][5] ), .D(\registers[867][5] ), .S0(n4214), .S1(n4447), 
        .Y(n3055) );
  MX4X1 U6596 ( .A(\registers[768][5] ), .B(\registers[769][5] ), .C(
        \registers[770][5] ), .D(\registers[771][5] ), .S0(n4216), .S1(n4449), 
        .Y(n3086) );
  MX4X1 U6597 ( .A(\registers[816][5] ), .B(\registers[817][5] ), .C(
        \registers[818][5] ), .D(\registers[819][5] ), .S0(n4215), .S1(n4448), 
        .Y(n3071) );
  MX4X1 U6598 ( .A(\registers[800][5] ), .B(\registers[801][5] ), .C(
        \registers[802][5] ), .D(\registers[803][5] ), .S0(n4215), .S1(n4449), 
        .Y(n3076) );
  MX4X1 U6599 ( .A(\registers[960][5] ), .B(\registers[961][5] ), .C(
        \registers[962][5] ), .D(\registers[963][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3023) );
  MX4X1 U6600 ( .A(\registers[1008][5] ), .B(\registers[1009][5] ), .C(
        \registers[1010][5] ), .D(\registers[1011][5] ), .S0(n4211), .S1(n4445), .Y(n3008) );
  MX4X1 U6601 ( .A(\registers[992][5] ), .B(\registers[993][5] ), .C(
        \registers[994][5] ), .D(\registers[995][5] ), .S0(n4211), .S1(n4445), 
        .Y(n3013) );
  MX4X1 U6602 ( .A(\registers[896][5] ), .B(\registers[897][5] ), .C(
        \registers[898][5] ), .D(\registers[899][5] ), .S0(n4213), .S1(n4447), 
        .Y(n3044) );
  MX4X1 U6603 ( .A(\registers[944][5] ), .B(\registers[945][5] ), .C(
        \registers[946][5] ), .D(\registers[947][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3029) );
  MX4X1 U6604 ( .A(\registers[928][5] ), .B(\registers[929][5] ), .C(
        \registers[930][5] ), .D(\registers[931][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3034) );
  MX4X1 U6605 ( .A(\registers[576][5] ), .B(\registers[577][5] ), .C(
        \registers[578][5] ), .D(\registers[579][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3150) );
  MX4X1 U6606 ( .A(\registers[624][5] ), .B(\registers[625][5] ), .C(
        \registers[626][5] ), .D(\registers[627][5] ), .S0(n4219), .S1(n4452), 
        .Y(n3135) );
  MX4X1 U6607 ( .A(\registers[608][5] ), .B(\registers[609][5] ), .C(
        \registers[610][5] ), .D(\registers[611][5] ), .S0(n4219), .S1(n4452), 
        .Y(n3140) );
  MX4X1 U6608 ( .A(\registers[512][5] ), .B(\registers[513][5] ), .C(
        \registers[514][5] ), .D(\registers[515][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3171) );
  MX4X1 U6609 ( .A(\registers[560][5] ), .B(\registers[561][5] ), .C(
        \registers[562][5] ), .D(\registers[563][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3156) );
  MX4X1 U6610 ( .A(\registers[544][5] ), .B(\registers[545][5] ), .C(
        \registers[546][5] ), .D(\registers[547][5] ), .S0(n4220), .S1(n4454), 
        .Y(n3161) );
  MX4X1 U6611 ( .A(\registers[704][5] ), .B(\registers[705][5] ), .C(
        \registers[706][5] ), .D(\registers[707][5] ), .S0(n4217), .S1(n4451), 
        .Y(n3108) );
  MX4X1 U6612 ( .A(\registers[752][5] ), .B(\registers[753][5] ), .C(
        \registers[754][5] ), .D(\registers[755][5] ), .S0(n4216), .S1(n4450), 
        .Y(n3093) );
  MX4X1 U6613 ( .A(\registers[736][5] ), .B(\registers[737][5] ), .C(
        \registers[738][5] ), .D(\registers[739][5] ), .S0(n4216), .S1(n4450), 
        .Y(n3098) );
  MX4X1 U6614 ( .A(\registers[640][5] ), .B(\registers[641][5] ), .C(
        \registers[642][5] ), .D(\registers[643][5] ), .S0(n4218), .S1(n4452), 
        .Y(n3129) );
  MX4X1 U6615 ( .A(\registers[688][5] ), .B(\registers[689][5] ), .C(
        \registers[690][5] ), .D(\registers[691][5] ), .S0(n4217), .S1(n4451), 
        .Y(n3114) );
  MX4X1 U6616 ( .A(\registers[672][5] ), .B(\registers[673][5] ), .C(
        \registers[674][5] ), .D(\registers[675][5] ), .S0(n4218), .S1(n4451), 
        .Y(n3119) );
  MX4X1 U6617 ( .A(\registers[320][6] ), .B(\registers[321][6] ), .C(
        \registers[322][6] ), .D(\registers[323][6] ), .S0(n4246), .S1(n4478), 
        .Y(n3575) );
  MX4X1 U6618 ( .A(\registers[368][6] ), .B(\registers[369][6] ), .C(
        \registers[370][6] ), .D(\registers[371][6] ), .S0(n4245), .S1(n4477), 
        .Y(n3560) );
  MX4X1 U6619 ( .A(\registers[352][6] ), .B(\registers[353][6] ), .C(
        \registers[354][6] ), .D(\registers[355][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3565) );
  MX4X1 U6620 ( .A(\registers[64][6] ), .B(\registers[65][6] ), .C(
        \registers[66][6] ), .D(\registers[67][6] ), .S0(n4252), .S1(n4483), 
        .Y(n3660) );
  MX4X1 U6621 ( .A(\registers[112][6] ), .B(\registers[113][6] ), .C(
        \registers[114][6] ), .D(\registers[115][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3645) );
  MX4X1 U6622 ( .A(\registers[96][6] ), .B(\registers[97][6] ), .C(
        \registers[98][6] ), .D(\registers[99][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3650) );
  MX4X1 U6623 ( .A(\registers[0][6] ), .B(\registers[1][6] ), .C(
        \registers[2][6] ), .D(\registers[3][6] ), .S0(n4253), .S1(n4484), .Y(
        n3681) );
  MX4X1 U6624 ( .A(\registers[48][6] ), .B(\registers[49][6] ), .C(
        \registers[50][6] ), .D(\registers[51][6] ), .S0(n4252), .S1(n4483), 
        .Y(n3666) );
  MX4X1 U6625 ( .A(\registers[32][6] ), .B(\registers[33][6] ), .C(
        \registers[34][6] ), .D(\registers[35][6] ), .S0(n4252), .S1(n4483), 
        .Y(n3671) );
  MX4X1 U6626 ( .A(\registers[192][6] ), .B(\registers[193][6] ), .C(
        \registers[194][6] ), .D(\registers[195][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3618) );
  MX4X1 U6627 ( .A(\registers[240][6] ), .B(\registers[241][6] ), .C(
        \registers[242][6] ), .D(\registers[243][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3603) );
  MX4X1 U6628 ( .A(\registers[224][6] ), .B(\registers[225][6] ), .C(
        \registers[226][6] ), .D(\registers[227][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3608) );
  MX4X1 U6629 ( .A(\registers[128][6] ), .B(\registers[129][6] ), .C(
        \registers[130][6] ), .D(\registers[131][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3639) );
  MX4X1 U6630 ( .A(\registers[176][6] ), .B(\registers[177][6] ), .C(
        \registers[178][6] ), .D(\registers[179][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3624) );
  MX4X1 U6631 ( .A(\registers[160][6] ), .B(\registers[161][6] ), .C(
        \registers[162][6] ), .D(\registers[163][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3629) );
  MX4X1 U6632 ( .A(\registers[832][6] ), .B(\registers[833][6] ), .C(
        \registers[834][6] ), .D(\registers[835][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3405) );
  MX4X1 U6633 ( .A(\registers[880][6] ), .B(\registers[881][6] ), .C(
        \registers[882][6] ), .D(\registers[883][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3390) );
  MX4X1 U6634 ( .A(\registers[864][6] ), .B(\registers[865][6] ), .C(
        \registers[866][6] ), .D(\registers[867][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3395) );
  MX4X1 U6635 ( .A(\registers[768][6] ), .B(\registers[769][6] ), .C(
        \registers[770][6] ), .D(\registers[771][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3426) );
  MX4X1 U6636 ( .A(\registers[816][6] ), .B(\registers[817][6] ), .C(
        \registers[818][6] ), .D(\registers[819][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3411) );
  MX4X1 U6637 ( .A(\registers[800][6] ), .B(\registers[801][6] ), .C(
        \registers[802][6] ), .D(\registers[803][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3416) );
  MX4X1 U6638 ( .A(\registers[960][6] ), .B(\registers[961][6] ), .C(
        \registers[962][6] ), .D(\registers[963][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3363) );
  MX4X1 U6639 ( .A(\registers[1008][6] ), .B(\registers[1009][6] ), .C(
        \registers[1010][6] ), .D(\registers[1011][6] ), .S0(n4232), .S1(n4464), .Y(n3348) );
  MX4X1 U6640 ( .A(\registers[992][6] ), .B(\registers[993][6] ), .C(
        \registers[994][6] ), .D(\registers[995][6] ), .S0(n4232), .S1(n4465), 
        .Y(n3353) );
  MX4X1 U6641 ( .A(\registers[896][6] ), .B(\registers[897][6] ), .C(
        \registers[898][6] ), .D(\registers[899][6] ), .S0(n4234), .S1(n4467), 
        .Y(n3384) );
  MX4X1 U6642 ( .A(\registers[944][6] ), .B(\registers[945][6] ), .C(
        \registers[946][6] ), .D(\registers[947][6] ), .S0(n4233), .S1(n4466), 
        .Y(n3369) );
  MX4X1 U6643 ( .A(\registers[928][6] ), .B(\registers[929][6] ), .C(
        \registers[930][6] ), .D(\registers[931][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3374) );
  MX4X1 U6644 ( .A(\registers[576][6] ), .B(\registers[577][6] ), .C(
        \registers[578][6] ), .D(\registers[579][6] ), .S0(n4241), .S1(n4473), 
        .Y(n3490) );
  MX4X1 U6645 ( .A(\registers[624][6] ), .B(\registers[625][6] ), .C(
        \registers[626][6] ), .D(\registers[627][6] ), .S0(n4240), .S1(n4472), 
        .Y(n3475) );
  MX4X1 U6646 ( .A(\registers[608][6] ), .B(\registers[609][6] ), .C(
        \registers[610][6] ), .D(\registers[611][6] ), .S0(n4240), .S1(n4472), 
        .Y(n3480) );
  MX4X1 U6647 ( .A(\registers[512][6] ), .B(\registers[513][6] ), .C(
        \registers[514][6] ), .D(\registers[515][6] ), .S0(n4242), .S1(n4474), 
        .Y(n3511) );
  MX4X1 U6648 ( .A(\registers[560][6] ), .B(\registers[561][6] ), .C(
        \registers[562][6] ), .D(\registers[563][6] ), .S0(n4241), .S1(n4473), 
        .Y(n3496) );
  MX4X1 U6649 ( .A(\registers[544][6] ), .B(\registers[545][6] ), .C(
        \registers[546][6] ), .D(\registers[547][6] ), .S0(n4242), .S1(n4473), 
        .Y(n3501) );
  MX4X1 U6650 ( .A(\registers[704][6] ), .B(\registers[705][6] ), .C(
        \registers[706][6] ), .D(\registers[707][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3448) );
  MX4X1 U6651 ( .A(\registers[752][6] ), .B(\registers[753][6] ), .C(
        \registers[754][6] ), .D(\registers[755][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3433) );
  MX4X1 U6652 ( .A(\registers[736][6] ), .B(\registers[737][6] ), .C(
        \registers[738][6] ), .D(\registers[739][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3438) );
  MX4X1 U6653 ( .A(\registers[640][6] ), .B(\registers[641][6] ), .C(
        \registers[642][6] ), .D(\registers[643][6] ), .S0(n4240), .S1(n4471), 
        .Y(n3469) );
  MX4X1 U6654 ( .A(\registers[688][6] ), .B(\registers[689][6] ), .C(
        \registers[690][6] ), .D(\registers[691][6] ), .S0(n4239), .S1(n4471), 
        .Y(n3454) );
  MX4X1 U6655 ( .A(\registers[672][6] ), .B(\registers[673][6] ), .C(
        \registers[674][6] ), .D(\registers[675][6] ), .S0(n4239), .S1(n4471), 
        .Y(n3459) );
  MX4X1 U6656 ( .A(\registers[320][7] ), .B(\registers[321][7] ), .C(
        \registers[322][7] ), .D(\registers[323][7] ), .S0(n4268), .S1(n4490), 
        .Y(n3915) );
  MX4X1 U6657 ( .A(\registers[368][7] ), .B(\registers[369][7] ), .C(
        \registers[370][7] ), .D(\registers[371][7] ), .S0(n4267), .S1(n4496), 
        .Y(n3900) );
  MX4X1 U6658 ( .A(\registers[352][7] ), .B(\registers[353][7] ), .C(
        \registers[354][7] ), .D(\registers[355][7] ), .S0(n4267), .S1(n4472), 
        .Y(n3905) );
  MX4X1 U6659 ( .A(\registers[64][7] ), .B(\registers[65][7] ), .C(
        \registers[66][7] ), .D(\registers[67][7] ), .S0(n4273), .S1(n4299), 
        .Y(n4000) );
  MX4X1 U6660 ( .A(\registers[112][7] ), .B(\registers[113][7] ), .C(
        \registers[114][7] ), .D(\registers[115][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3985) );
  MX4X1 U6661 ( .A(\registers[96][7] ), .B(\registers[97][7] ), .C(
        \registers[98][7] ), .D(\registers[99][7] ), .S0(n4272), .S1(n4298), 
        .Y(n3990) );
  MX4X1 U6662 ( .A(\registers[0][7] ), .B(\registers[1][7] ), .C(
        \registers[2][7] ), .D(\registers[3][7] ), .S0(n4274), .S1(n4501), .Y(
        n4021) );
  MX4X1 U6663 ( .A(\registers[48][7] ), .B(\registers[49][7] ), .C(
        \registers[50][7] ), .D(\registers[51][7] ), .S0(n4273), .S1(n4501), 
        .Y(n4006) );
  MX4X1 U6664 ( .A(\registers[32][7] ), .B(\registers[33][7] ), .C(
        \registers[34][7] ), .D(\registers[35][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4011) );
  MX4X1 U6665 ( .A(\registers[192][7] ), .B(\registers[193][7] ), .C(
        \registers[194][7] ), .D(\registers[195][7] ), .S0(n4270), .S1(n4499), 
        .Y(n3958) );
  MX4X1 U6666 ( .A(\registers[240][7] ), .B(\registers[241][7] ), .C(
        \registers[242][7] ), .D(\registers[243][7] ), .S0(n4269), .S1(n4498), 
        .Y(n3943) );
  MX4X1 U6667 ( .A(\registers[224][7] ), .B(\registers[225][7] ), .C(
        \registers[226][7] ), .D(\registers[227][7] ), .S0(n4270), .S1(n4498), 
        .Y(n3948) );
  MX4X1 U6668 ( .A(\registers[128][7] ), .B(\registers[129][7] ), .C(
        \registers[130][7] ), .D(\registers[131][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3979) );
  MX4X1 U6669 ( .A(\registers[176][7] ), .B(\registers[177][7] ), .C(
        \registers[178][7] ), .D(\registers[179][7] ), .S0(n4271), .S1(n4499), 
        .Y(n3964) );
  MX4X1 U6670 ( .A(\registers[160][7] ), .B(\registers[161][7] ), .C(
        \registers[162][7] ), .D(\registers[163][7] ), .S0(n4271), .S1(n4499), 
        .Y(n3969) );
  MX4X1 U6671 ( .A(\registers[832][7] ), .B(\registers[833][7] ), .C(
        \registers[834][7] ), .D(\registers[835][7] ), .S0(n4257), .S1(n4487), 
        .Y(n3745) );
  MX4X1 U6672 ( .A(\registers[880][7] ), .B(\registers[881][7] ), .C(
        \registers[882][7] ), .D(\registers[883][7] ), .S0(n4256), .S1(n4487), 
        .Y(n3730) );
  MX4X1 U6673 ( .A(\registers[864][7] ), .B(\registers[865][7] ), .C(
        \registers[866][7] ), .D(\registers[867][7] ), .S0(n4256), .S1(n4487), 
        .Y(n3735) );
  MX4X1 U6674 ( .A(\registers[768][7] ), .B(\registers[769][7] ), .C(
        \registers[770][7] ), .D(\registers[771][7] ), .S0(n4258), .S1(n4489), 
        .Y(n3766) );
  MX4X1 U6675 ( .A(\registers[816][7] ), .B(\registers[817][7] ), .C(
        \registers[818][7] ), .D(\registers[819][7] ), .S0(n4257), .S1(n4488), 
        .Y(n3751) );
  MX4X1 U6676 ( .A(\registers[800][7] ), .B(\registers[801][7] ), .C(
        \registers[802][7] ), .D(\registers[803][7] ), .S0(n4258), .S1(n4488), 
        .Y(n3756) );
  MX4X1 U6677 ( .A(\registers[960][7] ), .B(\registers[961][7] ), .C(
        \registers[962][7] ), .D(\registers[963][7] ), .S0(n4254), .S1(n4485), 
        .Y(n3703) );
  MX4X1 U6678 ( .A(\registers[1008][7] ), .B(\registers[1009][7] ), .C(
        \registers[1010][7] ), .D(\registers[1011][7] ), .S0(n4253), .S1(n4484), .Y(n3688) );
  MX4X1 U6679 ( .A(\registers[992][7] ), .B(\registers[993][7] ), .C(
        \registers[994][7] ), .D(\registers[995][7] ), .S0(n4254), .S1(n4484), 
        .Y(n3693) );
  MX4X1 U6680 ( .A(\registers[896][7] ), .B(\registers[897][7] ), .C(
        \registers[898][7] ), .D(\registers[899][7] ), .S0(n4256), .S1(n4486), 
        .Y(n3724) );
  MX4X1 U6681 ( .A(\registers[944][7] ), .B(\registers[945][7] ), .C(
        \registers[946][7] ), .D(\registers[947][7] ), .S0(n4255), .S1(n4485), 
        .Y(n3709) );
  MX4X1 U6682 ( .A(\registers[928][7] ), .B(\registers[929][7] ), .C(
        \registers[930][7] ), .D(\registers[931][7] ), .S0(n4255), .S1(n4486), 
        .Y(n3714) );
  MX4X1 U6683 ( .A(\registers[576][7] ), .B(\registers[577][7] ), .C(
        \registers[578][7] ), .D(\registers[579][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3830) );
  MX4X1 U6684 ( .A(\registers[624][7] ), .B(\registers[625][7] ), .C(
        \registers[626][7] ), .D(\registers[627][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3815) );
  MX4X1 U6685 ( .A(\registers[608][7] ), .B(\registers[609][7] ), .C(
        \registers[610][7] ), .D(\registers[611][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3820) );
  MX4X1 U6686 ( .A(\registers[512][7] ), .B(\registers[513][7] ), .C(
        \registers[514][7] ), .D(\registers[515][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3851) );
  MX4X1 U6687 ( .A(\registers[560][7] ), .B(\registers[561][7] ), .C(
        \registers[562][7] ), .D(\registers[563][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3836) );
  MX4X1 U6688 ( .A(\registers[544][7] ), .B(\registers[545][7] ), .C(
        \registers[546][7] ), .D(\registers[547][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3841) );
  MX4X1 U6689 ( .A(\registers[704][7] ), .B(\registers[705][7] ), .C(
        \registers[706][7] ), .D(\registers[707][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3788) );
  MX4X1 U6690 ( .A(\registers[752][7] ), .B(\registers[753][7] ), .C(
        \registers[754][7] ), .D(\registers[755][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3773) );
  MX4X1 U6691 ( .A(\registers[736][7] ), .B(\registers[737][7] ), .C(
        \registers[738][7] ), .D(\registers[739][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3778) );
  MX4X1 U6692 ( .A(\registers[640][7] ), .B(\registers[641][7] ), .C(
        \registers[642][7] ), .D(\registers[643][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3809) );
  MX4X1 U6693 ( .A(\registers[688][7] ), .B(\registers[689][7] ), .C(
        \registers[690][7] ), .D(\registers[691][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3794) );
  MX4X1 U6694 ( .A(\registers[672][7] ), .B(\registers[673][7] ), .C(
        \registers[674][7] ), .D(\registers[675][7] ), .S0(n4260), .S1(n4491), 
        .Y(n3799) );
  MX4X1 U6695 ( .A(\registers[320][0] ), .B(\registers[321][0] ), .C(
        \registers[322][0] ), .D(\registers[323][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4880) );
  MX4X1 U6696 ( .A(\registers[368][0] ), .B(\registers[369][0] ), .C(
        \registers[370][0] ), .D(\registers[371][0] ), .S0(n7460), .S1(n7703), 
        .Y(n4865) );
  MX4X1 U6697 ( .A(\registers[352][0] ), .B(\registers[353][0] ), .C(
        \registers[354][0] ), .D(\registers[355][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4870) );
  MX4X1 U6698 ( .A(\registers[64][0] ), .B(\registers[65][0] ), .C(
        \registers[66][0] ), .D(\registers[67][0] ), .S0(n7467), .S1(n7708), 
        .Y(n4965) );
  MX4X1 U6699 ( .A(\registers[112][0] ), .B(\registers[113][0] ), .C(
        \registers[114][0] ), .D(\registers[115][0] ), .S0(n7466), .S1(n7707), 
        .Y(n4950) );
  MX4X1 U6700 ( .A(\registers[96][0] ), .B(\registers[97][0] ), .C(
        \registers[98][0] ), .D(\registers[99][0] ), .S0(n7466), .S1(n7708), 
        .Y(n4955) );
  MX4X1 U6701 ( .A(\registers[0][0] ), .B(\registers[1][0] ), .C(
        \registers[2][0] ), .D(\registers[3][0] ), .S0(n7468), .S1(n7710), .Y(
        n4986) );
  MX4X1 U6702 ( .A(\registers[48][0] ), .B(\registers[49][0] ), .C(
        \registers[50][0] ), .D(\registers[51][0] ), .S0(n7467), .S1(n7709), 
        .Y(n4971) );
  MX4X1 U6703 ( .A(\registers[32][0] ), .B(\registers[33][0] ), .C(
        \registers[34][0] ), .D(\registers[35][0] ), .S0(n7467), .S1(n7709), 
        .Y(n4976) );
  MX4X1 U6704 ( .A(\registers[192][0] ), .B(\registers[193][0] ), .C(
        \registers[194][0] ), .D(\registers[195][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4923) );
  MX4X1 U6705 ( .A(\registers[240][0] ), .B(\registers[241][0] ), .C(
        \registers[242][0] ), .D(\registers[243][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4908) );
  MX4X1 U6706 ( .A(\registers[224][0] ), .B(\registers[225][0] ), .C(
        \registers[226][0] ), .D(\registers[227][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4913) );
  MX4X1 U6707 ( .A(\registers[128][0] ), .B(\registers[129][0] ), .C(
        \registers[130][0] ), .D(\registers[131][0] ), .S0(n7465), .S1(n7707), 
        .Y(n4944) );
  MX4X1 U6708 ( .A(\registers[176][0] ), .B(\registers[177][0] ), .C(
        \registers[178][0] ), .D(\registers[179][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4929) );
  MX4X1 U6709 ( .A(\registers[160][0] ), .B(\registers[161][0] ), .C(
        \registers[162][0] ), .D(\registers[163][0] ), .S0(n7465), .S1(n7707), 
        .Y(n4934) );
  MX4X1 U6710 ( .A(\registers[832][0] ), .B(\registers[833][0] ), .C(
        \registers[834][0] ), .D(\registers[835][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4710) );
  MX4X1 U6711 ( .A(\registers[880][0] ), .B(\registers[881][0] ), .C(
        \registers[882][0] ), .D(\registers[883][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4695) );
  MX4X1 U6712 ( .A(\registers[864][0] ), .B(\registers[865][0] ), .C(
        \registers[866][0] ), .D(\registers[867][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4700) );
  MX4X1 U6713 ( .A(\registers[768][0] ), .B(\registers[769][0] ), .C(
        \registers[770][0] ), .D(\registers[771][0] ), .S0(n7452), .S1(n7695), 
        .Y(n4731) );
  MX4X1 U6714 ( .A(\registers[816][0] ), .B(\registers[817][0] ), .C(
        \registers[818][0] ), .D(\registers[819][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4716) );
  MX4X1 U6715 ( .A(\registers[800][0] ), .B(\registers[801][0] ), .C(
        \registers[802][0] ), .D(\registers[803][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4721) );
  MX4X1 U6716 ( .A(\registers[960][0] ), .B(\registers[961][0] ), .C(
        \registers[962][0] ), .D(\registers[963][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4668) );
  MX4X1 U6717 ( .A(\registers[896][0] ), .B(\registers[897][0] ), .C(
        \registers[898][0] ), .D(\registers[899][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4689) );
  MX4X1 U6718 ( .A(\registers[944][0] ), .B(\registers[945][0] ), .C(
        \registers[946][0] ), .D(\registers[947][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4674) );
  MX4X1 U6719 ( .A(\registers[928][0] ), .B(\registers[929][0] ), .C(
        \registers[930][0] ), .D(\registers[931][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4679) );
  MX4X1 U6720 ( .A(\registers[576][0] ), .B(\registers[577][0] ), .C(
        \registers[578][0] ), .D(\registers[579][0] ), .S0(n7456), .S1(n7699), 
        .Y(n4795) );
  MX4X1 U6721 ( .A(\registers[624][0] ), .B(\registers[625][0] ), .C(
        \registers[626][0] ), .D(\registers[627][0] ), .S0(n7455), .S1(n7698), 
        .Y(n4780) );
  MX4X1 U6722 ( .A(\registers[608][0] ), .B(\registers[609][0] ), .C(
        \registers[610][0] ), .D(\registers[611][0] ), .S0(n7455), .S1(n7698), 
        .Y(n4785) );
  MX4X1 U6723 ( .A(\registers[512][0] ), .B(\registers[513][0] ), .C(
        \registers[514][0] ), .D(\registers[515][0] ), .S0(n7457), .S1(n7700), 
        .Y(n4816) );
  MX4X1 U6724 ( .A(\registers[560][0] ), .B(\registers[561][0] ), .C(
        \registers[562][0] ), .D(\registers[563][0] ), .S0(n7456), .S1(n7699), 
        .Y(n4801) );
  MX4X1 U6725 ( .A(\registers[544][0] ), .B(\registers[545][0] ), .C(
        \registers[546][0] ), .D(\registers[547][0] ), .S0(n7457), .S1(n7699), 
        .Y(n4806) );
  MX4X1 U6726 ( .A(\registers[704][0] ), .B(\registers[705][0] ), .C(
        \registers[706][0] ), .D(\registers[707][0] ), .S0(n7453), .S1(n7696), 
        .Y(n4753) );
  MX4X1 U6727 ( .A(\registers[752][0] ), .B(\registers[753][0] ), .C(
        \registers[754][0] ), .D(\registers[755][0] ), .S0(n7452), .S1(n7695), 
        .Y(n4738) );
  MX4X1 U6728 ( .A(\registers[736][0] ), .B(\registers[737][0] ), .C(
        \registers[738][0] ), .D(\registers[739][0] ), .S0(n7453), .S1(n7695), 
        .Y(n4743) );
  MX4X1 U6729 ( .A(\registers[640][0] ), .B(\registers[641][0] ), .C(
        \registers[642][0] ), .D(\registers[643][0] ), .S0(n7455), .S1(n7697), 
        .Y(n4774) );
  MX4X1 U6730 ( .A(\registers[688][0] ), .B(\registers[689][0] ), .C(
        \registers[690][0] ), .D(\registers[691][0] ), .S0(n7454), .S1(n7696), 
        .Y(n4759) );
  MX4X1 U6731 ( .A(\registers[672][0] ), .B(\registers[673][0] ), .C(
        \registers[674][0] ), .D(\registers[675][0] ), .S0(n7454), .S1(n7697), 
        .Y(n4764) );
  MX4X1 U6732 ( .A(\registers[320][1] ), .B(\registers[321][1] ), .C(
        \registers[322][1] ), .D(\registers[323][1] ), .S0(n7483), .S1(n7723), 
        .Y(n5220) );
  MX4X1 U6733 ( .A(\registers[368][1] ), .B(\registers[369][1] ), .C(
        \registers[370][1] ), .D(\registers[371][1] ), .S0(n7482), .S1(n7722), 
        .Y(n5205) );
  MX4X1 U6734 ( .A(\registers[352][1] ), .B(\registers[353][1] ), .C(
        \registers[354][1] ), .D(\registers[355][1] ), .S0(n7482), .S1(n7723), 
        .Y(n5210) );
  MX4X1 U6735 ( .A(\registers[64][1] ), .B(\registers[65][1] ), .C(
        \registers[66][1] ), .D(\registers[67][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5305) );
  MX4X1 U6736 ( .A(\registers[112][1] ), .B(\registers[113][1] ), .C(
        \registers[114][1] ), .D(\registers[115][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5290) );
  MX4X1 U6737 ( .A(\registers[96][1] ), .B(\registers[97][1] ), .C(
        \registers[98][1] ), .D(\registers[99][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5295) );
  MX4X1 U6738 ( .A(\registers[0][1] ), .B(\registers[1][1] ), .C(
        \registers[2][1] ), .D(\registers[3][1] ), .S0(n7489), .S1(n7729), .Y(
        n5326) );
  MX4X1 U6739 ( .A(\registers[48][1] ), .B(\registers[49][1] ), .C(
        \registers[50][1] ), .D(\registers[51][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5311) );
  MX4X1 U6740 ( .A(\registers[32][1] ), .B(\registers[33][1] ), .C(
        \registers[34][1] ), .D(\registers[35][1] ), .S0(n7489), .S1(n7729), 
        .Y(n5316) );
  MX4X1 U6741 ( .A(\registers[192][1] ), .B(\registers[193][1] ), .C(
        \registers[194][1] ), .D(\registers[195][1] ), .S0(n7485), .S1(n7726), 
        .Y(n5263) );
  MX4X1 U6742 ( .A(\registers[240][1] ), .B(\registers[241][1] ), .C(
        \registers[242][1] ), .D(\registers[243][1] ), .S0(n7484), .S1(n7725), 
        .Y(n5248) );
  MX4X1 U6743 ( .A(\registers[224][1] ), .B(\registers[225][1] ), .C(
        \registers[226][1] ), .D(\registers[227][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5253) );
  MX4X1 U6744 ( .A(\registers[128][1] ), .B(\registers[129][1] ), .C(
        \registers[130][1] ), .D(\registers[131][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5284) );
  MX4X1 U6745 ( .A(\registers[176][1] ), .B(\registers[177][1] ), .C(
        \registers[178][1] ), .D(\registers[179][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5269) );
  MX4X1 U6746 ( .A(\registers[160][1] ), .B(\registers[161][1] ), .C(
        \registers[162][1] ), .D(\registers[163][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5274) );
  MX4X1 U6747 ( .A(\registers[832][1] ), .B(\registers[833][1] ), .C(
        \registers[834][1] ), .D(\registers[835][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5050) );
  MX4X1 U6748 ( .A(\registers[880][1] ), .B(\registers[881][1] ), .C(
        \registers[882][1] ), .D(\registers[883][1] ), .S0(n7471), .S1(n7712), 
        .Y(n5035) );
  MX4X1 U6749 ( .A(\registers[864][1] ), .B(\registers[865][1] ), .C(
        \registers[866][1] ), .D(\registers[867][1] ), .S0(n7471), .S1(n7713), 
        .Y(n5040) );
  MX4X1 U6750 ( .A(\registers[768][1] ), .B(\registers[769][1] ), .C(
        \registers[770][1] ), .D(\registers[771][1] ), .S0(n7473), .S1(n7715), 
        .Y(n5071) );
  MX4X1 U6751 ( .A(\registers[816][1] ), .B(\registers[817][1] ), .C(
        \registers[818][1] ), .D(\registers[819][1] ), .S0(n7472), .S1(n7714), 
        .Y(n5056) );
  MX4X1 U6752 ( .A(\registers[800][1] ), .B(\registers[801][1] ), .C(
        \registers[802][1] ), .D(\registers[803][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5061) );
  MX4X1 U6753 ( .A(\registers[960][1] ), .B(\registers[961][1] ), .C(
        \registers[962][1] ), .D(\registers[963][1] ), .S0(n7469), .S1(n7711), 
        .Y(n5008) );
  MX4X1 U6754 ( .A(\registers[1008][1] ), .B(\registers[1009][1] ), .C(
        \registers[1010][1] ), .D(\registers[1011][1] ), .S0(n7468), .S1(n7710), .Y(n4993) );
  MX4X1 U6755 ( .A(\registers[992][1] ), .B(\registers[993][1] ), .C(
        \registers[994][1] ), .D(\registers[995][1] ), .S0(n7469), .S1(n7710), 
        .Y(n4998) );
  MX4X1 U6756 ( .A(\registers[896][1] ), .B(\registers[897][1] ), .C(
        \registers[898][1] ), .D(\registers[899][1] ), .S0(n7471), .S1(n7712), 
        .Y(n5029) );
  MX4X1 U6757 ( .A(\registers[944][1] ), .B(\registers[945][1] ), .C(
        \registers[946][1] ), .D(\registers[947][1] ), .S0(n7470), .S1(n7711), 
        .Y(n5014) );
  MX4X1 U6758 ( .A(\registers[928][1] ), .B(\registers[929][1] ), .C(
        \registers[930][1] ), .D(\registers[931][1] ), .S0(n7470), .S1(n7711), 
        .Y(n5019) );
  MX4X1 U6759 ( .A(\registers[576][1] ), .B(\registers[577][1] ), .C(
        \registers[578][1] ), .D(\registers[579][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5135) );
  MX4X1 U6760 ( .A(\registers[624][1] ), .B(\registers[625][1] ), .C(
        \registers[626][1] ), .D(\registers[627][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5120) );
  MX4X1 U6761 ( .A(\registers[608][1] ), .B(\registers[609][1] ), .C(
        \registers[610][1] ), .D(\registers[611][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5125) );
  MX4X1 U6762 ( .A(\registers[512][1] ), .B(\registers[513][1] ), .C(
        \registers[514][1] ), .D(\registers[515][1] ), .S0(n7479), .S1(n7719), 
        .Y(n5156) );
  MX4X1 U6763 ( .A(\registers[560][1] ), .B(\registers[561][1] ), .C(
        \registers[562][1] ), .D(\registers[563][1] ), .S0(n7478), .S1(n7719), 
        .Y(n5141) );
  MX4X1 U6764 ( .A(\registers[544][1] ), .B(\registers[545][1] ), .C(
        \registers[546][1] ), .D(\registers[547][1] ), .S0(n7478), .S1(n7719), 
        .Y(n5146) );
  MX4X1 U6765 ( .A(\registers[704][1] ), .B(\registers[705][1] ), .C(
        \registers[706][1] ), .D(\registers[707][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5093) );
  MX4X1 U6766 ( .A(\registers[752][1] ), .B(\registers[753][1] ), .C(
        \registers[754][1] ), .D(\registers[755][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5078) );
  MX4X1 U6767 ( .A(\registers[736][1] ), .B(\registers[737][1] ), .C(
        \registers[738][1] ), .D(\registers[739][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5083) );
  MX4X1 U6768 ( .A(\registers[640][1] ), .B(\registers[641][1] ), .C(
        \registers[642][1] ), .D(\registers[643][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5114) );
  MX4X1 U6769 ( .A(\registers[688][1] ), .B(\registers[689][1] ), .C(
        \registers[690][1] ), .D(\registers[691][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5099) );
  MX4X1 U6770 ( .A(\registers[672][1] ), .B(\registers[673][1] ), .C(
        \registers[674][1] ), .D(\registers[675][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5104) );
  MX4X1 U6771 ( .A(\registers[320][2] ), .B(\registers[321][2] ), .C(
        \registers[322][2] ), .D(\registers[323][2] ), .S0(n7504), .S1(n7743), 
        .Y(n5560) );
  MX4X1 U6772 ( .A(\registers[368][2] ), .B(\registers[369][2] ), .C(
        \registers[370][2] ), .D(\registers[371][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5545) );
  MX4X1 U6773 ( .A(\registers[352][2] ), .B(\registers[353][2] ), .C(
        \registers[354][2] ), .D(\registers[355][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5550) );
  MX4X1 U6774 ( .A(\registers[64][2] ), .B(\registers[65][2] ), .C(
        \registers[66][2] ), .D(\registers[67][2] ), .S0(n7509), .S1(n7748), 
        .Y(n5645) );
  MX4X1 U6775 ( .A(\registers[112][2] ), .B(\registers[113][2] ), .C(
        \registers[114][2] ), .D(\registers[115][2] ), .S0(n7508), .S1(n7747), 
        .Y(n5630) );
  MX4X1 U6776 ( .A(\registers[96][2] ), .B(\registers[97][2] ), .C(
        \registers[98][2] ), .D(\registers[99][2] ), .S0(n7509), .S1(n7747), 
        .Y(n5635) );
  MX4X1 U6777 ( .A(\registers[0][2] ), .B(\registers[1][2] ), .C(
        \registers[2][2] ), .D(\registers[3][2] ), .S0(n7511), .S1(n7749), .Y(
        n5666) );
  MX4X1 U6778 ( .A(\registers[48][2] ), .B(\registers[49][2] ), .C(
        \registers[50][2] ), .D(\registers[51][2] ), .S0(n7510), .S1(n7748), 
        .Y(n5651) );
  MX4X1 U6779 ( .A(\registers[32][2] ), .B(\registers[33][2] ), .C(
        \registers[34][2] ), .D(\registers[35][2] ), .S0(n7510), .S1(n7748), 
        .Y(n5656) );
  MX4X1 U6780 ( .A(\registers[192][2] ), .B(\registers[193][2] ), .C(
        \registers[194][2] ), .D(\registers[195][2] ), .S0(n7507), .S1(n7745), 
        .Y(n5603) );
  MX4X1 U6781 ( .A(\registers[240][2] ), .B(\registers[241][2] ), .C(
        \registers[242][2] ), .D(\registers[243][2] ), .S0(n7506), .S1(n7744), 
        .Y(n5588) );
  MX4X1 U6782 ( .A(\registers[224][2] ), .B(\registers[225][2] ), .C(
        \registers[226][2] ), .D(\registers[227][2] ), .S0(n7506), .S1(n7745), 
        .Y(n5593) );
  MX4X1 U6783 ( .A(\registers[128][2] ), .B(\registers[129][2] ), .C(
        \registers[130][2] ), .D(\registers[131][2] ), .S0(n7508), .S1(n7747), 
        .Y(n5624) );
  MX4X1 U6784 ( .A(\registers[176][2] ), .B(\registers[177][2] ), .C(
        \registers[178][2] ), .D(\registers[179][2] ), .S0(n7507), .S1(n7746), 
        .Y(n5609) );
  MX4X1 U6785 ( .A(\registers[160][2] ), .B(\registers[161][2] ), .C(
        \registers[162][2] ), .D(\registers[163][2] ), .S0(n7507), .S1(n7746), 
        .Y(n5614) );
  MX4X1 U6786 ( .A(\registers[832][2] ), .B(\registers[833][2] ), .C(
        \registers[834][2] ), .D(\registers[835][2] ), .S0(n7493), .S1(n7733), 
        .Y(n5390) );
  MX4X1 U6787 ( .A(\registers[880][2] ), .B(\registers[881][2] ), .C(
        \registers[882][2] ), .D(\registers[883][2] ), .S0(n7492), .S1(n7732), 
        .Y(n5375) );
  MX4X1 U6788 ( .A(\registers[864][2] ), .B(\registers[865][2] ), .C(
        \registers[866][2] ), .D(\registers[867][2] ), .S0(n7493), .S1(n7732), 
        .Y(n5380) );
  MX4X1 U6789 ( .A(\registers[768][2] ), .B(\registers[769][2] ), .C(
        \registers[770][2] ), .D(\registers[771][2] ), .S0(n7495), .S1(n7734), 
        .Y(n5411) );
  MX4X1 U6790 ( .A(\registers[816][2] ), .B(\registers[817][2] ), .C(
        \registers[818][2] ), .D(\registers[819][2] ), .S0(n7494), .S1(n7733), 
        .Y(n5396) );
  MX4X1 U6791 ( .A(\registers[800][2] ), .B(\registers[801][2] ), .C(
        \registers[802][2] ), .D(\registers[803][2] ), .S0(n7494), .S1(n7734), 
        .Y(n5401) );
  MX4X1 U6792 ( .A(\registers[960][2] ), .B(\registers[961][2] ), .C(
        \registers[962][2] ), .D(\registers[963][2] ), .S0(n7491), .S1(n7731), 
        .Y(n5348) );
  MX4X1 U6793 ( .A(\registers[1008][2] ), .B(\registers[1009][2] ), .C(
        \registers[1010][2] ), .D(\registers[1011][2] ), .S0(n7490), .S1(n7730), .Y(n5333) );
  MX4X1 U6794 ( .A(\registers[992][2] ), .B(\registers[993][2] ), .C(
        \registers[994][2] ), .D(\registers[995][2] ), .S0(n7490), .S1(n7730), 
        .Y(n5338) );
  MX4X1 U6795 ( .A(\registers[896][2] ), .B(\registers[897][2] ), .C(
        \registers[898][2] ), .D(\registers[899][2] ), .S0(n7492), .S1(n7732), 
        .Y(n5369) );
  MX4X1 U6796 ( .A(\registers[944][2] ), .B(\registers[945][2] ), .C(
        \registers[946][2] ), .D(\registers[947][2] ), .S0(n7491), .S1(n7731), 
        .Y(n5354) );
  MX4X1 U6797 ( .A(\registers[928][2] ), .B(\registers[929][2] ), .C(
        \registers[930][2] ), .D(\registers[931][2] ), .S0(n7491), .S1(n7731), 
        .Y(n5359) );
  MX4X1 U6798 ( .A(\registers[576][2] ), .B(\registers[577][2] ), .C(
        \registers[578][2] ), .D(\registers[579][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5475) );
  MX4X1 U6799 ( .A(\registers[624][2] ), .B(\registers[625][2] ), .C(
        \registers[626][2] ), .D(\registers[627][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5460) );
  MX4X1 U6800 ( .A(\registers[608][2] ), .B(\registers[609][2] ), .C(
        \registers[610][2] ), .D(\registers[611][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5465) );
  MX4X1 U6801 ( .A(\registers[512][2] ), .B(\registers[513][2] ), .C(
        \registers[514][2] ), .D(\registers[515][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5496) );
  MX4X1 U6802 ( .A(\registers[560][2] ), .B(\registers[561][2] ), .C(
        \registers[562][2] ), .D(\registers[563][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5481) );
  MX4X1 U6803 ( .A(\registers[544][2] ), .B(\registers[545][2] ), .C(
        \registers[546][2] ), .D(\registers[547][2] ), .S0(n7499), .S1(n7739), 
        .Y(n5486) );
  MX4X1 U6804 ( .A(\registers[704][2] ), .B(\registers[705][2] ), .C(
        \registers[706][2] ), .D(\registers[707][2] ), .S0(n7496), .S1(n7735), 
        .Y(n5433) );
  MX4X1 U6805 ( .A(\registers[752][2] ), .B(\registers[753][2] ), .C(
        \registers[754][2] ), .D(\registers[755][2] ), .S0(n7495), .S1(n7735), 
        .Y(n5418) );
  MX4X1 U6806 ( .A(\registers[736][2] ), .B(\registers[737][2] ), .C(
        \registers[738][2] ), .D(\registers[739][2] ), .S0(n7495), .S1(n7735), 
        .Y(n5423) );
  MX4X1 U6807 ( .A(\registers[640][2] ), .B(\registers[641][2] ), .C(
        \registers[642][2] ), .D(\registers[643][2] ), .S0(n7497), .S1(n7737), 
        .Y(n5454) );
  MX4X1 U6808 ( .A(\registers[688][2] ), .B(\registers[689][2] ), .C(
        \registers[690][2] ), .D(\registers[691][2] ), .S0(n7496), .S1(n7736), 
        .Y(n5439) );
  MX4X1 U6809 ( .A(\registers[672][2] ), .B(\registers[673][2] ), .C(
        \registers[674][2] ), .D(\registers[675][2] ), .S0(n7497), .S1(n7736), 
        .Y(n5444) );
  MX4X1 U6810 ( .A(\registers[320][3] ), .B(\registers[321][3] ), .C(
        \registers[322][3] ), .D(\registers[323][3] ), .S0(n7525), .S1(n7763), 
        .Y(n5900) );
  MX4X1 U6811 ( .A(\registers[368][3] ), .B(\registers[369][3] ), .C(
        \registers[370][3] ), .D(\registers[371][3] ), .S0(n7524), .S1(n7762), 
        .Y(n5885) );
  MX4X1 U6812 ( .A(\registers[352][3] ), .B(\registers[353][3] ), .C(
        \registers[354][3] ), .D(\registers[355][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5890) );
  MX4X1 U6813 ( .A(\registers[64][3] ), .B(\registers[65][3] ), .C(
        \registers[66][3] ), .D(\registers[67][3] ), .S0(n7531), .S1(n7767), 
        .Y(n5985) );
  MX4X1 U6814 ( .A(\registers[112][3] ), .B(\registers[113][3] ), .C(
        \registers[114][3] ), .D(\registers[115][3] ), .S0(n7530), .S1(n7767), 
        .Y(n5970) );
  MX4X1 U6815 ( .A(\registers[96][3] ), .B(\registers[97][3] ), .C(
        \registers[98][3] ), .D(\registers[99][3] ), .S0(n7530), .S1(n7767), 
        .Y(n5975) );
  MX4X1 U6816 ( .A(\registers[0][3] ), .B(\registers[1][3] ), .C(
        \registers[2][3] ), .D(\registers[3][3] ), .S0(n7532), .S1(n7769), .Y(
        n6006) );
  MX4X1 U6817 ( .A(\registers[48][3] ), .B(\registers[49][3] ), .C(
        \registers[50][3] ), .D(\registers[51][3] ), .S0(n7531), .S1(n7768), 
        .Y(n5991) );
  MX4X1 U6818 ( .A(\registers[32][3] ), .B(\registers[33][3] ), .C(
        \registers[34][3] ), .D(\registers[35][3] ), .S0(n7531), .S1(n7768), 
        .Y(n5996) );
  MX4X1 U6819 ( .A(\registers[192][3] ), .B(\registers[193][3] ), .C(
        \registers[194][3] ), .D(\registers[195][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5943) );
  MX4X1 U6820 ( .A(\registers[240][3] ), .B(\registers[241][3] ), .C(
        \registers[242][3] ), .D(\registers[243][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5928) );
  MX4X1 U6821 ( .A(\registers[224][3] ), .B(\registers[225][3] ), .C(
        \registers[226][3] ), .D(\registers[227][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5933) );
  MX4X1 U6822 ( .A(\registers[128][3] ), .B(\registers[129][3] ), .C(
        \registers[130][3] ), .D(\registers[131][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5964) );
  MX4X1 U6823 ( .A(\registers[176][3] ), .B(\registers[177][3] ), .C(
        \registers[178][3] ), .D(\registers[179][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5949) );
  MX4X1 U6824 ( .A(\registers[160][3] ), .B(\registers[161][3] ), .C(
        \registers[162][3] ), .D(\registers[163][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5954) );
  MX4X1 U6825 ( .A(\registers[832][3] ), .B(\registers[833][3] ), .C(
        \registers[834][3] ), .D(\registers[835][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5730) );
  MX4X1 U6826 ( .A(\registers[880][3] ), .B(\registers[881][3] ), .C(
        \registers[882][3] ), .D(\registers[883][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5715) );
  MX4X1 U6827 ( .A(\registers[864][3] ), .B(\registers[865][3] ), .C(
        \registers[866][3] ), .D(\registers[867][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5720) );
  MX4X1 U6828 ( .A(\registers[768][3] ), .B(\registers[769][3] ), .C(
        \registers[770][3] ), .D(\registers[771][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5751) );
  MX4X1 U6829 ( .A(\registers[816][3] ), .B(\registers[817][3] ), .C(
        \registers[818][3] ), .D(\registers[819][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5736) );
  MX4X1 U6830 ( .A(\registers[800][3] ), .B(\registers[801][3] ), .C(
        \registers[802][3] ), .D(\registers[803][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5741) );
  MX4X1 U6831 ( .A(\registers[960][3] ), .B(\registers[961][3] ), .C(
        \registers[962][3] ), .D(\registers[963][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5688) );
  MX4X1 U6832 ( .A(\registers[1008][3] ), .B(\registers[1009][3] ), .C(
        \registers[1010][3] ), .D(\registers[1011][3] ), .S0(n7511), .S1(n7749), .Y(n5673) );
  MX4X1 U6833 ( .A(\registers[992][3] ), .B(\registers[993][3] ), .C(
        \registers[994][3] ), .D(\registers[995][3] ), .S0(n7511), .S1(n7750), 
        .Y(n5678) );
  MX4X1 U6834 ( .A(\registers[896][3] ), .B(\registers[897][3] ), .C(
        \registers[898][3] ), .D(\registers[899][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5709) );
  MX4X1 U6835 ( .A(\registers[944][3] ), .B(\registers[945][3] ), .C(
        \registers[946][3] ), .D(\registers[947][3] ), .S0(n7512), .S1(n7751), 
        .Y(n5694) );
  MX4X1 U6836 ( .A(\registers[928][3] ), .B(\registers[929][3] ), .C(
        \registers[930][3] ), .D(\registers[931][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5699) );
  MX4X1 U6837 ( .A(\registers[576][3] ), .B(\registers[577][3] ), .C(
        \registers[578][3] ), .D(\registers[579][3] ), .S0(n7520), .S1(n7758), 
        .Y(n5815) );
  MX4X1 U6838 ( .A(\registers[624][3] ), .B(\registers[625][3] ), .C(
        \registers[626][3] ), .D(\registers[627][3] ), .S0(n7519), .S1(n7757), 
        .Y(n5800) );
  MX4X1 U6839 ( .A(\registers[608][3] ), .B(\registers[609][3] ), .C(
        \registers[610][3] ), .D(\registers[611][3] ), .S0(n7519), .S1(n7757), 
        .Y(n5805) );
  MX4X1 U6840 ( .A(\registers[512][3] ), .B(\registers[513][3] ), .C(
        \registers[514][3] ), .D(\registers[515][3] ), .S0(n7521), .S1(n7759), 
        .Y(n5836) );
  MX4X1 U6841 ( .A(\registers[560][3] ), .B(\registers[561][3] ), .C(
        \registers[562][3] ), .D(\registers[563][3] ), .S0(n7520), .S1(n7758), 
        .Y(n5821) );
  MX4X1 U6842 ( .A(\registers[544][3] ), .B(\registers[545][3] ), .C(
        \registers[546][3] ), .D(\registers[547][3] ), .S0(n7521), .S1(n7758), 
        .Y(n5826) );
  MX4X1 U6843 ( .A(\registers[704][3] ), .B(\registers[705][3] ), .C(
        \registers[706][3] ), .D(\registers[707][3] ), .S0(n7517), .S1(n7755), 
        .Y(n5773) );
  MX4X1 U6844 ( .A(\registers[752][3] ), .B(\registers[753][3] ), .C(
        \registers[754][3] ), .D(\registers[755][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5758) );
  MX4X1 U6845 ( .A(\registers[736][3] ), .B(\registers[737][3] ), .C(
        \registers[738][3] ), .D(\registers[739][3] ), .S0(n7517), .S1(n7755), 
        .Y(n5763) );
  MX4X1 U6846 ( .A(\registers[640][3] ), .B(\registers[641][3] ), .C(
        \registers[642][3] ), .D(\registers[643][3] ), .S0(n7519), .S1(n7756), 
        .Y(n5794) );
  MX4X1 U6847 ( .A(\registers[688][3] ), .B(\registers[689][3] ), .C(
        \registers[690][3] ), .D(\registers[691][3] ), .S0(n7518), .S1(n7755), 
        .Y(n5779) );
  MX4X1 U6848 ( .A(\registers[672][3] ), .B(\registers[673][3] ), .C(
        \registers[674][3] ), .D(\registers[675][3] ), .S0(n7518), .S1(n7756), 
        .Y(n5784) );
  MX4X1 U6849 ( .A(\registers[320][4] ), .B(\registers[321][4] ), .C(
        \registers[322][4] ), .D(\registers[323][4] ), .S0(n7547), .S1(n7782), 
        .Y(n6240) );
  MX4X1 U6850 ( .A(\registers[368][4] ), .B(\registers[369][4] ), .C(
        \registers[370][4] ), .D(\registers[371][4] ), .S0(n7546), .S1(n7781), 
        .Y(n6225) );
  MX4X1 U6851 ( .A(\registers[352][4] ), .B(\registers[353][4] ), .C(
        \registers[354][4] ), .D(\registers[355][4] ), .S0(n7546), .S1(n7782), 
        .Y(n6230) );
  MX4X1 U6852 ( .A(\registers[64][4] ), .B(\registers[65][4] ), .C(
        \registers[66][4] ), .D(\registers[67][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6325) );
  MX4X1 U6853 ( .A(\registers[112][4] ), .B(\registers[113][4] ), .C(
        \registers[114][4] ), .D(\registers[115][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6310) );
  MX4X1 U6854 ( .A(\registers[96][4] ), .B(\registers[97][4] ), .C(
        \registers[98][4] ), .D(\registers[99][4] ), .S0(n7551), .S1(n7787), 
        .Y(n6315) );
  MX4X1 U6855 ( .A(\registers[0][4] ), .B(\registers[1][4] ), .C(
        \registers[2][4] ), .D(\registers[3][4] ), .S0(n7553), .S1(n7788), .Y(
        n6346) );
  MX4X1 U6856 ( .A(\registers[48][4] ), .B(\registers[49][4] ), .C(
        \registers[50][4] ), .D(\registers[51][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6331) );
  MX4X1 U6857 ( .A(\registers[32][4] ), .B(\registers[33][4] ), .C(
        \registers[34][4] ), .D(\registers[35][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6336) );
  MX4X1 U6858 ( .A(\registers[192][4] ), .B(\registers[193][4] ), .C(
        \registers[194][4] ), .D(\registers[195][4] ), .S0(n7549), .S1(n7785), 
        .Y(n6283) );
  MX4X1 U6859 ( .A(\registers[240][4] ), .B(\registers[241][4] ), .C(
        \registers[242][4] ), .D(\registers[243][4] ), .S0(n7548), .S1(n7784), 
        .Y(n6268) );
  MX4X1 U6860 ( .A(\registers[224][4] ), .B(\registers[225][4] ), .C(
        \registers[226][4] ), .D(\registers[227][4] ), .S0(n7549), .S1(n7784), 
        .Y(n6273) );
  MX4X1 U6861 ( .A(\registers[128][4] ), .B(\registers[129][4] ), .C(
        \registers[130][4] ), .D(\registers[131][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6304) );
  MX4X1 U6862 ( .A(\registers[176][4] ), .B(\registers[177][4] ), .C(
        \registers[178][4] ), .D(\registers[179][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6289) );
  MX4X1 U6863 ( .A(\registers[160][4] ), .B(\registers[161][4] ), .C(
        \registers[162][4] ), .D(\registers[163][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6294) );
  MX4X1 U6864 ( .A(\registers[832][4] ), .B(\registers[833][4] ), .C(
        \registers[834][4] ), .D(\registers[835][4] ), .S0(n7536), .S1(n7772), 
        .Y(n6070) );
  MX4X1 U6865 ( .A(\registers[880][4] ), .B(\registers[881][4] ), .C(
        \registers[882][4] ), .D(\registers[883][4] ), .S0(n7535), .S1(n7771), 
        .Y(n6055) );
  MX4X1 U6866 ( .A(\registers[864][4] ), .B(\registers[865][4] ), .C(
        \registers[866][4] ), .D(\registers[867][4] ), .S0(n7535), .S1(n7772), 
        .Y(n6060) );
  MX4X1 U6867 ( .A(\registers[768][4] ), .B(\registers[769][4] ), .C(
        \registers[770][4] ), .D(\registers[771][4] ), .S0(n7537), .S1(n7774), 
        .Y(n6091) );
  MX4X1 U6868 ( .A(\registers[816][4] ), .B(\registers[817][4] ), .C(
        \registers[818][4] ), .D(\registers[819][4] ), .S0(n7536), .S1(n7773), 
        .Y(n6076) );
  MX4X1 U6869 ( .A(\registers[800][4] ), .B(\registers[801][4] ), .C(
        \registers[802][4] ), .D(\registers[803][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6081) );
  MX4X1 U6870 ( .A(\registers[960][4] ), .B(\registers[961][4] ), .C(
        \registers[962][4] ), .D(\registers[963][4] ), .S0(n7533), .S1(n7770), 
        .Y(n6028) );
  MX4X1 U6871 ( .A(\registers[1008][4] ), .B(\registers[1009][4] ), .C(
        \registers[1010][4] ), .D(\registers[1011][4] ), .S0(n7532), .S1(n7769), .Y(n6013) );
  MX4X1 U6872 ( .A(\registers[992][4] ), .B(\registers[993][4] ), .C(
        \registers[994][4] ), .D(\registers[995][4] ), .S0(n7533), .S1(n7769), 
        .Y(n6018) );
  MX4X1 U6873 ( .A(\registers[896][4] ), .B(\registers[897][4] ), .C(
        \registers[898][4] ), .D(\registers[899][4] ), .S0(n7535), .S1(n7771), 
        .Y(n6049) );
  MX4X1 U6874 ( .A(\registers[944][4] ), .B(\registers[945][4] ), .C(
        \registers[946][4] ), .D(\registers[947][4] ), .S0(n7534), .S1(n7770), 
        .Y(n6034) );
  MX4X1 U6875 ( .A(\registers[928][4] ), .B(\registers[929][4] ), .C(
        \registers[930][4] ), .D(\registers[931][4] ), .S0(n7534), .S1(n7771), 
        .Y(n6039) );
  MX4X1 U6876 ( .A(\registers[576][4] ), .B(\registers[577][4] ), .C(
        \registers[578][4] ), .D(\registers[579][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6155) );
  MX4X1 U6877 ( .A(\registers[624][4] ), .B(\registers[625][4] ), .C(
        \registers[626][4] ), .D(\registers[627][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6140) );
  MX4X1 U6878 ( .A(\registers[608][4] ), .B(\registers[609][4] ), .C(
        \registers[610][4] ), .D(\registers[611][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6145) );
  MX4X1 U6879 ( .A(\registers[512][4] ), .B(\registers[513][4] ), .C(
        \registers[514][4] ), .D(\registers[515][4] ), .S0(n7543), .S1(n7779), 
        .Y(n6176) );
  MX4X1 U6880 ( .A(\registers[560][4] ), .B(\registers[561][4] ), .C(
        \registers[562][4] ), .D(\registers[563][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6161) );
  MX4X1 U6881 ( .A(\registers[544][4] ), .B(\registers[545][4] ), .C(
        \registers[546][4] ), .D(\registers[547][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6166) );
  MX4X1 U6882 ( .A(\registers[704][4] ), .B(\registers[705][4] ), .C(
        \registers[706][4] ), .D(\registers[707][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6113) );
  MX4X1 U6883 ( .A(\registers[752][4] ), .B(\registers[753][4] ), .C(
        \registers[754][4] ), .D(\registers[755][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6098) );
  MX4X1 U6884 ( .A(\registers[736][4] ), .B(\registers[737][4] ), .C(
        \registers[738][4] ), .D(\registers[739][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6103) );
  MX4X1 U6885 ( .A(\registers[640][4] ), .B(\registers[641][4] ), .C(
        \registers[642][4] ), .D(\registers[643][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6134) );
  MX4X1 U6886 ( .A(\registers[688][4] ), .B(\registers[689][4] ), .C(
        \registers[690][4] ), .D(\registers[691][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6119) );
  MX4X1 U6887 ( .A(\registers[672][4] ), .B(\registers[673][4] ), .C(
        \registers[674][4] ), .D(\registers[675][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6124) );
  MX4X1 U6888 ( .A(\registers[320][5] ), .B(\registers[321][5] ), .C(
        \registers[322][5] ), .D(\registers[323][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6580) );
  MX4X1 U6889 ( .A(\registers[368][5] ), .B(\registers[369][5] ), .C(
        \registers[370][5] ), .D(\registers[371][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6565) );
  MX4X1 U6890 ( .A(\registers[352][5] ), .B(\registers[353][5] ), .C(
        \registers[354][5] ), .D(\registers[355][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6570) );
  MX4X1 U6891 ( .A(\registers[64][5] ), .B(\registers[65][5] ), .C(
        \registers[66][5] ), .D(\registers[67][5] ), .S0(n7573), .S1(n7806), 
        .Y(n6665) );
  MX4X1 U6892 ( .A(\registers[112][5] ), .B(\registers[113][5] ), .C(
        \registers[114][5] ), .D(\registers[115][5] ), .S0(n7572), .S1(n7805), 
        .Y(n6650) );
  MX4X1 U6893 ( .A(\registers[96][5] ), .B(\registers[97][5] ), .C(
        \registers[98][5] ), .D(\registers[99][5] ), .S0(n7573), .S1(n7805), 
        .Y(n6655) );
  MX4X1 U6894 ( .A(\registers[0][5] ), .B(\registers[1][5] ), .C(
        \registers[2][5] ), .D(\registers[3][5] ), .S0(n7575), .S1(n7807), .Y(
        n6686) );
  MX4X1 U6895 ( .A(\registers[48][5] ), .B(\registers[49][5] ), .C(
        \registers[50][5] ), .D(\registers[51][5] ), .S0(n7574), .S1(n7806), 
        .Y(n6671) );
  MX4X1 U6896 ( .A(\registers[32][5] ), .B(\registers[33][5] ), .C(
        \registers[34][5] ), .D(\registers[35][5] ), .S0(n7574), .S1(n7806), 
        .Y(n6676) );
  MX4X1 U6897 ( .A(\registers[192][5] ), .B(\registers[193][5] ), .C(
        \registers[194][5] ), .D(\registers[195][5] ), .S0(n7571), .S1(n7693), 
        .Y(n6623) );
  MX4X1 U6898 ( .A(\registers[240][5] ), .B(\registers[241][5] ), .C(
        \registers[242][5] ), .D(\registers[243][5] ), .S0(n7570), .S1(n7803), 
        .Y(n6608) );
  MX4X1 U6899 ( .A(\registers[224][5] ), .B(\registers[225][5] ), .C(
        \registers[226][5] ), .D(\registers[227][5] ), .S0(n7570), .S1(n7799), 
        .Y(n6613) );
  MX4X1 U6900 ( .A(\registers[128][5] ), .B(\registers[129][5] ), .C(
        \registers[130][5] ), .D(\registers[131][5] ), .S0(n7572), .S1(n7805), 
        .Y(n6644) );
  MX4X1 U6901 ( .A(\registers[176][5] ), .B(\registers[177][5] ), .C(
        \registers[178][5] ), .D(\registers[179][5] ), .S0(n7571), .S1(n7804), 
        .Y(n6629) );
  MX4X1 U6902 ( .A(\registers[160][5] ), .B(\registers[161][5] ), .C(
        \registers[162][5] ), .D(\registers[163][5] ), .S0(n7571), .S1(n7804), 
        .Y(n6634) );
  MX4X1 U6903 ( .A(\registers[832][5] ), .B(\registers[833][5] ), .C(
        \registers[834][5] ), .D(\registers[835][5] ), .S0(n7557), .S1(n7792), 
        .Y(n6410) );
  MX4X1 U6904 ( .A(\registers[880][5] ), .B(\registers[881][5] ), .C(
        \registers[882][5] ), .D(\registers[883][5] ), .S0(n7556), .S1(n7791), 
        .Y(n6395) );
  MX4X1 U6905 ( .A(\registers[864][5] ), .B(\registers[865][5] ), .C(
        \registers[866][5] ), .D(\registers[867][5] ), .S0(n7557), .S1(n7791), 
        .Y(n6400) );
  MX4X1 U6906 ( .A(\registers[768][5] ), .B(\registers[769][5] ), .C(
        \registers[770][5] ), .D(\registers[771][5] ), .S0(n7559), .S1(n7793), 
        .Y(n6431) );
  MX4X1 U6907 ( .A(\registers[816][5] ), .B(\registers[817][5] ), .C(
        \registers[818][5] ), .D(\registers[819][5] ), .S0(n7558), .S1(n7792), 
        .Y(n6416) );
  MX4X1 U6908 ( .A(\registers[800][5] ), .B(\registers[801][5] ), .C(
        \registers[802][5] ), .D(\registers[803][5] ), .S0(n7558), .S1(n7793), 
        .Y(n6421) );
  MX4X1 U6909 ( .A(\registers[960][5] ), .B(\registers[961][5] ), .C(
        \registers[962][5] ), .D(\registers[963][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6368) );
  MX4X1 U6910 ( .A(\registers[1008][5] ), .B(\registers[1009][5] ), .C(
        \registers[1010][5] ), .D(\registers[1011][5] ), .S0(n7554), .S1(n7789), .Y(n6353) );
  MX4X1 U6911 ( .A(\registers[992][5] ), .B(\registers[993][5] ), .C(
        \registers[994][5] ), .D(\registers[995][5] ), .S0(n7554), .S1(n7789), 
        .Y(n6358) );
  MX4X1 U6912 ( .A(\registers[896][5] ), .B(\registers[897][5] ), .C(
        \registers[898][5] ), .D(\registers[899][5] ), .S0(n7556), .S1(n7791), 
        .Y(n6389) );
  MX4X1 U6913 ( .A(\registers[944][5] ), .B(\registers[945][5] ), .C(
        \registers[946][5] ), .D(\registers[947][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6374) );
  MX4X1 U6914 ( .A(\registers[928][5] ), .B(\registers[929][5] ), .C(
        \registers[930][5] ), .D(\registers[931][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6379) );
  MX4X1 U6915 ( .A(\registers[576][5] ), .B(\registers[577][5] ), .C(
        \registers[578][5] ), .D(\registers[579][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6495) );
  MX4X1 U6916 ( .A(\registers[624][5] ), .B(\registers[625][5] ), .C(
        \registers[626][5] ), .D(\registers[627][5] ), .S0(n7562), .S1(n7796), 
        .Y(n6480) );
  MX4X1 U6917 ( .A(\registers[608][5] ), .B(\registers[609][5] ), .C(
        \registers[610][5] ), .D(\registers[611][5] ), .S0(n7562), .S1(n7796), 
        .Y(n6485) );
  MX4X1 U6918 ( .A(\registers[512][5] ), .B(\registers[513][5] ), .C(
        \registers[514][5] ), .D(\registers[515][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6516) );
  MX4X1 U6919 ( .A(\registers[560][5] ), .B(\registers[561][5] ), .C(
        \registers[562][5] ), .D(\registers[563][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6501) );
  MX4X1 U6920 ( .A(\registers[544][5] ), .B(\registers[545][5] ), .C(
        \registers[546][5] ), .D(\registers[547][5] ), .S0(n7563), .S1(n7798), 
        .Y(n6506) );
  MX4X1 U6921 ( .A(\registers[704][5] ), .B(\registers[705][5] ), .C(
        \registers[706][5] ), .D(\registers[707][5] ), .S0(n7560), .S1(n7795), 
        .Y(n6453) );
  MX4X1 U6922 ( .A(\registers[752][5] ), .B(\registers[753][5] ), .C(
        \registers[754][5] ), .D(\registers[755][5] ), .S0(n7559), .S1(n7794), 
        .Y(n6438) );
  MX4X1 U6923 ( .A(\registers[736][5] ), .B(\registers[737][5] ), .C(
        \registers[738][5] ), .D(\registers[739][5] ), .S0(n7559), .S1(n7794), 
        .Y(n6443) );
  MX4X1 U6924 ( .A(\registers[640][5] ), .B(\registers[641][5] ), .C(
        \registers[642][5] ), .D(\registers[643][5] ), .S0(n7561), .S1(n7796), 
        .Y(n6474) );
  MX4X1 U6925 ( .A(\registers[688][5] ), .B(\registers[689][5] ), .C(
        \registers[690][5] ), .D(\registers[691][5] ), .S0(n7560), .S1(n7795), 
        .Y(n6459) );
  MX4X1 U6926 ( .A(\registers[672][5] ), .B(\registers[673][5] ), .C(
        \registers[674][5] ), .D(\registers[675][5] ), .S0(n7561), .S1(n7795), 
        .Y(n6464) );
  MX4X1 U6927 ( .A(\registers[320][6] ), .B(\registers[321][6] ), .C(
        \registers[322][6] ), .D(\registers[323][6] ), .S0(n7589), .S1(n7821), 
        .Y(n6920) );
  MX4X1 U6928 ( .A(\registers[368][6] ), .B(\registers[369][6] ), .C(
        \registers[370][6] ), .D(\registers[371][6] ), .S0(n7588), .S1(n7820), 
        .Y(n6905) );
  MX4X1 U6929 ( .A(\registers[352][6] ), .B(\registers[353][6] ), .C(
        \registers[354][6] ), .D(\registers[355][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6910) );
  MX4X1 U6930 ( .A(\registers[64][6] ), .B(\registers[65][6] ), .C(
        \registers[66][6] ), .D(\registers[67][6] ), .S0(n7595), .S1(n7826), 
        .Y(n7005) );
  MX4X1 U6931 ( .A(\registers[112][6] ), .B(\registers[113][6] ), .C(
        \registers[114][6] ), .D(\registers[115][6] ), .S0(n7594), .S1(n7825), 
        .Y(n6990) );
  MX4X1 U6932 ( .A(\registers[96][6] ), .B(\registers[97][6] ), .C(
        \registers[98][6] ), .D(\registers[99][6] ), .S0(n7594), .S1(n7825), 
        .Y(n6995) );
  MX4X1 U6933 ( .A(\registers[0][6] ), .B(\registers[1][6] ), .C(
        \registers[2][6] ), .D(\registers[3][6] ), .S0(n7596), .S1(n7827), .Y(
        n7026) );
  MX4X1 U6934 ( .A(\registers[48][6] ), .B(\registers[49][6] ), .C(
        \registers[50][6] ), .D(\registers[51][6] ), .S0(n7595), .S1(n7826), 
        .Y(n7011) );
  MX4X1 U6935 ( .A(\registers[32][6] ), .B(\registers[33][6] ), .C(
        \registers[34][6] ), .D(\registers[35][6] ), .S0(n7595), .S1(n7826), 
        .Y(n7016) );
  MX4X1 U6936 ( .A(\registers[192][6] ), .B(\registers[193][6] ), .C(
        \registers[194][6] ), .D(\registers[195][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6963) );
  MX4X1 U6937 ( .A(\registers[240][6] ), .B(\registers[241][6] ), .C(
        \registers[242][6] ), .D(\registers[243][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6948) );
  MX4X1 U6938 ( .A(\registers[224][6] ), .B(\registers[225][6] ), .C(
        \registers[226][6] ), .D(\registers[227][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6953) );
  MX4X1 U6939 ( .A(\registers[128][6] ), .B(\registers[129][6] ), .C(
        \registers[130][6] ), .D(\registers[131][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6984) );
  MX4X1 U6940 ( .A(\registers[176][6] ), .B(\registers[177][6] ), .C(
        \registers[178][6] ), .D(\registers[179][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6969) );
  MX4X1 U6941 ( .A(\registers[160][6] ), .B(\registers[161][6] ), .C(
        \registers[162][6] ), .D(\registers[163][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6974) );
  MX4X1 U6942 ( .A(\registers[832][6] ), .B(\registers[833][6] ), .C(
        \registers[834][6] ), .D(\registers[835][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6750) );
  MX4X1 U6943 ( .A(\registers[880][6] ), .B(\registers[881][6] ), .C(
        \registers[882][6] ), .D(\registers[883][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6735) );
  MX4X1 U6944 ( .A(\registers[864][6] ), .B(\registers[865][6] ), .C(
        \registers[866][6] ), .D(\registers[867][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6740) );
  MX4X1 U6945 ( .A(\registers[768][6] ), .B(\registers[769][6] ), .C(
        \registers[770][6] ), .D(\registers[771][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6771) );
  MX4X1 U6946 ( .A(\registers[816][6] ), .B(\registers[817][6] ), .C(
        \registers[818][6] ), .D(\registers[819][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6756) );
  MX4X1 U6947 ( .A(\registers[800][6] ), .B(\registers[801][6] ), .C(
        \registers[802][6] ), .D(\registers[803][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6761) );
  MX4X1 U6948 ( .A(\registers[960][6] ), .B(\registers[961][6] ), .C(
        \registers[962][6] ), .D(\registers[963][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6708) );
  MX4X1 U6949 ( .A(\registers[1008][6] ), .B(\registers[1009][6] ), .C(
        \registers[1010][6] ), .D(\registers[1011][6] ), .S0(n7575), .S1(n7807), .Y(n6693) );
  MX4X1 U6950 ( .A(\registers[992][6] ), .B(\registers[993][6] ), .C(
        \registers[994][6] ), .D(\registers[995][6] ), .S0(n7575), .S1(n7808), 
        .Y(n6698) );
  MX4X1 U6951 ( .A(\registers[896][6] ), .B(\registers[897][6] ), .C(
        \registers[898][6] ), .D(\registers[899][6] ), .S0(n7577), .S1(n7810), 
        .Y(n6729) );
  MX4X1 U6952 ( .A(\registers[944][6] ), .B(\registers[945][6] ), .C(
        \registers[946][6] ), .D(\registers[947][6] ), .S0(n7576), .S1(n7809), 
        .Y(n6714) );
  MX4X1 U6953 ( .A(\registers[928][6] ), .B(\registers[929][6] ), .C(
        \registers[930][6] ), .D(\registers[931][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6719) );
  MX4X1 U6954 ( .A(\registers[576][6] ), .B(\registers[577][6] ), .C(
        \registers[578][6] ), .D(\registers[579][6] ), .S0(n7584), .S1(n7816), 
        .Y(n6835) );
  MX4X1 U6955 ( .A(\registers[624][6] ), .B(\registers[625][6] ), .C(
        \registers[626][6] ), .D(\registers[627][6] ), .S0(n7583), .S1(n7815), 
        .Y(n6820) );
  MX4X1 U6956 ( .A(\registers[608][6] ), .B(\registers[609][6] ), .C(
        \registers[610][6] ), .D(\registers[611][6] ), .S0(n7583), .S1(n7815), 
        .Y(n6825) );
  MX4X1 U6957 ( .A(\registers[512][6] ), .B(\registers[513][6] ), .C(
        \registers[514][6] ), .D(\registers[515][6] ), .S0(n7585), .S1(n7817), 
        .Y(n6856) );
  MX4X1 U6958 ( .A(\registers[560][6] ), .B(\registers[561][6] ), .C(
        \registers[562][6] ), .D(\registers[563][6] ), .S0(n7584), .S1(n7816), 
        .Y(n6841) );
  MX4X1 U6959 ( .A(\registers[544][6] ), .B(\registers[545][6] ), .C(
        \registers[546][6] ), .D(\registers[547][6] ), .S0(n7585), .S1(n7816), 
        .Y(n6846) );
  MX4X1 U6960 ( .A(\registers[704][6] ), .B(\registers[705][6] ), .C(
        \registers[706][6] ), .D(\registers[707][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6793) );
  MX4X1 U6961 ( .A(\registers[752][6] ), .B(\registers[753][6] ), .C(
        \registers[754][6] ), .D(\registers[755][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6778) );
  MX4X1 U6962 ( .A(\registers[736][6] ), .B(\registers[737][6] ), .C(
        \registers[738][6] ), .D(\registers[739][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6783) );
  MX4X1 U6963 ( .A(\registers[640][6] ), .B(\registers[641][6] ), .C(
        \registers[642][6] ), .D(\registers[643][6] ), .S0(n7583), .S1(n7814), 
        .Y(n6814) );
  MX4X1 U6964 ( .A(\registers[688][6] ), .B(\registers[689][6] ), .C(
        \registers[690][6] ), .D(\registers[691][6] ), .S0(n7582), .S1(n7814), 
        .Y(n6799) );
  MX4X1 U6965 ( .A(\registers[672][6] ), .B(\registers[673][6] ), .C(
        \registers[674][6] ), .D(\registers[675][6] ), .S0(n7582), .S1(n7814), 
        .Y(n6804) );
  MX4X1 U6966 ( .A(\registers[320][7] ), .B(\registers[321][7] ), .C(
        \registers[322][7] ), .D(\registers[323][7] ), .S0(n7611), .S1(n7840), 
        .Y(n7260) );
  MX4X1 U6967 ( .A(\registers[368][7] ), .B(\registers[369][7] ), .C(
        \registers[370][7] ), .D(\registers[371][7] ), .S0(n7610), .S1(n7839), 
        .Y(n7245) );
  MX4X1 U6968 ( .A(\registers[352][7] ), .B(\registers[353][7] ), .C(
        \registers[354][7] ), .D(\registers[355][7] ), .S0(n7610), .S1(n7840), 
        .Y(n7250) );
  MX4X1 U6969 ( .A(\registers[192][7] ), .B(\registers[193][7] ), .C(
        \registers[194][7] ), .D(\registers[195][7] ), .S0(n7613), .S1(n7843), 
        .Y(n7303) );
  MX4X1 U6970 ( .A(\registers[240][7] ), .B(\registers[241][7] ), .C(
        \registers[242][7] ), .D(\registers[243][7] ), .S0(n7612), .S1(n7842), 
        .Y(n7288) );
  MX4X1 U6971 ( .A(\registers[224][7] ), .B(\registers[225][7] ), .C(
        \registers[226][7] ), .D(\registers[227][7] ), .S0(n7613), .S1(n7842), 
        .Y(n7293) );
  MX4X1 U6972 ( .A(\registers[64][7] ), .B(\registers[65][7] ), .C(
        \registers[66][7] ), .D(\registers[67][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7345) );
  MX4X1 U6973 ( .A(\registers[112][7] ), .B(\registers[113][7] ), .C(
        \registers[114][7] ), .D(\registers[115][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7330) );
  MX4X1 U6974 ( .A(\registers[96][7] ), .B(\registers[97][7] ), .C(
        \registers[98][7] ), .D(\registers[99][7] ), .S0(n7615), .S1(n7845), 
        .Y(n7335) );
  MX4X1 U6975 ( .A(\registers[0][7] ), .B(\registers[1][7] ), .C(
        \registers[2][7] ), .D(\registers[3][7] ), .S0(n7617), .S1(n7846), .Y(
        n7366) );
  MX4X1 U6976 ( .A(\registers[48][7] ), .B(\registers[49][7] ), .C(
        \registers[50][7] ), .D(\registers[51][7] ), .S0(n7616), .S1(n7846), 
        .Y(n7351) );
  MX4X1 U6977 ( .A(\registers[32][7] ), .B(\registers[33][7] ), .C(
        \registers[34][7] ), .D(\registers[35][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7356) );
  MX4X1 U6978 ( .A(\registers[128][7] ), .B(\registers[129][7] ), .C(
        \registers[130][7] ), .D(\registers[131][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7324) );
  MX4X1 U6979 ( .A(\registers[176][7] ), .B(\registers[177][7] ), .C(
        \registers[178][7] ), .D(\registers[179][7] ), .S0(n7614), .S1(n7843), 
        .Y(n7309) );
  MX4X1 U6980 ( .A(\registers[160][7] ), .B(\registers[161][7] ), .C(
        \registers[162][7] ), .D(\registers[163][7] ), .S0(n7614), .S1(n7843), 
        .Y(n7314) );
  MX4X1 U6981 ( .A(\registers[832][7] ), .B(\registers[833][7] ), .C(
        \registers[834][7] ), .D(\registers[835][7] ), .S0(n7600), .S1(n7830), 
        .Y(n7090) );
  MX4X1 U6982 ( .A(\registers[880][7] ), .B(\registers[881][7] ), .C(
        \registers[882][7] ), .D(\registers[883][7] ), .S0(n7599), .S1(n7830), 
        .Y(n7075) );
  MX4X1 U6983 ( .A(\registers[864][7] ), .B(\registers[865][7] ), .C(
        \registers[866][7] ), .D(\registers[867][7] ), .S0(n7599), .S1(n7830), 
        .Y(n7080) );
  MX4X1 U6984 ( .A(\registers[768][7] ), .B(\registers[769][7] ), .C(
        \registers[770][7] ), .D(\registers[771][7] ), .S0(n7601), .S1(n7832), 
        .Y(n7111) );
  MX4X1 U6985 ( .A(\registers[816][7] ), .B(\registers[817][7] ), .C(
        \registers[818][7] ), .D(\registers[819][7] ), .S0(n7600), .S1(n7831), 
        .Y(n7096) );
  MX4X1 U6986 ( .A(\registers[800][7] ), .B(\registers[801][7] ), .C(
        \registers[802][7] ), .D(\registers[803][7] ), .S0(n7601), .S1(n7831), 
        .Y(n7101) );
  MX4X1 U6987 ( .A(\registers[960][7] ), .B(\registers[961][7] ), .C(
        \registers[962][7] ), .D(\registers[963][7] ), .S0(n7597), .S1(n7828), 
        .Y(n7048) );
  MX4X1 U6988 ( .A(\registers[1008][7] ), .B(\registers[1009][7] ), .C(
        \registers[1010][7] ), .D(\registers[1011][7] ), .S0(n7596), .S1(n7827), .Y(n7033) );
  MX4X1 U6989 ( .A(\registers[992][7] ), .B(\registers[993][7] ), .C(
        \registers[994][7] ), .D(\registers[995][7] ), .S0(n7597), .S1(n7827), 
        .Y(n7038) );
  MX4X1 U6990 ( .A(\registers[896][7] ), .B(\registers[897][7] ), .C(
        \registers[898][7] ), .D(\registers[899][7] ), .S0(n7599), .S1(n7829), 
        .Y(n7069) );
  MX4X1 U6991 ( .A(\registers[944][7] ), .B(\registers[945][7] ), .C(
        \registers[946][7] ), .D(\registers[947][7] ), .S0(n7598), .S1(n7828), 
        .Y(n7054) );
  MX4X1 U6992 ( .A(\registers[928][7] ), .B(\registers[929][7] ), .C(
        \registers[930][7] ), .D(\registers[931][7] ), .S0(n7598), .S1(n7829), 
        .Y(n7059) );
  MX4X1 U6993 ( .A(\registers[576][7] ), .B(\registers[577][7] ), .C(
        \registers[578][7] ), .D(\registers[579][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7175) );
  MX4X1 U6994 ( .A(\registers[624][7] ), .B(\registers[625][7] ), .C(
        \registers[626][7] ), .D(\registers[627][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7160) );
  MX4X1 U6995 ( .A(\registers[608][7] ), .B(\registers[609][7] ), .C(
        \registers[610][7] ), .D(\registers[611][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7165) );
  MX4X1 U6996 ( .A(\registers[512][7] ), .B(\registers[513][7] ), .C(
        \registers[514][7] ), .D(\registers[515][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7196) );
  MX4X1 U6997 ( .A(\registers[560][7] ), .B(\registers[561][7] ), .C(
        \registers[562][7] ), .D(\registers[563][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7181) );
  MX4X1 U6998 ( .A(\registers[544][7] ), .B(\registers[545][7] ), .C(
        \registers[546][7] ), .D(\registers[547][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7186) );
  MX4X1 U6999 ( .A(\registers[704][7] ), .B(\registers[705][7] ), .C(
        \registers[706][7] ), .D(\registers[707][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7133) );
  MX4X1 U7000 ( .A(\registers[752][7] ), .B(\registers[753][7] ), .C(
        \registers[754][7] ), .D(\registers[755][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7118) );
  MX4X1 U7001 ( .A(\registers[736][7] ), .B(\registers[737][7] ), .C(
        \registers[738][7] ), .D(\registers[739][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7123) );
  MX4X1 U7002 ( .A(\registers[640][7] ), .B(\registers[641][7] ), .C(
        \registers[642][7] ), .D(\registers[643][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7154) );
  MX4X1 U7003 ( .A(\registers[688][7] ), .B(\registers[689][7] ), .C(
        \registers[690][7] ), .D(\registers[691][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7139) );
  MX4X1 U7004 ( .A(\registers[672][7] ), .B(\registers[673][7] ), .C(
        \registers[674][7] ), .D(\registers[675][7] ), .S0(n7603), .S1(n7834), 
        .Y(n7144) );
  MX4X1 U7005 ( .A(n3256), .B(n3254), .C(n3255), .D(n3253), .S0(n4613), .S1(
        n4552), .Y(n3257) );
  MX4X1 U7006 ( .A(\registers[264][5] ), .B(\registers[265][5] ), .C(
        \registers[266][5] ), .D(\registers[267][5] ), .S0(n4226), .S1(n4459), 
        .Y(n3254) );
  MX4X1 U7007 ( .A(\registers[268][5] ), .B(\registers[269][5] ), .C(
        \registers[270][5] ), .D(\registers[271][5] ), .S0(n4226), .S1(n4459), 
        .Y(n3253) );
  MX4X1 U7008 ( .A(\registers[256][5] ), .B(\registers[257][5] ), .C(
        \registers[258][5] ), .D(\registers[259][5] ), .S0(n4226), .S1(n4459), 
        .Y(n3256) );
  MX4X1 U7009 ( .A(n3193), .B(n3191), .C(n3192), .D(n3190), .S0(n4612), .S1(
        n4551), .Y(n3194) );
  MX4X1 U7010 ( .A(\registers[456][5] ), .B(\registers[457][5] ), .C(
        \registers[458][5] ), .D(\registers[459][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3191) );
  MX4X1 U7011 ( .A(\registers[460][5] ), .B(\registers[461][5] ), .C(
        \registers[462][5] ), .D(\registers[463][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3190) );
  MX4X1 U7012 ( .A(\registers[448][5] ), .B(\registers[449][5] ), .C(
        \registers[450][5] ), .D(\registers[451][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3193) );
  MX4X1 U7013 ( .A(n3214), .B(n3212), .C(n3213), .D(n3211), .S0(n4613), .S1(
        n4552), .Y(n3215) );
  MX4X1 U7014 ( .A(\registers[392][5] ), .B(\registers[393][5] ), .C(
        \registers[394][5] ), .D(\registers[395][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3212) );
  MX4X1 U7015 ( .A(\registers[396][5] ), .B(\registers[397][5] ), .C(
        \registers[398][5] ), .D(\registers[399][5] ), .S0(n4224), .S1(n4456), 
        .Y(n3211) );
  MX4X1 U7016 ( .A(\registers[384][5] ), .B(\registers[385][5] ), .C(
        \registers[386][5] ), .D(\registers[387][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3214) );
  MX4X1 U7017 ( .A(n3596), .B(n3594), .C(n3595), .D(n3593), .S0(n4619), .S1(
        n4557), .Y(n3597) );
  MX4X1 U7018 ( .A(\registers[264][6] ), .B(\registers[265][6] ), .C(
        \registers[266][6] ), .D(\registers[267][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3594) );
  MX4X1 U7019 ( .A(\registers[268][6] ), .B(\registers[269][6] ), .C(
        \registers[270][6] ), .D(\registers[271][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3593) );
  MX4X1 U7020 ( .A(\registers[256][6] ), .B(\registers[257][6] ), .C(
        \registers[258][6] ), .D(\registers[259][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3596) );
  MX4X1 U7021 ( .A(n3533), .B(n3531), .C(n3532), .D(n3530), .S0(n4618), .S1(
        n4556), .Y(n3534) );
  MX4X1 U7022 ( .A(\registers[456][6] ), .B(\registers[457][6] ), .C(
        \registers[458][6] ), .D(\registers[459][6] ), .S0(n4244), .S1(n4475), 
        .Y(n3531) );
  MX4X1 U7023 ( .A(\registers[460][6] ), .B(\registers[461][6] ), .C(
        \registers[462][6] ), .D(\registers[463][6] ), .S0(n4244), .S1(n4475), 
        .Y(n3530) );
  MX4X1 U7024 ( .A(\registers[448][6] ), .B(\registers[449][6] ), .C(
        \registers[450][6] ), .D(\registers[451][6] ), .S0(n4244), .S1(n4475), 
        .Y(n3533) );
  MX4X1 U7025 ( .A(n3554), .B(n3552), .C(n3553), .D(n3551), .S0(n4618), .S1(
        n4557), .Y(n3555) );
  MX4X1 U7026 ( .A(\registers[392][6] ), .B(\registers[393][6] ), .C(
        \registers[394][6] ), .D(\registers[395][6] ), .S0(n4245), .S1(n4476), 
        .Y(n3552) );
  MX4X1 U7027 ( .A(\registers[396][6] ), .B(\registers[397][6] ), .C(
        \registers[398][6] ), .D(\registers[399][6] ), .S0(n4245), .S1(n4476), 
        .Y(n3551) );
  MX4X1 U7028 ( .A(\registers[384][6] ), .B(\registers[385][6] ), .C(
        \registers[386][6] ), .D(\registers[387][6] ), .S0(n4245), .S1(n4476), 
        .Y(n3554) );
  MX4X1 U7029 ( .A(n3936), .B(n3934), .C(n3935), .D(n3933), .S0(n4624), .S1(
        n4558), .Y(n3937) );
  MX4X1 U7030 ( .A(\registers[264][7] ), .B(\registers[265][7] ), .C(
        \registers[266][7] ), .D(\registers[267][7] ), .S0(n4269), .S1(n4497), 
        .Y(n3934) );
  MX4X1 U7031 ( .A(\registers[268][7] ), .B(\registers[269][7] ), .C(
        \registers[270][7] ), .D(\registers[271][7] ), .S0(n4269), .S1(n4497), 
        .Y(n3933) );
  MX4X1 U7032 ( .A(\registers[256][7] ), .B(\registers[257][7] ), .C(
        \registers[258][7] ), .D(\registers[259][7] ), .S0(n4269), .S1(n4498), 
        .Y(n3936) );
  MX4X1 U7033 ( .A(n3873), .B(n3871), .C(n3872), .D(n3870), .S0(n4623), .S1(
        n4526), .Y(n3874) );
  MX4X1 U7034 ( .A(\registers[456][7] ), .B(\registers[457][7] ), .C(
        \registers[458][7] ), .D(\registers[459][7] ), .S0(n4265), .S1(n4495), 
        .Y(n3871) );
  MX4X1 U7035 ( .A(\registers[460][7] ), .B(\registers[461][7] ), .C(
        \registers[462][7] ), .D(\registers[463][7] ), .S0(n4265), .S1(n4495), 
        .Y(n3870) );
  MX4X1 U7036 ( .A(\registers[448][7] ), .B(\registers[449][7] ), .C(
        \registers[450][7] ), .D(\registers[451][7] ), .S0(n4265), .S1(n4495), 
        .Y(n3873) );
  MX4X1 U7037 ( .A(n3894), .B(n3892), .C(n3893), .D(n3891), .S0(n4623), .S1(
        n4558), .Y(n3895) );
  MX4X1 U7038 ( .A(\registers[392][7] ), .B(\registers[393][7] ), .C(
        \registers[394][7] ), .D(\registers[395][7] ), .S0(n4266), .S1(n4496), 
        .Y(n3892) );
  MX4X1 U7039 ( .A(\registers[396][7] ), .B(\registers[397][7] ), .C(
        \registers[398][7] ), .D(\registers[399][7] ), .S0(n4266), .S1(n4496), 
        .Y(n3891) );
  MX4X1 U7040 ( .A(\registers[384][7] ), .B(\registers[385][7] ), .C(
        \registers[386][7] ), .D(\registers[387][7] ), .S0(n4266), .S1(n4496), 
        .Y(n3894) );
  MX4X1 U7041 ( .A(n4901), .B(n4899), .C(n4900), .D(n4898), .S0(n7930), .S1(
        n7870), .Y(n4902) );
  MX4X1 U7042 ( .A(\registers[264][0] ), .B(\registers[265][0] ), .C(
        \registers[266][0] ), .D(\registers[267][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4899) );
  MX4X1 U7043 ( .A(\registers[268][0] ), .B(\registers[269][0] ), .C(
        \registers[270][0] ), .D(\registers[271][0] ), .S0(n7463), .S1(n7704), 
        .Y(n4898) );
  MX4X1 U7044 ( .A(\registers[256][0] ), .B(\registers[257][0] ), .C(
        \registers[258][0] ), .D(\registers[259][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4901) );
  MX4X1 U7045 ( .A(n4838), .B(n4836), .C(n4837), .D(n4835), .S0(n7955), .S1(
        n7869), .Y(n4839) );
  MX4X1 U7046 ( .A(\registers[456][0] ), .B(\registers[457][0] ), .C(
        \registers[458][0] ), .D(\registers[459][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4836) );
  MX4X1 U7047 ( .A(\registers[460][0] ), .B(\registers[461][0] ), .C(
        \registers[462][0] ), .D(\registers[463][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4835) );
  MX4X1 U7048 ( .A(\registers[448][0] ), .B(\registers[449][0] ), .C(
        \registers[450][0] ), .D(\registers[451][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4838) );
  MX4X1 U7049 ( .A(n4859), .B(n4857), .C(n4858), .D(n4856), .S0(n7934), .S1(
        n7869), .Y(n4860) );
  MX4X1 U7050 ( .A(\registers[392][0] ), .B(\registers[393][0] ), .C(
        \registers[394][0] ), .D(\registers[395][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4857) );
  MX4X1 U7051 ( .A(\registers[396][0] ), .B(\registers[397][0] ), .C(
        \registers[398][0] ), .D(\registers[399][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4856) );
  MX4X1 U7052 ( .A(\registers[384][0] ), .B(\registers[385][0] ), .C(
        \registers[386][0] ), .D(\registers[387][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4859) );
  MX4X1 U7053 ( .A(n5241), .B(n5239), .C(n5240), .D(n5238), .S0(n7935), .S1(
        n7875), .Y(n5242) );
  MX4X1 U7054 ( .A(\registers[264][1] ), .B(\registers[265][1] ), .C(
        \registers[266][1] ), .D(\registers[267][1] ), .S0(n7484), .S1(n7724), 
        .Y(n5239) );
  MX4X1 U7055 ( .A(\registers[268][1] ), .B(\registers[269][1] ), .C(
        \registers[270][1] ), .D(\registers[271][1] ), .S0(n7484), .S1(n7724), 
        .Y(n5238) );
  MX4X1 U7056 ( .A(\registers[256][1] ), .B(\registers[257][1] ), .C(
        \registers[258][1] ), .D(\registers[259][1] ), .S0(n7484), .S1(n7724), 
        .Y(n5241) );
  MX4X1 U7057 ( .A(n5178), .B(n5176), .C(n5177), .D(n5175), .S0(n7934), .S1(
        n7874), .Y(n5179) );
  MX4X1 U7058 ( .A(\registers[456][1] ), .B(\registers[457][1] ), .C(
        \registers[458][1] ), .D(\registers[459][1] ), .S0(n7480), .S1(n7721), 
        .Y(n5176) );
  MX4X1 U7059 ( .A(\registers[460][1] ), .B(\registers[461][1] ), .C(
        \registers[462][1] ), .D(\registers[463][1] ), .S0(n7480), .S1(n7720), 
        .Y(n5175) );
  MX4X1 U7060 ( .A(\registers[448][1] ), .B(\registers[449][1] ), .C(
        \registers[450][1] ), .D(\registers[451][1] ), .S0(n7480), .S1(n7721), 
        .Y(n5178) );
  MX4X1 U7061 ( .A(n5199), .B(n5197), .C(n5198), .D(n5196), .S0(n7934), .S1(
        n7874), .Y(n5200) );
  MX4X1 U7062 ( .A(\registers[392][1] ), .B(\registers[393][1] ), .C(
        \registers[394][1] ), .D(\registers[395][1] ), .S0(n7481), .S1(n7722), 
        .Y(n5197) );
  MX4X1 U7063 ( .A(\registers[396][1] ), .B(\registers[397][1] ), .C(
        \registers[398][1] ), .D(\registers[399][1] ), .S0(n7481), .S1(n7722), 
        .Y(n5196) );
  MX4X1 U7064 ( .A(\registers[384][1] ), .B(\registers[385][1] ), .C(
        \registers[386][1] ), .D(\registers[387][1] ), .S0(n7481), .S1(n7722), 
        .Y(n5199) );
  MX4X1 U7065 ( .A(n5581), .B(n5579), .C(n5580), .D(n5578), .S0(n7940), .S1(
        n7880), .Y(n5582) );
  MX4X1 U7066 ( .A(\registers[264][2] ), .B(\registers[265][2] ), .C(
        \registers[266][2] ), .D(\registers[267][2] ), .S0(n7505), .S1(n7744), 
        .Y(n5579) );
  MX4X1 U7067 ( .A(\registers[268][2] ), .B(\registers[269][2] ), .C(
        \registers[270][2] ), .D(\registers[271][2] ), .S0(n7505), .S1(n7744), 
        .Y(n5578) );
  MX4X1 U7068 ( .A(\registers[256][2] ), .B(\registers[257][2] ), .C(
        \registers[258][2] ), .D(\registers[259][2] ), .S0(n7505), .S1(n7744), 
        .Y(n5581) );
  MX4X1 U7069 ( .A(n5518), .B(n5516), .C(n5517), .D(n5515), .S0(n7939), .S1(
        n7879), .Y(n5519) );
  MX4X1 U7070 ( .A(\registers[456][2] ), .B(\registers[457][2] ), .C(
        \registers[458][2] ), .D(\registers[459][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5516) );
  MX4X1 U7071 ( .A(\registers[460][2] ), .B(\registers[461][2] ), .C(
        \registers[462][2] ), .D(\registers[463][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5515) );
  MX4X1 U7072 ( .A(\registers[448][2] ), .B(\registers[449][2] ), .C(
        \registers[450][2] ), .D(\registers[451][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5518) );
  MX4X1 U7073 ( .A(n5539), .B(n5537), .C(n5538), .D(n5536), .S0(n7940), .S1(
        n7879), .Y(n5540) );
  MX4X1 U7074 ( .A(\registers[392][2] ), .B(\registers[393][2] ), .C(
        \registers[394][2] ), .D(\registers[395][2] ), .S0(n7503), .S1(n7741), 
        .Y(n5537) );
  MX4X1 U7075 ( .A(\registers[396][2] ), .B(\registers[397][2] ), .C(
        \registers[398][2] ), .D(\registers[399][2] ), .S0(n7503), .S1(n7741), 
        .Y(n5536) );
  MX4X1 U7076 ( .A(\registers[384][2] ), .B(\registers[385][2] ), .C(
        \registers[386][2] ), .D(\registers[387][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5539) );
  MX4X1 U7077 ( .A(n5921), .B(n5919), .C(n5920), .D(n5918), .S0(n7946), .S1(
        n7885), .Y(n5922) );
  MX4X1 U7078 ( .A(\registers[264][3] ), .B(\registers[265][3] ), .C(
        \registers[266][3] ), .D(\registers[267][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5919) );
  MX4X1 U7079 ( .A(\registers[268][3] ), .B(\registers[269][3] ), .C(
        \registers[270][3] ), .D(\registers[271][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5918) );
  MX4X1 U7080 ( .A(\registers[256][3] ), .B(\registers[257][3] ), .C(
        \registers[258][3] ), .D(\registers[259][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5921) );
  MX4X1 U7081 ( .A(n5858), .B(n5856), .C(n5857), .D(n5855), .S0(n7945), .S1(
        n7884), .Y(n5859) );
  MX4X1 U7082 ( .A(\registers[456][3] ), .B(\registers[457][3] ), .C(
        \registers[458][3] ), .D(\registers[459][3] ), .S0(n7523), .S1(n7760), 
        .Y(n5856) );
  MX4X1 U7083 ( .A(\registers[460][3] ), .B(\registers[461][3] ), .C(
        \registers[462][3] ), .D(\registers[463][3] ), .S0(n7523), .S1(n7760), 
        .Y(n5855) );
  MX4X1 U7084 ( .A(\registers[448][3] ), .B(\registers[449][3] ), .C(
        \registers[450][3] ), .D(\registers[451][3] ), .S0(n7523), .S1(n7760), 
        .Y(n5858) );
  MX4X1 U7085 ( .A(n5879), .B(n5877), .C(n5878), .D(n5876), .S0(n7945), .S1(
        n7884), .Y(n5880) );
  MX4X1 U7086 ( .A(\registers[392][3] ), .B(\registers[393][3] ), .C(
        \registers[394][3] ), .D(\registers[395][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5877) );
  MX4X1 U7087 ( .A(\registers[396][3] ), .B(\registers[397][3] ), .C(
        \registers[398][3] ), .D(\registers[399][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5876) );
  MX4X1 U7088 ( .A(\registers[384][3] ), .B(\registers[385][3] ), .C(
        \registers[386][3] ), .D(\registers[387][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5879) );
  MX4X1 U7089 ( .A(n6261), .B(n6259), .C(n6260), .D(n6258), .S0(n7951), .S1(
        n7889), .Y(n6262) );
  MX4X1 U7090 ( .A(\registers[264][4] ), .B(\registers[265][4] ), .C(
        \registers[266][4] ), .D(\registers[267][4] ), .S0(n7548), .S1(n7783), 
        .Y(n6259) );
  MX4X1 U7091 ( .A(\registers[268][4] ), .B(\registers[269][4] ), .C(
        \registers[270][4] ), .D(\registers[271][4] ), .S0(n7548), .S1(n7783), 
        .Y(n6258) );
  MX4X1 U7092 ( .A(\registers[256][4] ), .B(\registers[257][4] ), .C(
        \registers[258][4] ), .D(\registers[259][4] ), .S0(n7548), .S1(n7783), 
        .Y(n6261) );
  MX4X1 U7093 ( .A(n6198), .B(n6196), .C(n6197), .D(n6195), .S0(n7950), .S1(
        n7889), .Y(n6199) );
  MX4X1 U7094 ( .A(\registers[456][4] ), .B(\registers[457][4] ), .C(
        \registers[458][4] ), .D(\registers[459][4] ), .S0(n7544), .S1(n7780), 
        .Y(n6196) );
  MX4X1 U7095 ( .A(\registers[460][4] ), .B(\registers[461][4] ), .C(
        \registers[462][4] ), .D(\registers[463][4] ), .S0(n7544), .S1(n7780), 
        .Y(n6195) );
  MX4X1 U7096 ( .A(\registers[448][4] ), .B(\registers[449][4] ), .C(
        \registers[450][4] ), .D(\registers[451][4] ), .S0(n7544), .S1(n7780), 
        .Y(n6198) );
  MX4X1 U7097 ( .A(n6219), .B(n6217), .C(n6218), .D(n6216), .S0(n7950), .S1(
        n7889), .Y(n6220) );
  MX4X1 U7098 ( .A(\registers[392][4] ), .B(\registers[393][4] ), .C(
        \registers[394][4] ), .D(\registers[395][4] ), .S0(n7545), .S1(n7781), 
        .Y(n6217) );
  MX4X1 U7099 ( .A(\registers[396][4] ), .B(\registers[397][4] ), .C(
        \registers[398][4] ), .D(\registers[399][4] ), .S0(n7545), .S1(n7781), 
        .Y(n6216) );
  MX4X1 U7100 ( .A(\registers[384][4] ), .B(\registers[385][4] ), .C(
        \registers[386][4] ), .D(\registers[387][4] ), .S0(n7545), .S1(n7781), 
        .Y(n6219) );
  MX4X1 U7101 ( .A(n6601), .B(n6599), .C(n6600), .D(n6598), .S0(n7956), .S1(
        n7894), .Y(n6602) );
  MX4X1 U7102 ( .A(\registers[264][5] ), .B(\registers[265][5] ), .C(
        \registers[266][5] ), .D(\registers[267][5] ), .S0(n7569), .S1(n7803), 
        .Y(n6599) );
  MX4X1 U7103 ( .A(\registers[268][5] ), .B(\registers[269][5] ), .C(
        \registers[270][5] ), .D(\registers[271][5] ), .S0(n7569), .S1(n7803), 
        .Y(n6598) );
  MX4X1 U7104 ( .A(\registers[256][5] ), .B(\registers[257][5] ), .C(
        \registers[258][5] ), .D(\registers[259][5] ), .S0(n7569), .S1(n7803), 
        .Y(n6601) );
  MX4X1 U7105 ( .A(n6538), .B(n6536), .C(n6537), .D(n6535), .S0(n7955), .S1(
        n7893), .Y(n6539) );
  MX4X1 U7106 ( .A(\registers[456][5] ), .B(\registers[457][5] ), .C(
        \registers[458][5] ), .D(\registers[459][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6536) );
  MX4X1 U7107 ( .A(\registers[460][5] ), .B(\registers[461][5] ), .C(
        \registers[462][5] ), .D(\registers[463][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6535) );
  MX4X1 U7108 ( .A(\registers[448][5] ), .B(\registers[449][5] ), .C(
        \registers[450][5] ), .D(\registers[451][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6538) );
  MX4X1 U7109 ( .A(n6559), .B(n6557), .C(n6558), .D(n6556), .S0(n7956), .S1(
        n7894), .Y(n6560) );
  MX4X1 U7110 ( .A(\registers[392][5] ), .B(\registers[393][5] ), .C(
        \registers[394][5] ), .D(\registers[395][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6557) );
  MX4X1 U7111 ( .A(\registers[396][5] ), .B(\registers[397][5] ), .C(
        \registers[398][5] ), .D(\registers[399][5] ), .S0(n7567), .S1(n7800), 
        .Y(n6556) );
  MX4X1 U7112 ( .A(\registers[384][5] ), .B(\registers[385][5] ), .C(
        \registers[386][5] ), .D(\registers[387][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6559) );
  MX4X1 U7113 ( .A(n6941), .B(n6939), .C(n6940), .D(n6938), .S0(n7962), .S1(
        n7897), .Y(n6942) );
  MX4X1 U7114 ( .A(\registers[264][6] ), .B(\registers[265][6] ), .C(
        \registers[266][6] ), .D(\registers[267][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6939) );
  MX4X1 U7115 ( .A(\registers[268][6] ), .B(\registers[269][6] ), .C(
        \registers[270][6] ), .D(\registers[271][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6938) );
  MX4X1 U7116 ( .A(\registers[256][6] ), .B(\registers[257][6] ), .C(
        \registers[258][6] ), .D(\registers[259][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6941) );
  MX4X1 U7117 ( .A(n6878), .B(n6876), .C(n6877), .D(n6875), .S0(n7961), .S1(
        n7893), .Y(n6879) );
  MX4X1 U7118 ( .A(\registers[456][6] ), .B(\registers[457][6] ), .C(
        \registers[458][6] ), .D(\registers[459][6] ), .S0(n7587), .S1(n7818), 
        .Y(n6876) );
  MX4X1 U7119 ( .A(\registers[460][6] ), .B(\registers[461][6] ), .C(
        \registers[462][6] ), .D(\registers[463][6] ), .S0(n7587), .S1(n7818), 
        .Y(n6875) );
  MX4X1 U7120 ( .A(\registers[448][6] ), .B(\registers[449][6] ), .C(
        \registers[450][6] ), .D(\registers[451][6] ), .S0(n7587), .S1(n7818), 
        .Y(n6878) );
  MX4X1 U7121 ( .A(n6899), .B(n6897), .C(n6898), .D(n6896), .S0(n7961), .S1(
        n7897), .Y(n6900) );
  MX4X1 U7122 ( .A(\registers[392][6] ), .B(\registers[393][6] ), .C(
        \registers[394][6] ), .D(\registers[395][6] ), .S0(n7588), .S1(n7819), 
        .Y(n6897) );
  MX4X1 U7123 ( .A(\registers[396][6] ), .B(\registers[397][6] ), .C(
        \registers[398][6] ), .D(\registers[399][6] ), .S0(n7588), .S1(n7819), 
        .Y(n6896) );
  MX4X1 U7124 ( .A(\registers[384][6] ), .B(\registers[385][6] ), .C(
        \registers[386][6] ), .D(\registers[387][6] ), .S0(n7588), .S1(n7819), 
        .Y(n6899) );
  MX4X1 U7125 ( .A(n7218), .B(n7216), .C(n7217), .D(n7215), .S0(n7966), .S1(
        n7901), .Y(n7219) );
  MX4X1 U7126 ( .A(\registers[456][7] ), .B(\registers[457][7] ), .C(
        \registers[458][7] ), .D(\registers[459][7] ), .S0(n7608), .S1(n7838), 
        .Y(n7216) );
  MX4X1 U7127 ( .A(\registers[460][7] ), .B(\registers[461][7] ), .C(
        \registers[462][7] ), .D(\registers[463][7] ), .S0(n7608), .S1(n7838), 
        .Y(n7215) );
  MX4X1 U7128 ( .A(\registers[448][7] ), .B(\registers[449][7] ), .C(
        \registers[450][7] ), .D(\registers[451][7] ), .S0(n7608), .S1(n7838), 
        .Y(n7218) );
  MX4X1 U7129 ( .A(n7239), .B(n7237), .C(n7238), .D(n7236), .S0(n7966), .S1(
        n7902), .Y(n7240) );
  MX4X1 U7130 ( .A(\registers[392][7] ), .B(\registers[393][7] ), .C(
        \registers[394][7] ), .D(\registers[395][7] ), .S0(n7609), .S1(n7839), 
        .Y(n7237) );
  MX4X1 U7131 ( .A(\registers[396][7] ), .B(\registers[397][7] ), .C(
        \registers[398][7] ), .D(\registers[399][7] ), .S0(n7609), .S1(n7839), 
        .Y(n7236) );
  MX4X1 U7132 ( .A(\registers[384][7] ), .B(\registers[385][7] ), .C(
        \registers[386][7] ), .D(\registers[387][7] ), .S0(n7609), .S1(n7839), 
        .Y(n7239) );
  MX4X1 U7133 ( .A(n7281), .B(n7279), .C(n7280), .D(n7278), .S0(n7967), .S1(
        n7898), .Y(n7282) );
  MX4X1 U7134 ( .A(\registers[264][7] ), .B(\registers[265][7] ), .C(
        \registers[266][7] ), .D(\registers[267][7] ), .S0(n7612), .S1(n7841), 
        .Y(n7279) );
  MX4X1 U7135 ( .A(\registers[268][7] ), .B(\registers[269][7] ), .C(
        \registers[270][7] ), .D(\registers[271][7] ), .S0(n7612), .S1(n7841), 
        .Y(n7278) );
  MX4X1 U7136 ( .A(\registers[256][7] ), .B(\registers[257][7] ), .C(
        \registers[258][7] ), .D(\registers[259][7] ), .S0(n7612), .S1(n7842), 
        .Y(n7281) );
  MX4X1 U7137 ( .A(\registers[1020][0] ), .B(\registers[1021][0] ), .C(
        \registers[1022][0] ), .D(\registers[1023][0] ), .S0(n4105), .S1(n4349), .Y(n1045) );
  MX4X1 U7138 ( .A(\registers[1004][0] ), .B(\registers[1005][0] ), .C(
        \registers[1006][0] ), .D(\registers[1007][0] ), .S0(n4231), .S1(n4349), .Y(n1050) );
  MX4X1 U7139 ( .A(\registers[1020][0] ), .B(\registers[1021][0] ), .C(
        \registers[1022][0] ), .D(\registers[1023][0] ), .S0(n7575), .S1(n7807), .Y(n4650) );
  MX4X1 U7140 ( .A(\registers[1004][0] ), .B(\registers[1005][0] ), .C(
        \registers[1006][0] ), .D(\registers[1007][0] ), .S0(n7556), .S1(n7805), .Y(n4655) );
  MX4X1 U7141 ( .A(\registers[332][0] ), .B(\registers[333][0] ), .C(
        \registers[334][0] ), .D(\registers[335][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1428) );
  MX4X1 U7142 ( .A(\registers[380][0] ), .B(\registers[381][0] ), .C(
        \registers[382][0] ), .D(\registers[383][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1413) );
  MX4X1 U7143 ( .A(\registers[364][0] ), .B(\registers[365][0] ), .C(
        \registers[366][0] ), .D(\registers[367][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1418) );
  MX4X1 U7144 ( .A(\registers[76][0] ), .B(\registers[77][0] ), .C(
        \registers[78][0] ), .D(\registers[79][0] ), .S0(n4124), .S1(n4364), 
        .Y(n1519) );
  MX4X1 U7145 ( .A(\registers[124][0] ), .B(\registers[125][0] ), .C(
        \registers[126][0] ), .D(\registers[127][0] ), .S0(n4123), .S1(n4363), 
        .Y(n1502) );
  MX4X1 U7146 ( .A(\registers[108][0] ), .B(\registers[109][0] ), .C(
        \registers[110][0] ), .D(\registers[111][0] ), .S0(n4123), .S1(n4364), 
        .Y(n1509) );
  MX4X1 U7147 ( .A(\registers[12][0] ), .B(\registers[13][0] ), .C(
        \registers[14][0] ), .D(\registers[15][0] ), .S0(n4125), .S1(n4365), 
        .Y(n1542) );
  MX4X1 U7148 ( .A(\registers[60][0] ), .B(\registers[61][0] ), .C(
        \registers[62][0] ), .D(\registers[63][0] ), .S0(n4124), .S1(n4364), 
        .Y(n1525) );
  MX4X1 U7149 ( .A(\registers[44][0] ), .B(\registers[45][0] ), .C(
        \registers[46][0] ), .D(\registers[47][0] ), .S0(n4124), .S1(n4365), 
        .Y(n1530) );
  MX4X1 U7150 ( .A(\registers[204][0] ), .B(\registers[205][0] ), .C(
        \registers[206][0] ), .D(\registers[207][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1475) );
  MX4X1 U7151 ( .A(\registers[252][0] ), .B(\registers[253][0] ), .C(
        \registers[254][0] ), .D(\registers[255][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1458) );
  MX4X1 U7152 ( .A(\registers[236][0] ), .B(\registers[237][0] ), .C(
        \registers[238][0] ), .D(\registers[239][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1463) );
  MX4X1 U7153 ( .A(\registers[140][0] ), .B(\registers[141][0] ), .C(
        \registers[142][0] ), .D(\registers[143][0] ), .S0(n4122), .S1(n4363), 
        .Y(n1496) );
  MX4X1 U7154 ( .A(\registers[188][0] ), .B(\registers[189][0] ), .C(
        \registers[190][0] ), .D(\registers[191][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1481) );
  MX4X1 U7155 ( .A(\registers[172][0] ), .B(\registers[173][0] ), .C(
        \registers[174][0] ), .D(\registers[175][0] ), .S0(n4122), .S1(n4362), 
        .Y(n1486) );
  MX4X1 U7156 ( .A(\registers[844][0] ), .B(\registers[845][0] ), .C(
        \registers[846][0] ), .D(\registers[847][0] ), .S0(n4108), .S1(n4485), 
        .Y(n1102) );
  MX4X1 U7157 ( .A(\registers[892][0] ), .B(\registers[893][0] ), .C(
        \registers[894][0] ), .D(\registers[895][0] ), .S0(n4107), .S1(n4350), 
        .Y(n1087) );
  MX4X1 U7158 ( .A(\registers[876][0] ), .B(\registers[877][0] ), .C(
        \registers[878][0] ), .D(\registers[879][0] ), .S0(n4107), .S1(n4494), 
        .Y(n1092) );
  MX4X1 U7159 ( .A(\registers[780][0] ), .B(\registers[781][0] ), .C(
        \registers[782][0] ), .D(\registers[783][0] ), .S0(n4109), .S1(n4351), 
        .Y(n1165) );
  MX4X1 U7160 ( .A(\registers[828][0] ), .B(\registers[829][0] ), .C(
        \registers[830][0] ), .D(\registers[831][0] ), .S0(n4108), .S1(n4501), 
        .Y(n1150) );
  MX4X1 U7161 ( .A(\registers[812][0] ), .B(\registers[813][0] ), .C(
        \registers[814][0] ), .D(\registers[815][0] ), .S0(n4108), .S1(n4464), 
        .Y(n1155) );
  MX4X1 U7162 ( .A(\registers[972][0] ), .B(\registers[973][0] ), .C(
        \registers[974][0] ), .D(\registers[975][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1060) );
  MX4X1 U7163 ( .A(\registers[908][0] ), .B(\registers[909][0] ), .C(
        \registers[910][0] ), .D(\registers[911][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1081) );
  MX4X1 U7164 ( .A(\registers[956][0] ), .B(\registers[957][0] ), .C(
        \registers[958][0] ), .D(\registers[959][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1066) );
  MX4X1 U7165 ( .A(\registers[940][0] ), .B(\registers[941][0] ), .C(
        \registers[942][0] ), .D(\registers[943][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1071) );
  MX4X1 U7166 ( .A(\registers[588][0] ), .B(\registers[589][0] ), .C(
        \registers[590][0] ), .D(\registers[591][0] ), .S0(n4113), .S1(n4354), 
        .Y(n1338) );
  MX4X1 U7167 ( .A(\registers[636][0] ), .B(\registers[637][0] ), .C(
        \registers[638][0] ), .D(\registers[639][0] ), .S0(n4112), .S1(n4353), 
        .Y(n1311) );
  MX4X1 U7168 ( .A(\registers[620][0] ), .B(\registers[621][0] ), .C(
        \registers[622][0] ), .D(\registers[623][0] ), .S0(n4112), .S1(n4354), 
        .Y(n1321) );
  MX4X1 U7169 ( .A(\registers[524][0] ), .B(\registers[525][0] ), .C(
        \registers[526][0] ), .D(\registers[527][0] ), .S0(n4114), .S1(n4356), 
        .Y(n1359) );
  MX4X1 U7170 ( .A(\registers[572][0] ), .B(\registers[573][0] ), .C(
        \registers[574][0] ), .D(\registers[575][0] ), .S0(n4113), .S1(n4355), 
        .Y(n1344) );
  MX4X1 U7171 ( .A(\registers[556][0] ), .B(\registers[557][0] ), .C(
        \registers[558][0] ), .D(\registers[559][0] ), .S0(n4114), .S1(n4355), 
        .Y(n1349) );
  MX4X1 U7172 ( .A(\registers[716][0] ), .B(\registers[717][0] ), .C(
        \registers[718][0] ), .D(\registers[719][0] ), .S0(n4110), .S1(n4352), 
        .Y(n1201) );
  MX4X1 U7173 ( .A(\registers[764][0] ), .B(\registers[765][0] ), .C(
        \registers[766][0] ), .D(\registers[767][0] ), .S0(n4109), .S1(n4351), 
        .Y(n1172) );
  MX4X1 U7174 ( .A(\registers[748][0] ), .B(\registers[749][0] ), .C(
        \registers[750][0] ), .D(\registers[751][0] ), .S0(n4110), .S1(n4351), 
        .Y(n1177) );
  MX4X1 U7175 ( .A(\registers[652][0] ), .B(\registers[653][0] ), .C(
        \registers[654][0] ), .D(\registers[655][0] ), .S0(n4112), .S1(n4353), 
        .Y(n1299) );
  MX4X1 U7176 ( .A(\registers[700][0] ), .B(\registers[701][0] ), .C(
        \registers[702][0] ), .D(\registers[703][0] ), .S0(n4111), .S1(n4352), 
        .Y(n1210) );
  MX4X1 U7177 ( .A(\registers[684][0] ), .B(\registers[685][0] ), .C(
        \registers[686][0] ), .D(\registers[687][0] ), .S0(n4111), .S1(n4352), 
        .Y(n1279) );
  MX4X1 U7178 ( .A(\registers[332][1] ), .B(\registers[333][1] ), .C(
        \registers[334][1] ), .D(\registers[335][1] ), .S0(n4140), .S1(n4379), 
        .Y(n1786) );
  MX4X1 U7179 ( .A(\registers[380][1] ), .B(\registers[381][1] ), .C(
        \registers[382][1] ), .D(\registers[383][1] ), .S0(n4139), .S1(n4378), 
        .Y(n1770) );
  MX4X1 U7180 ( .A(\registers[364][1] ), .B(\registers[365][1] ), .C(
        \registers[366][1] ), .D(\registers[367][1] ), .S0(n4139), .S1(n4378), 
        .Y(n1776) );
  MX4X1 U7181 ( .A(\registers[76][1] ), .B(\registers[77][1] ), .C(
        \registers[78][1] ), .D(\registers[79][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1875) );
  MX4X1 U7182 ( .A(\registers[124][1] ), .B(\registers[125][1] ), .C(
        \registers[126][1] ), .D(\registers[127][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1858) );
  MX4X1 U7183 ( .A(\registers[108][1] ), .B(\registers[109][1] ), .C(
        \registers[110][1] ), .D(\registers[111][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1863) );
  MX4X1 U7184 ( .A(\registers[12][1] ), .B(\registers[13][1] ), .C(
        \registers[14][1] ), .D(\registers[15][1] ), .S0(n4146), .S1(n4385), 
        .Y(n1896) );
  MX4X1 U7185 ( .A(\registers[60][1] ), .B(\registers[61][1] ), .C(
        \registers[62][1] ), .D(\registers[63][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1881) );
  MX4X1 U7186 ( .A(\registers[44][1] ), .B(\registers[45][1] ), .C(
        \registers[46][1] ), .D(\registers[47][1] ), .S0(n4146), .S1(n4384), 
        .Y(n1886) );
  MX4X1 U7187 ( .A(\registers[204][1] ), .B(\registers[205][1] ), .C(
        \registers[206][1] ), .D(\registers[207][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1830) );
  MX4X1 U7188 ( .A(\registers[252][1] ), .B(\registers[253][1] ), .C(
        \registers[254][1] ), .D(\registers[255][1] ), .S0(n4141), .S1(n4380), 
        .Y(n1815) );
  MX4X1 U7189 ( .A(\registers[236][1] ), .B(\registers[237][1] ), .C(
        \registers[238][1] ), .D(\registers[239][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1820) );
  MX4X1 U7190 ( .A(\registers[140][1] ), .B(\registers[141][1] ), .C(
        \registers[142][1] ), .D(\registers[143][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1852) );
  MX4X1 U7191 ( .A(\registers[188][1] ), .B(\registers[189][1] ), .C(
        \registers[190][1] ), .D(\registers[191][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1836) );
  MX4X1 U7192 ( .A(\registers[172][1] ), .B(\registers[173][1] ), .C(
        \registers[174][1] ), .D(\registers[175][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1842) );
  MX4X1 U7193 ( .A(\registers[844][1] ), .B(\registers[845][1] ), .C(
        \registers[846][1] ), .D(\registers[847][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1611) );
  MX4X1 U7194 ( .A(\registers[892][1] ), .B(\registers[893][1] ), .C(
        \registers[894][1] ), .D(\registers[895][1] ), .S0(n4128), .S1(n4368), 
        .Y(n1593) );
  MX4X1 U7195 ( .A(\registers[876][1] ), .B(\registers[877][1] ), .C(
        \registers[878][1] ), .D(\registers[879][1] ), .S0(n4128), .S1(n4368), 
        .Y(n1598) );
  MX4X1 U7196 ( .A(\registers[780][1] ), .B(\registers[781][1] ), .C(
        \registers[782][1] ), .D(\registers[783][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1632) );
  MX4X1 U7197 ( .A(\registers[828][1] ), .B(\registers[829][1] ), .C(
        \registers[830][1] ), .D(\registers[831][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1617) );
  MX4X1 U7198 ( .A(\registers[812][1] ), .B(\registers[813][1] ), .C(
        \registers[814][1] ), .D(\registers[815][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1622) );
  MX4X1 U7199 ( .A(\registers[972][1] ), .B(\registers[973][1] ), .C(
        \registers[974][1] ), .D(\registers[975][1] ), .S0(n4126), .S1(n4367), 
        .Y(n1564) );
  MX4X1 U7200 ( .A(\registers[1020][1] ), .B(\registers[1021][1] ), .C(
        \registers[1022][1] ), .D(\registers[1023][1] ), .S0(n4125), .S1(n4366), .Y(n1549) );
  MX4X1 U7201 ( .A(\registers[1004][1] ), .B(\registers[1005][1] ), .C(
        \registers[1006][1] ), .D(\registers[1007][1] ), .S0(n4126), .S1(n4366), .Y(n1554) );
  MX4X1 U7202 ( .A(\registers[908][1] ), .B(\registers[909][1] ), .C(
        \registers[910][1] ), .D(\registers[911][1] ), .S0(n4128), .S1(n4368), 
        .Y(n1587) );
  MX4X1 U7203 ( .A(\registers[956][1] ), .B(\registers[957][1] ), .C(
        \registers[958][1] ), .D(\registers[959][1] ), .S0(n4127), .S1(n4367), 
        .Y(n1570) );
  MX4X1 U7204 ( .A(\registers[940][1] ), .B(\registers[941][1] ), .C(
        \registers[942][1] ), .D(\registers[943][1] ), .S0(n4127), .S1(n4367), 
        .Y(n1577) );
  MX4X1 U7205 ( .A(\registers[588][1] ), .B(\registers[589][1] ), .C(
        \registers[590][1] ), .D(\registers[591][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1698) );
  MX4X1 U7206 ( .A(\registers[636][1] ), .B(\registers[637][1] ), .C(
        \registers[638][1] ), .D(\registers[639][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1683) );
  MX4X1 U7207 ( .A(\registers[620][1] ), .B(\registers[621][1] ), .C(
        \registers[622][1] ), .D(\registers[623][1] ), .S0(n4134), .S1(n4373), 
        .Y(n1688) );
  MX4X1 U7208 ( .A(\registers[524][1] ), .B(\registers[525][1] ), .C(
        \registers[526][1] ), .D(\registers[527][1] ), .S0(n4136), .S1(n4375), 
        .Y(n1720) );
  MX4X1 U7209 ( .A(\registers[572][1] ), .B(\registers[573][1] ), .C(
        \registers[574][1] ), .D(\registers[575][1] ), .S0(n4135), .S1(n4374), 
        .Y(n1704) );
  MX4X1 U7210 ( .A(\registers[556][1] ), .B(\registers[557][1] ), .C(
        \registers[558][1] ), .D(\registers[559][1] ), .S0(n4135), .S1(n4375), 
        .Y(n1710) );
  MX4X1 U7211 ( .A(\registers[716][1] ), .B(\registers[717][1] ), .C(
        \registers[718][1] ), .D(\registers[719][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1655) );
  MX4X1 U7212 ( .A(\registers[764][1] ), .B(\registers[765][1] ), .C(
        \registers[766][1] ), .D(\registers[767][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1639) );
  MX4X1 U7213 ( .A(\registers[748][1] ), .B(\registers[749][1] ), .C(
        \registers[750][1] ), .D(\registers[751][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1645) );
  MX4X1 U7214 ( .A(\registers[652][1] ), .B(\registers[653][1] ), .C(
        \registers[654][1] ), .D(\registers[655][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1677) );
  MX4X1 U7215 ( .A(\registers[700][1] ), .B(\registers[701][1] ), .C(
        \registers[702][1] ), .D(\registers[703][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1661) );
  MX4X1 U7216 ( .A(\registers[684][1] ), .B(\registers[685][1] ), .C(
        \registers[686][1] ), .D(\registers[687][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1666) );
  MX4X1 U7217 ( .A(\registers[332][2] ), .B(\registers[333][2] ), .C(
        \registers[334][2] ), .D(\registers[335][2] ), .S0(n4161), .S1(n4399), 
        .Y(n2139) );
  MX4X1 U7218 ( .A(\registers[380][2] ), .B(\registers[381][2] ), .C(
        \registers[382][2] ), .D(\registers[383][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2122) );
  MX4X1 U7219 ( .A(\registers[364][2] ), .B(\registers[365][2] ), .C(
        \registers[366][2] ), .D(\registers[367][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2127) );
  MX4X1 U7220 ( .A(\registers[76][2] ), .B(\registers[77][2] ), .C(
        \registers[78][2] ), .D(\registers[79][2] ), .S0(n4166), .S1(n4404), 
        .Y(n2226) );
  MX4X1 U7221 ( .A(\registers[124][2] ), .B(\registers[125][2] ), .C(
        \registers[126][2] ), .D(\registers[127][2] ), .S0(n4165), .S1(n4403), 
        .Y(n2211) );
  MX4X1 U7222 ( .A(\registers[108][2] ), .B(\registers[109][2] ), .C(
        \registers[110][2] ), .D(\registers[111][2] ), .S0(n4166), .S1(n4403), 
        .Y(n2216) );
  MX4X1 U7223 ( .A(\registers[12][2] ), .B(\registers[13][2] ), .C(
        \registers[14][2] ), .D(\registers[15][2] ), .S0(n4168), .S1(n4405), 
        .Y(n2248) );
  MX4X1 U7224 ( .A(\registers[60][2] ), .B(\registers[61][2] ), .C(
        \registers[62][2] ), .D(\registers[63][2] ), .S0(n4167), .S1(n4404), 
        .Y(n2232) );
  MX4X1 U7225 ( .A(\registers[44][2] ), .B(\registers[45][2] ), .C(
        \registers[46][2] ), .D(\registers[47][2] ), .S0(n4167), .S1(n4404), 
        .Y(n2238) );
  MX4X1 U7226 ( .A(\registers[204][2] ), .B(\registers[205][2] ), .C(
        \registers[206][2] ), .D(\registers[207][2] ), .S0(n4164), .S1(n4401), 
        .Y(n2183) );
  MX4X1 U7227 ( .A(\registers[252][2] ), .B(\registers[253][2] ), .C(
        \registers[254][2] ), .D(\registers[255][2] ), .S0(n4163), .S1(n4400), 
        .Y(n2167) );
  MX4X1 U7228 ( .A(\registers[236][2] ), .B(\registers[237][2] ), .C(
        \registers[238][2] ), .D(\registers[239][2] ), .S0(n4163), .S1(n4400), 
        .Y(n2173) );
  MX4X1 U7229 ( .A(\registers[140][2] ), .B(\registers[141][2] ), .C(
        \registers[142][2] ), .D(\registers[143][2] ), .S0(n4165), .S1(n4402), 
        .Y(n2205) );
  MX4X1 U7230 ( .A(\registers[188][2] ), .B(\registers[189][2] ), .C(
        \registers[190][2] ), .D(\registers[191][2] ), .S0(n4164), .S1(n4401), 
        .Y(n2189) );
  MX4X1 U7231 ( .A(\registers[172][2] ), .B(\registers[173][2] ), .C(
        \registers[174][2] ), .D(\registers[175][2] ), .S0(n4164), .S1(n4402), 
        .Y(n2194) );
  MX4X1 U7232 ( .A(\registers[844][2] ), .B(\registers[845][2] ), .C(
        \registers[846][2] ), .D(\registers[847][2] ), .S0(n4150), .S1(n4389), 
        .Y(n1962) );
  MX4X1 U7233 ( .A(\registers[892][2] ), .B(\registers[893][2] ), .C(
        \registers[894][2] ), .D(\registers[895][2] ), .S0(n4149), .S1(n4388), 
        .Y(n1947) );
  MX4X1 U7234 ( .A(\registers[876][2] ), .B(\registers[877][2] ), .C(
        \registers[878][2] ), .D(\registers[879][2] ), .S0(n4150), .S1(n4388), 
        .Y(n1952) );
  MX4X1 U7235 ( .A(\registers[780][2] ), .B(\registers[781][2] ), .C(
        \registers[782][2] ), .D(\registers[783][2] ), .S0(n4152), .S1(n4390), 
        .Y(n1984) );
  MX4X1 U7236 ( .A(\registers[828][2] ), .B(\registers[829][2] ), .C(
        \registers[830][2] ), .D(\registers[831][2] ), .S0(n4151), .S1(n4389), 
        .Y(n1968) );
  MX4X1 U7237 ( .A(\registers[812][2] ), .B(\registers[813][2] ), .C(
        \registers[814][2] ), .D(\registers[815][2] ), .S0(n4151), .S1(n4389), 
        .Y(n1974) );
  MX4X1 U7238 ( .A(\registers[972][2] ), .B(\registers[973][2] ), .C(
        \registers[974][2] ), .D(\registers[975][2] ), .S0(n4148), .S1(n4386), 
        .Y(n1919) );
  MX4X1 U7239 ( .A(\registers[1020][2] ), .B(\registers[1021][2] ), .C(
        \registers[1022][2] ), .D(\registers[1023][2] ), .S0(n4147), .S1(n4385), .Y(n1903) );
  MX4X1 U7240 ( .A(\registers[1004][2] ), .B(\registers[1005][2] ), .C(
        \registers[1006][2] ), .D(\registers[1007][2] ), .S0(n4147), .S1(n4386), .Y(n1909) );
  MX4X1 U7241 ( .A(\registers[908][2] ), .B(\registers[909][2] ), .C(
        \registers[910][2] ), .D(\registers[911][2] ), .S0(n4149), .S1(n4388), 
        .Y(n1941) );
  MX4X1 U7242 ( .A(\registers[956][2] ), .B(\registers[957][2] ), .C(
        \registers[958][2] ), .D(\registers[959][2] ), .S0(n4148), .S1(n4387), 
        .Y(n1925) );
  MX4X1 U7243 ( .A(\registers[940][2] ), .B(\registers[941][2] ), .C(
        \registers[942][2] ), .D(\registers[943][2] ), .S0(n4148), .S1(n4387), 
        .Y(n1930) );
  MX4X1 U7244 ( .A(\registers[588][2] ), .B(\registers[589][2] ), .C(
        \registers[590][2] ), .D(\registers[591][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2050) );
  MX4X1 U7245 ( .A(\registers[636][2] ), .B(\registers[637][2] ), .C(
        \registers[638][2] ), .D(\registers[639][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2034) );
  MX4X1 U7246 ( .A(\registers[620][2] ), .B(\registers[621][2] ), .C(
        \registers[622][2] ), .D(\registers[623][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2040) );
  MX4X1 U7247 ( .A(\registers[524][2] ), .B(\registers[525][2] ), .C(
        \registers[526][2] ), .D(\registers[527][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2072) );
  MX4X1 U7248 ( .A(\registers[572][2] ), .B(\registers[573][2] ), .C(
        \registers[574][2] ), .D(\registers[575][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2056) );
  MX4X1 U7249 ( .A(\registers[556][2] ), .B(\registers[557][2] ), .C(
        \registers[558][2] ), .D(\registers[559][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2061) );
  MX4X1 U7250 ( .A(\registers[716][2] ), .B(\registers[717][2] ), .C(
        \registers[718][2] ), .D(\registers[719][2] ), .S0(n4153), .S1(n4391), 
        .Y(n2007) );
  MX4X1 U7251 ( .A(\registers[764][2] ), .B(\registers[765][2] ), .C(
        \registers[766][2] ), .D(\registers[767][2] ), .S0(n4152), .S1(n4390), 
        .Y(n1991) );
  MX4X1 U7252 ( .A(\registers[748][2] ), .B(\registers[749][2] ), .C(
        \registers[750][2] ), .D(\registers[751][2] ), .S0(n4152), .S1(n4391), 
        .Y(n1996) );
  MX4X1 U7253 ( .A(\registers[652][2] ), .B(\registers[653][2] ), .C(
        \registers[654][2] ), .D(\registers[655][2] ), .S0(n4154), .S1(n4392), 
        .Y(n2028) );
  MX4X1 U7254 ( .A(\registers[700][2] ), .B(\registers[701][2] ), .C(
        \registers[702][2] ), .D(\registers[703][2] ), .S0(n4153), .S1(n4392), 
        .Y(n2013) );
  MX4X1 U7255 ( .A(\registers[684][2] ), .B(\registers[685][2] ), .C(
        \registers[686][2] ), .D(\registers[687][2] ), .S0(n4154), .S1(n4392), 
        .Y(n2018) );
  MX4X1 U7256 ( .A(\registers[332][3] ), .B(\registers[333][3] ), .C(
        \registers[334][3] ), .D(\registers[335][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2552) );
  MX4X1 U7257 ( .A(\registers[380][3] ), .B(\registers[381][3] ), .C(
        \registers[382][3] ), .D(\registers[383][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2537) );
  MX4X1 U7258 ( .A(\registers[364][3] ), .B(\registers[365][3] ), .C(
        \registers[366][3] ), .D(\registers[367][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2542) );
  MX4X1 U7259 ( .A(\registers[76][3] ), .B(\registers[77][3] ), .C(
        \registers[78][3] ), .D(\registers[79][3] ), .S0(n4188), .S1(n4423), 
        .Y(n2637) );
  MX4X1 U7260 ( .A(\registers[124][3] ), .B(\registers[125][3] ), .C(
        \registers[126][3] ), .D(\registers[127][3] ), .S0(n4187), .S1(n4422), 
        .Y(n2622) );
  MX4X1 U7261 ( .A(\registers[108][3] ), .B(\registers[109][3] ), .C(
        \registers[110][3] ), .D(\registers[111][3] ), .S0(n4187), .S1(n4423), 
        .Y(n2627) );
  MX4X1 U7262 ( .A(\registers[12][3] ), .B(\registers[13][3] ), .C(
        \registers[14][3] ), .D(\registers[15][3] ), .S0(n4189), .S1(n4424), 
        .Y(n2658) );
  MX4X1 U7263 ( .A(\registers[60][3] ), .B(\registers[61][3] ), .C(
        \registers[62][3] ), .D(\registers[63][3] ), .S0(n4188), .S1(n4424), 
        .Y(n2643) );
  MX4X1 U7264 ( .A(\registers[44][3] ), .B(\registers[45][3] ), .C(
        \registers[46][3] ), .D(\registers[47][3] ), .S0(n4188), .S1(n4424), 
        .Y(n2648) );
  MX4X1 U7265 ( .A(\registers[204][3] ), .B(\registers[205][3] ), .C(
        \registers[206][3] ), .D(\registers[207][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2595) );
  MX4X1 U7266 ( .A(\registers[252][3] ), .B(\registers[253][3] ), .C(
        \registers[254][3] ), .D(\registers[255][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2580) );
  MX4X1 U7267 ( .A(\registers[236][3] ), .B(\registers[237][3] ), .C(
        \registers[238][3] ), .D(\registers[239][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2585) );
  MX4X1 U7268 ( .A(\registers[140][3] ), .B(\registers[141][3] ), .C(
        \registers[142][3] ), .D(\registers[143][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2616) );
  MX4X1 U7269 ( .A(\registers[188][3] ), .B(\registers[189][3] ), .C(
        \registers[190][3] ), .D(\registers[191][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2601) );
  MX4X1 U7270 ( .A(\registers[172][3] ), .B(\registers[173][3] ), .C(
        \registers[174][3] ), .D(\registers[175][3] ), .S0(n4186), .S1(n4421), 
        .Y(n2606) );
  MX4X1 U7271 ( .A(\registers[844][3] ), .B(\registers[845][3] ), .C(
        \registers[846][3] ), .D(\registers[847][3] ), .S0(n4172), .S1(n4408), 
        .Y(n2314) );
  MX4X1 U7272 ( .A(\registers[892][3] ), .B(\registers[893][3] ), .C(
        \registers[894][3] ), .D(\registers[895][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2298) );
  MX4X1 U7273 ( .A(\registers[876][3] ), .B(\registers[877][3] ), .C(
        \registers[878][3] ), .D(\registers[879][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2304) );
  MX4X1 U7274 ( .A(\registers[780][3] ), .B(\registers[781][3] ), .C(
        \registers[782][3] ), .D(\registers[783][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2335) );
  MX4X1 U7275 ( .A(\registers[828][3] ), .B(\registers[829][3] ), .C(
        \registers[830][3] ), .D(\registers[831][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2320) );
  MX4X1 U7276 ( .A(\registers[812][3] ), .B(\registers[813][3] ), .C(
        \registers[814][3] ), .D(\registers[815][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2325) );
  MX4X1 U7277 ( .A(\registers[972][3] ), .B(\registers[973][3] ), .C(
        \registers[974][3] ), .D(\registers[975][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2271) );
  MX4X1 U7278 ( .A(\registers[1020][3] ), .B(\registers[1021][3] ), .C(
        \registers[1022][3] ), .D(\registers[1023][3] ), .S0(n4168), .S1(n4405), .Y(n2255) );
  MX4X1 U7279 ( .A(\registers[1004][3] ), .B(\registers[1005][3] ), .C(
        \registers[1006][3] ), .D(\registers[1007][3] ), .S0(n4168), .S1(n4405), .Y(n2260) );
  MX4X1 U7280 ( .A(\registers[908][3] ), .B(\registers[909][3] ), .C(
        \registers[910][3] ), .D(\registers[911][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2292) );
  MX4X1 U7281 ( .A(\registers[956][3] ), .B(\registers[957][3] ), .C(
        \registers[958][3] ), .D(\registers[959][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2277) );
  MX4X1 U7282 ( .A(\registers[940][3] ), .B(\registers[941][3] ), .C(
        \registers[942][3] ), .D(\registers[943][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2282) );
  MX4X1 U7283 ( .A(\registers[588][3] ), .B(\registers[589][3] ), .C(
        \registers[590][3] ), .D(\registers[591][3] ), .S0(n4177), .S1(n4413), 
        .Y(n2467) );
  MX4X1 U7284 ( .A(\registers[636][3] ), .B(\registers[637][3] ), .C(
        \registers[638][3] ), .D(\registers[639][3] ), .S0(n4176), .S1(n4412), 
        .Y(n2452) );
  MX4X1 U7285 ( .A(\registers[620][3] ), .B(\registers[621][3] ), .C(
        \registers[622][3] ), .D(\registers[623][3] ), .S0(n4176), .S1(n4413), 
        .Y(n2457) );
  MX4X1 U7286 ( .A(\registers[524][3] ), .B(\registers[525][3] ), .C(
        \registers[526][3] ), .D(\registers[527][3] ), .S0(n4178), .S1(n4415), 
        .Y(n2488) );
  MX4X1 U7287 ( .A(\registers[572][3] ), .B(\registers[573][3] ), .C(
        \registers[574][3] ), .D(\registers[575][3] ), .S0(n4177), .S1(n4414), 
        .Y(n2473) );
  MX4X1 U7288 ( .A(\registers[556][3] ), .B(\registers[557][3] ), .C(
        \registers[558][3] ), .D(\registers[559][3] ), .S0(n4178), .S1(n4414), 
        .Y(n2478) );
  MX4X1 U7289 ( .A(\registers[716][3] ), .B(\registers[717][3] ), .C(
        \registers[718][3] ), .D(\registers[719][3] ), .S0(n4174), .S1(n4411), 
        .Y(n2369) );
  MX4X1 U7290 ( .A(\registers[764][3] ), .B(\registers[765][3] ), .C(
        \registers[766][3] ), .D(\registers[767][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2351) );
  MX4X1 U7291 ( .A(\registers[748][3] ), .B(\registers[749][3] ), .C(
        \registers[750][3] ), .D(\registers[751][3] ), .S0(n4174), .S1(n4410), 
        .Y(n2358) );
  MX4X1 U7292 ( .A(\registers[652][3] ), .B(\registers[653][3] ), .C(
        \registers[654][3] ), .D(\registers[655][3] ), .S0(n4176), .S1(n4412), 
        .Y(n2446) );
  MX4X1 U7293 ( .A(\registers[700][3] ), .B(\registers[701][3] ), .C(
        \registers[702][3] ), .D(\registers[703][3] ), .S0(n4175), .S1(n4411), 
        .Y(n2376) );
  MX4X1 U7294 ( .A(\registers[684][3] ), .B(\registers[685][3] ), .C(
        \registers[686][3] ), .D(\registers[687][3] ), .S0(n4175), .S1(n4412), 
        .Y(n2382) );
  MX4X1 U7295 ( .A(\registers[332][4] ), .B(\registers[333][4] ), .C(
        \registers[334][4] ), .D(\registers[335][4] ), .S0(n4204), .S1(n4438), 
        .Y(n2892) );
  MX4X1 U7296 ( .A(\registers[380][4] ), .B(\registers[381][4] ), .C(
        \registers[382][4] ), .D(\registers[383][4] ), .S0(n4203), .S1(n4437), 
        .Y(n2877) );
  MX4X1 U7297 ( .A(\registers[364][4] ), .B(\registers[365][4] ), .C(
        \registers[366][4] ), .D(\registers[367][4] ), .S0(n4203), .S1(n4437), 
        .Y(n2882) );
  MX4X1 U7298 ( .A(\registers[76][4] ), .B(\registers[77][4] ), .C(
        \registers[78][4] ), .D(\registers[79][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2977) );
  MX4X1 U7299 ( .A(\registers[124][4] ), .B(\registers[125][4] ), .C(
        \registers[126][4] ), .D(\registers[127][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2962) );
  MX4X1 U7300 ( .A(\registers[108][4] ), .B(\registers[109][4] ), .C(
        \registers[110][4] ), .D(\registers[111][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2967) );
  MX4X1 U7301 ( .A(\registers[12][4] ), .B(\registers[13][4] ), .C(
        \registers[14][4] ), .D(\registers[15][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2998) );
  MX4X1 U7302 ( .A(\registers[60][4] ), .B(\registers[61][4] ), .C(
        \registers[62][4] ), .D(\registers[63][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2983) );
  MX4X1 U7303 ( .A(\registers[44][4] ), .B(\registers[45][4] ), .C(
        \registers[46][4] ), .D(\registers[47][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2988) );
  MX4X1 U7304 ( .A(\registers[204][4] ), .B(\registers[205][4] ), .C(
        \registers[206][4] ), .D(\registers[207][4] ), .S0(n4206), .S1(n4440), 
        .Y(n2935) );
  MX4X1 U7305 ( .A(\registers[252][4] ), .B(\registers[253][4] ), .C(
        \registers[254][4] ), .D(\registers[255][4] ), .S0(n4205), .S1(n4440), 
        .Y(n2920) );
  MX4X1 U7306 ( .A(\registers[236][4] ), .B(\registers[237][4] ), .C(
        \registers[238][4] ), .D(\registers[239][4] ), .S0(n4206), .S1(n4440), 
        .Y(n2925) );
  MX4X1 U7307 ( .A(\registers[140][4] ), .B(\registers[141][4] ), .C(
        \registers[142][4] ), .D(\registers[143][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2956) );
  MX4X1 U7308 ( .A(\registers[188][4] ), .B(\registers[189][4] ), .C(
        \registers[190][4] ), .D(\registers[191][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2941) );
  MX4X1 U7309 ( .A(\registers[172][4] ), .B(\registers[173][4] ), .C(
        \registers[174][4] ), .D(\registers[175][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2946) );
  MX4X1 U7310 ( .A(\registers[844][4] ), .B(\registers[845][4] ), .C(
        \registers[846][4] ), .D(\registers[847][4] ), .S0(n4193), .S1(n4428), 
        .Y(n2722) );
  MX4X1 U7311 ( .A(\registers[892][4] ), .B(\registers[893][4] ), .C(
        \registers[894][4] ), .D(\registers[895][4] ), .S0(n4192), .S1(n4427), 
        .Y(n2707) );
  MX4X1 U7312 ( .A(\registers[876][4] ), .B(\registers[877][4] ), .C(
        \registers[878][4] ), .D(\registers[879][4] ), .S0(n4192), .S1(n4428), 
        .Y(n2712) );
  MX4X1 U7313 ( .A(\registers[780][4] ), .B(\registers[781][4] ), .C(
        \registers[782][4] ), .D(\registers[783][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2743) );
  MX4X1 U7314 ( .A(\registers[828][4] ), .B(\registers[829][4] ), .C(
        \registers[830][4] ), .D(\registers[831][4] ), .S0(n4193), .S1(n4428), 
        .Y(n2728) );
  MX4X1 U7315 ( .A(\registers[812][4] ), .B(\registers[813][4] ), .C(
        \registers[814][4] ), .D(\registers[815][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2733) );
  MX4X1 U7316 ( .A(\registers[972][4] ), .B(\registers[973][4] ), .C(
        \registers[974][4] ), .D(\registers[975][4] ), .S0(n4190), .S1(n4426), 
        .Y(n2680) );
  MX4X1 U7317 ( .A(\registers[1020][4] ), .B(\registers[1021][4] ), .C(
        \registers[1022][4] ), .D(\registers[1023][4] ), .S0(n4189), .S1(n4425), .Y(n2665) );
  MX4X1 U7318 ( .A(\registers[1004][4] ), .B(\registers[1005][4] ), .C(
        \registers[1006][4] ), .D(\registers[1007][4] ), .S0(n4190), .S1(n4425), .Y(n2670) );
  MX4X1 U7319 ( .A(\registers[908][4] ), .B(\registers[909][4] ), .C(
        \registers[910][4] ), .D(\registers[911][4] ), .S0(n4192), .S1(n4427), 
        .Y(n2701) );
  MX4X1 U7320 ( .A(\registers[956][4] ), .B(\registers[957][4] ), .C(
        \registers[958][4] ), .D(\registers[959][4] ), .S0(n4191), .S1(n4426), 
        .Y(n2686) );
  MX4X1 U7321 ( .A(\registers[940][4] ), .B(\registers[941][4] ), .C(
        \registers[942][4] ), .D(\registers[943][4] ), .S0(n4191), .S1(n4426), 
        .Y(n2691) );
  MX4X1 U7322 ( .A(\registers[588][4] ), .B(\registers[589][4] ), .C(
        \registers[590][4] ), .D(\registers[591][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2807) );
  MX4X1 U7323 ( .A(\registers[636][4] ), .B(\registers[637][4] ), .C(
        \registers[638][4] ), .D(\registers[639][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2792) );
  MX4X1 U7324 ( .A(\registers[620][4] ), .B(\registers[621][4] ), .C(
        \registers[622][4] ), .D(\registers[623][4] ), .S0(n4198), .S1(n4432), 
        .Y(n2797) );
  MX4X1 U7325 ( .A(\registers[524][4] ), .B(\registers[525][4] ), .C(
        \registers[526][4] ), .D(\registers[527][4] ), .S0(n4200), .S1(n4434), 
        .Y(n2828) );
  MX4X1 U7326 ( .A(\registers[572][4] ), .B(\registers[573][4] ), .C(
        \registers[574][4] ), .D(\registers[575][4] ), .S0(n4199), .S1(n4433), 
        .Y(n2813) );
  MX4X1 U7327 ( .A(\registers[556][4] ), .B(\registers[557][4] ), .C(
        \registers[558][4] ), .D(\registers[559][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2818) );
  MX4X1 U7328 ( .A(\registers[716][4] ), .B(\registers[717][4] ), .C(
        \registers[718][4] ), .D(\registers[719][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2765) );
  MX4X1 U7329 ( .A(\registers[764][4] ), .B(\registers[765][4] ), .C(
        \registers[766][4] ), .D(\registers[767][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2750) );
  MX4X1 U7330 ( .A(\registers[748][4] ), .B(\registers[749][4] ), .C(
        \registers[750][4] ), .D(\registers[751][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2755) );
  MX4X1 U7331 ( .A(\registers[652][4] ), .B(\registers[653][4] ), .C(
        \registers[654][4] ), .D(\registers[655][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2786) );
  MX4X1 U7332 ( .A(\registers[700][4] ), .B(\registers[701][4] ), .C(
        \registers[702][4] ), .D(\registers[703][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2771) );
  MX4X1 U7333 ( .A(\registers[684][4] ), .B(\registers[685][4] ), .C(
        \registers[686][4] ), .D(\registers[687][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2776) );
  MX4X1 U7334 ( .A(\registers[332][5] ), .B(\registers[333][5] ), .C(
        \registers[334][5] ), .D(\registers[335][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3232) );
  MX4X1 U7335 ( .A(\registers[380][5] ), .B(\registers[381][5] ), .C(
        \registers[382][5] ), .D(\registers[383][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3217) );
  MX4X1 U7336 ( .A(\registers[364][5] ), .B(\registers[365][5] ), .C(
        \registers[366][5] ), .D(\registers[367][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3222) );
  MX4X1 U7337 ( .A(\registers[76][5] ), .B(\registers[77][5] ), .C(
        \registers[78][5] ), .D(\registers[79][5] ), .S0(n4230), .S1(n4463), 
        .Y(n3317) );
  MX4X1 U7338 ( .A(\registers[124][5] ), .B(\registers[125][5] ), .C(
        \registers[126][5] ), .D(\registers[127][5] ), .S0(n4229), .S1(n4462), 
        .Y(n3302) );
  MX4X1 U7339 ( .A(\registers[108][5] ), .B(\registers[109][5] ), .C(
        \registers[110][5] ), .D(\registers[111][5] ), .S0(n4230), .S1(n4462), 
        .Y(n3307) );
  MX4X1 U7340 ( .A(\registers[12][5] ), .B(\registers[13][5] ), .C(
        \registers[14][5] ), .D(\registers[15][5] ), .S0(n4232), .S1(n4464), 
        .Y(n3338) );
  MX4X1 U7341 ( .A(\registers[60][5] ), .B(\registers[61][5] ), .C(
        \registers[62][5] ), .D(\registers[63][5] ), .S0(n4231), .S1(n4463), 
        .Y(n3323) );
  MX4X1 U7342 ( .A(\registers[44][5] ), .B(\registers[45][5] ), .C(
        \registers[46][5] ), .D(\registers[47][5] ), .S0(n4231), .S1(n4463), 
        .Y(n3328) );
  MX4X1 U7343 ( .A(\registers[204][5] ), .B(\registers[205][5] ), .C(
        \registers[206][5] ), .D(\registers[207][5] ), .S0(n4228), .S1(n4460), 
        .Y(n3275) );
  MX4X1 U7344 ( .A(\registers[252][5] ), .B(\registers[253][5] ), .C(
        \registers[254][5] ), .D(\registers[255][5] ), .S0(n4227), .S1(n4459), 
        .Y(n3260) );
  MX4X1 U7345 ( .A(\registers[236][5] ), .B(\registers[237][5] ), .C(
        \registers[238][5] ), .D(\registers[239][5] ), .S0(n4227), .S1(n4460), 
        .Y(n3265) );
  MX4X1 U7346 ( .A(\registers[140][5] ), .B(\registers[141][5] ), .C(
        \registers[142][5] ), .D(\registers[143][5] ), .S0(n4229), .S1(n4461), 
        .Y(n3296) );
  MX4X1 U7347 ( .A(\registers[188][5] ), .B(\registers[189][5] ), .C(
        \registers[190][5] ), .D(\registers[191][5] ), .S0(n4228), .S1(n4460), 
        .Y(n3281) );
  MX4X1 U7348 ( .A(\registers[172][5] ), .B(\registers[173][5] ), .C(
        \registers[174][5] ), .D(\registers[175][5] ), .S0(n4228), .S1(n4461), 
        .Y(n3286) );
  MX4X1 U7349 ( .A(\registers[844][5] ), .B(\registers[845][5] ), .C(
        \registers[846][5] ), .D(\registers[847][5] ), .S0(n4214), .S1(n4448), 
        .Y(n3062) );
  MX4X1 U7350 ( .A(\registers[892][5] ), .B(\registers[893][5] ), .C(
        \registers[894][5] ), .D(\registers[895][5] ), .S0(n4213), .S1(n4447), 
        .Y(n3047) );
  MX4X1 U7351 ( .A(\registers[876][5] ), .B(\registers[877][5] ), .C(
        \registers[878][5] ), .D(\registers[879][5] ), .S0(n4214), .S1(n4447), 
        .Y(n3052) );
  MX4X1 U7352 ( .A(\registers[780][5] ), .B(\registers[781][5] ), .C(
        \registers[782][5] ), .D(\registers[783][5] ), .S0(n4216), .S1(n4449), 
        .Y(n3083) );
  MX4X1 U7353 ( .A(\registers[828][5] ), .B(\registers[829][5] ), .C(
        \registers[830][5] ), .D(\registers[831][5] ), .S0(n4215), .S1(n4448), 
        .Y(n3068) );
  MX4X1 U7354 ( .A(\registers[812][5] ), .B(\registers[813][5] ), .C(
        \registers[814][5] ), .D(\registers[815][5] ), .S0(n4215), .S1(n4448), 
        .Y(n3073) );
  MX4X1 U7355 ( .A(\registers[972][5] ), .B(\registers[973][5] ), .C(
        \registers[974][5] ), .D(\registers[975][5] ), .S0(n4212), .S1(n4445), 
        .Y(n3020) );
  MX4X1 U7356 ( .A(\registers[1020][5] ), .B(\registers[1021][5] ), .C(
        \registers[1022][5] ), .D(\registers[1023][5] ), .S0(n4211), .S1(n4444), .Y(n3005) );
  MX4X1 U7357 ( .A(\registers[1004][5] ), .B(\registers[1005][5] ), .C(
        \registers[1006][5] ), .D(\registers[1007][5] ), .S0(n4211), .S1(n4445), .Y(n3010) );
  MX4X1 U7358 ( .A(\registers[908][5] ), .B(\registers[909][5] ), .C(
        \registers[910][5] ), .D(\registers[911][5] ), .S0(n4213), .S1(n4447), 
        .Y(n3041) );
  MX4X1 U7359 ( .A(\registers[956][5] ), .B(\registers[957][5] ), .C(
        \registers[958][5] ), .D(\registers[959][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3026) );
  MX4X1 U7360 ( .A(\registers[940][5] ), .B(\registers[941][5] ), .C(
        \registers[942][5] ), .D(\registers[943][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3031) );
  MX4X1 U7361 ( .A(\registers[588][5] ), .B(\registers[589][5] ), .C(
        \registers[590][5] ), .D(\registers[591][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3147) );
  MX4X1 U7362 ( .A(\registers[636][5] ), .B(\registers[637][5] ), .C(
        \registers[638][5] ), .D(\registers[639][5] ), .S0(n4219), .S1(n4452), 
        .Y(n3132) );
  MX4X1 U7363 ( .A(\registers[620][5] ), .B(\registers[621][5] ), .C(
        \registers[622][5] ), .D(\registers[623][5] ), .S0(n4219), .S1(n4452), 
        .Y(n3137) );
  MX4X1 U7364 ( .A(\registers[524][5] ), .B(\registers[525][5] ), .C(
        \registers[526][5] ), .D(\registers[527][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3168) );
  MX4X1 U7365 ( .A(\registers[572][5] ), .B(\registers[573][5] ), .C(
        \registers[574][5] ), .D(\registers[575][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3153) );
  MX4X1 U7366 ( .A(\registers[556][5] ), .B(\registers[557][5] ), .C(
        \registers[558][5] ), .D(\registers[559][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3158) );
  MX4X1 U7367 ( .A(\registers[716][5] ), .B(\registers[717][5] ), .C(
        \registers[718][5] ), .D(\registers[719][5] ), .S0(n4217), .S1(n4450), 
        .Y(n3105) );
  MX4X1 U7368 ( .A(\registers[764][5] ), .B(\registers[765][5] ), .C(
        \registers[766][5] ), .D(\registers[767][5] ), .S0(n4216), .S1(n4449), 
        .Y(n3090) );
  MX4X1 U7369 ( .A(\registers[748][5] ), .B(\registers[749][5] ), .C(
        \registers[750][5] ), .D(\registers[751][5] ), .S0(n4216), .S1(n4450), 
        .Y(n3095) );
  MX4X1 U7370 ( .A(\registers[652][5] ), .B(\registers[653][5] ), .C(
        \registers[654][5] ), .D(\registers[655][5] ), .S0(n4218), .S1(n4452), 
        .Y(n3126) );
  MX4X1 U7371 ( .A(\registers[700][5] ), .B(\registers[701][5] ), .C(
        \registers[702][5] ), .D(\registers[703][5] ), .S0(n4217), .S1(n4451), 
        .Y(n3111) );
  MX4X1 U7372 ( .A(\registers[684][5] ), .B(\registers[685][5] ), .C(
        \registers[686][5] ), .D(\registers[687][5] ), .S0(n4218), .S1(n4451), 
        .Y(n3116) );
  MX4X1 U7373 ( .A(\registers[332][6] ), .B(\registers[333][6] ), .C(
        \registers[334][6] ), .D(\registers[335][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3572) );
  MX4X1 U7374 ( .A(\registers[380][6] ), .B(\registers[381][6] ), .C(
        \registers[382][6] ), .D(\registers[383][6] ), .S0(n4245), .S1(n4476), 
        .Y(n3557) );
  MX4X1 U7375 ( .A(\registers[364][6] ), .B(\registers[365][6] ), .C(
        \registers[366][6] ), .D(\registers[367][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3562) );
  MX4X1 U7376 ( .A(\registers[76][6] ), .B(\registers[77][6] ), .C(
        \registers[78][6] ), .D(\registers[79][6] ), .S0(n4252), .S1(n4482), 
        .Y(n3657) );
  MX4X1 U7377 ( .A(\registers[124][6] ), .B(\registers[125][6] ), .C(
        \registers[126][6] ), .D(\registers[127][6] ), .S0(n4251), .S1(n4481), 
        .Y(n3642) );
  MX4X1 U7378 ( .A(\registers[108][6] ), .B(\registers[109][6] ), .C(
        \registers[110][6] ), .D(\registers[111][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3647) );
  MX4X1 U7379 ( .A(\registers[12][6] ), .B(\registers[13][6] ), .C(
        \registers[14][6] ), .D(\registers[15][6] ), .S0(n4253), .S1(n4484), 
        .Y(n3678) );
  MX4X1 U7380 ( .A(\registers[60][6] ), .B(\registers[61][6] ), .C(
        \registers[62][6] ), .D(\registers[63][6] ), .S0(n4252), .S1(n4483), 
        .Y(n3663) );
  MX4X1 U7381 ( .A(\registers[44][6] ), .B(\registers[45][6] ), .C(
        \registers[46][6] ), .D(\registers[47][6] ), .S0(n4252), .S1(n4483), 
        .Y(n3668) );
  MX4X1 U7382 ( .A(\registers[204][6] ), .B(\registers[205][6] ), .C(
        \registers[206][6] ), .D(\registers[207][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3615) );
  MX4X1 U7383 ( .A(\registers[252][6] ), .B(\registers[253][6] ), .C(
        \registers[254][6] ), .D(\registers[255][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3600) );
  MX4X1 U7384 ( .A(\registers[236][6] ), .B(\registers[237][6] ), .C(
        \registers[238][6] ), .D(\registers[239][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3605) );
  MX4X1 U7385 ( .A(\registers[140][6] ), .B(\registers[141][6] ), .C(
        \registers[142][6] ), .D(\registers[143][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3636) );
  MX4X1 U7386 ( .A(\registers[188][6] ), .B(\registers[189][6] ), .C(
        \registers[190][6] ), .D(\registers[191][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3621) );
  MX4X1 U7387 ( .A(\registers[172][6] ), .B(\registers[173][6] ), .C(
        \registers[174][6] ), .D(\registers[175][6] ), .S0(n4250), .S1(n4480), 
        .Y(n3626) );
  MX4X1 U7388 ( .A(\registers[844][6] ), .B(\registers[845][6] ), .C(
        \registers[846][6] ), .D(\registers[847][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3402) );
  MX4X1 U7389 ( .A(\registers[892][6] ), .B(\registers[893][6] ), .C(
        \registers[894][6] ), .D(\registers[895][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3387) );
  MX4X1 U7390 ( .A(\registers[876][6] ), .B(\registers[877][6] ), .C(
        \registers[878][6] ), .D(\registers[879][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3392) );
  MX4X1 U7391 ( .A(\registers[780][6] ), .B(\registers[781][6] ), .C(
        \registers[782][6] ), .D(\registers[783][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3423) );
  MX4X1 U7392 ( .A(\registers[828][6] ), .B(\registers[829][6] ), .C(
        \registers[830][6] ), .D(\registers[831][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3408) );
  MX4X1 U7393 ( .A(\registers[812][6] ), .B(\registers[813][6] ), .C(
        \registers[814][6] ), .D(\registers[815][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3413) );
  MX4X1 U7394 ( .A(\registers[972][6] ), .B(\registers[973][6] ), .C(
        \registers[974][6] ), .D(\registers[975][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3360) );
  MX4X1 U7395 ( .A(\registers[1020][6] ), .B(\registers[1021][6] ), .C(
        \registers[1022][6] ), .D(\registers[1023][6] ), .S0(n4232), .S1(n4464), .Y(n3345) );
  MX4X1 U7396 ( .A(\registers[1004][6] ), .B(\registers[1005][6] ), .C(
        \registers[1006][6] ), .D(\registers[1007][6] ), .S0(n4232), .S1(n4464), .Y(n3350) );
  MX4X1 U7397 ( .A(\registers[908][6] ), .B(\registers[909][6] ), .C(
        \registers[910][6] ), .D(\registers[911][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3381) );
  MX4X1 U7398 ( .A(\registers[956][6] ), .B(\registers[957][6] ), .C(
        \registers[958][6] ), .D(\registers[959][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3366) );
  MX4X1 U7399 ( .A(\registers[940][6] ), .B(\registers[941][6] ), .C(
        \registers[942][6] ), .D(\registers[943][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3371) );
  MX4X1 U7400 ( .A(\registers[588][6] ), .B(\registers[589][6] ), .C(
        \registers[590][6] ), .D(\registers[591][6] ), .S0(n4241), .S1(n4472), 
        .Y(n3487) );
  MX4X1 U7401 ( .A(\registers[636][6] ), .B(\registers[637][6] ), .C(
        \registers[638][6] ), .D(\registers[639][6] ), .S0(n4240), .S1(n4472), 
        .Y(n3472) );
  MX4X1 U7402 ( .A(\registers[620][6] ), .B(\registers[621][6] ), .C(
        \registers[622][6] ), .D(\registers[623][6] ), .S0(n4240), .S1(n4472), 
        .Y(n3477) );
  MX4X1 U7403 ( .A(\registers[524][6] ), .B(\registers[525][6] ), .C(
        \registers[526][6] ), .D(\registers[527][6] ), .S0(n4242), .S1(n4474), 
        .Y(n3508) );
  MX4X1 U7404 ( .A(\registers[572][6] ), .B(\registers[573][6] ), .C(
        \registers[574][6] ), .D(\registers[575][6] ), .S0(n4241), .S1(n4473), 
        .Y(n3493) );
  MX4X1 U7405 ( .A(\registers[556][6] ), .B(\registers[557][6] ), .C(
        \registers[558][6] ), .D(\registers[559][6] ), .S0(n4242), .S1(n4473), 
        .Y(n3498) );
  MX4X1 U7406 ( .A(\registers[716][6] ), .B(\registers[717][6] ), .C(
        \registers[718][6] ), .D(\registers[719][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3445) );
  MX4X1 U7407 ( .A(\registers[764][6] ), .B(\registers[765][6] ), .C(
        \registers[766][6] ), .D(\registers[767][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3430) );
  MX4X1 U7408 ( .A(\registers[748][6] ), .B(\registers[749][6] ), .C(
        \registers[750][6] ), .D(\registers[751][6] ), .S0(n4238), .S1(n4469), 
        .Y(n3435) );
  MX4X1 U7409 ( .A(\registers[652][6] ), .B(\registers[653][6] ), .C(
        \registers[654][6] ), .D(\registers[655][6] ), .S0(n4240), .S1(n4471), 
        .Y(n3466) );
  MX4X1 U7410 ( .A(\registers[700][6] ), .B(\registers[701][6] ), .C(
        \registers[702][6] ), .D(\registers[703][6] ), .S0(n4239), .S1(n4470), 
        .Y(n3451) );
  MX4X1 U7411 ( .A(\registers[684][6] ), .B(\registers[685][6] ), .C(
        \registers[686][6] ), .D(\registers[687][6] ), .S0(n4239), .S1(n4471), 
        .Y(n3456) );
  MX4X1 U7412 ( .A(\registers[332][7] ), .B(\registers[333][7] ), .C(
        \registers[334][7] ), .D(\registers[335][7] ), .S0(n4268), .S1(n4480), 
        .Y(n3912) );
  MX4X1 U7413 ( .A(\registers[380][7] ), .B(\registers[381][7] ), .C(
        \registers[382][7] ), .D(\registers[383][7] ), .S0(n4267), .S1(n4496), 
        .Y(n3897) );
  MX4X1 U7414 ( .A(\registers[364][7] ), .B(\registers[365][7] ), .C(
        \registers[366][7] ), .D(\registers[367][7] ), .S0(n4267), .S1(n4496), 
        .Y(n3902) );
  MX4X1 U7415 ( .A(\registers[76][7] ), .B(\registers[77][7] ), .C(
        \registers[78][7] ), .D(\registers[79][7] ), .S0(n4273), .S1(n4451), 
        .Y(n3997) );
  MX4X1 U7416 ( .A(\registers[124][7] ), .B(\registers[125][7] ), .C(
        \registers[126][7] ), .D(\registers[127][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3982) );
  MX4X1 U7417 ( .A(\registers[108][7] ), .B(\registers[109][7] ), .C(
        \registers[110][7] ), .D(\registers[111][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3987) );
  MX4X1 U7418 ( .A(\registers[12][7] ), .B(\registers[13][7] ), .C(
        \registers[14][7] ), .D(\registers[15][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4018) );
  MX4X1 U7419 ( .A(\registers[60][7] ), .B(\registers[61][7] ), .C(
        \registers[62][7] ), .D(\registers[63][7] ), .S0(n4273), .S1(n4453), 
        .Y(n4003) );
  MX4X1 U7420 ( .A(\registers[44][7] ), .B(\registers[45][7] ), .C(
        \registers[46][7] ), .D(\registers[47][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4008) );
  MX4X1 U7421 ( .A(\registers[204][7] ), .B(\registers[205][7] ), .C(
        \registers[206][7] ), .D(\registers[207][7] ), .S0(n4270), .S1(n4499), 
        .Y(n3955) );
  MX4X1 U7422 ( .A(\registers[252][7] ), .B(\registers[253][7] ), .C(
        \registers[254][7] ), .D(\registers[255][7] ), .S0(n4269), .S1(n4498), 
        .Y(n3940) );
  MX4X1 U7423 ( .A(\registers[236][7] ), .B(\registers[237][7] ), .C(
        \registers[238][7] ), .D(\registers[239][7] ), .S0(n4270), .S1(n4498), 
        .Y(n3945) );
  MX4X1 U7424 ( .A(\registers[140][7] ), .B(\registers[141][7] ), .C(
        \registers[142][7] ), .D(\registers[143][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3976) );
  MX4X1 U7425 ( .A(\registers[188][7] ), .B(\registers[189][7] ), .C(
        \registers[190][7] ), .D(\registers[191][7] ), .S0(n4271), .S1(n4499), 
        .Y(n3961) );
  MX4X1 U7426 ( .A(\registers[172][7] ), .B(\registers[173][7] ), .C(
        \registers[174][7] ), .D(\registers[175][7] ), .S0(n4271), .S1(n4499), 
        .Y(n3966) );
  MX4X1 U7427 ( .A(\registers[844][7] ), .B(\registers[845][7] ), .C(
        \registers[846][7] ), .D(\registers[847][7] ), .S0(n4257), .S1(n4487), 
        .Y(n3742) );
  MX4X1 U7428 ( .A(\registers[892][7] ), .B(\registers[893][7] ), .C(
        \registers[894][7] ), .D(\registers[895][7] ), .S0(n4256), .S1(n4486), 
        .Y(n3727) );
  MX4X1 U7429 ( .A(\registers[876][7] ), .B(\registers[877][7] ), .C(
        \registers[878][7] ), .D(\registers[879][7] ), .S0(n4256), .S1(n4487), 
        .Y(n3732) );
  MX4X1 U7430 ( .A(\registers[780][7] ), .B(\registers[781][7] ), .C(
        \registers[782][7] ), .D(\registers[783][7] ), .S0(n4258), .S1(n4488), 
        .Y(n3763) );
  MX4X1 U7431 ( .A(\registers[828][7] ), .B(\registers[829][7] ), .C(
        \registers[830][7] ), .D(\registers[831][7] ), .S0(n4257), .S1(n4488), 
        .Y(n3748) );
  MX4X1 U7432 ( .A(\registers[812][7] ), .B(\registers[813][7] ), .C(
        \registers[814][7] ), .D(\registers[815][7] ), .S0(n4258), .S1(n4488), 
        .Y(n3753) );
  MX4X1 U7433 ( .A(\registers[972][7] ), .B(\registers[973][7] ), .C(
        \registers[974][7] ), .D(\registers[975][7] ), .S0(n4254), .S1(n4485), 
        .Y(n3700) );
  MX4X1 U7434 ( .A(\registers[1020][7] ), .B(\registers[1021][7] ), .C(
        \registers[1022][7] ), .D(\registers[1023][7] ), .S0(n4253), .S1(n4484), .Y(n3685) );
  MX4X1 U7435 ( .A(\registers[1004][7] ), .B(\registers[1005][7] ), .C(
        \registers[1006][7] ), .D(\registers[1007][7] ), .S0(n4254), .S1(n4484), .Y(n3690) );
  MX4X1 U7436 ( .A(\registers[908][7] ), .B(\registers[909][7] ), .C(
        \registers[910][7] ), .D(\registers[911][7] ), .S0(n4256), .S1(n4486), 
        .Y(n3721) );
  MX4X1 U7437 ( .A(\registers[956][7] ), .B(\registers[957][7] ), .C(
        \registers[958][7] ), .D(\registers[959][7] ), .S0(n4255), .S1(n4485), 
        .Y(n3706) );
  MX4X1 U7438 ( .A(\registers[940][7] ), .B(\registers[941][7] ), .C(
        \registers[942][7] ), .D(\registers[943][7] ), .S0(n4255), .S1(n4485), 
        .Y(n3711) );
  MX4X1 U7439 ( .A(\registers[588][7] ), .B(\registers[589][7] ), .C(
        \registers[590][7] ), .D(\registers[591][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3827) );
  MX4X1 U7440 ( .A(\registers[636][7] ), .B(\registers[637][7] ), .C(
        \registers[638][7] ), .D(\registers[639][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3812) );
  MX4X1 U7441 ( .A(\registers[620][7] ), .B(\registers[621][7] ), .C(
        \registers[622][7] ), .D(\registers[623][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3817) );
  MX4X1 U7442 ( .A(\registers[524][7] ), .B(\registers[525][7] ), .C(
        \registers[526][7] ), .D(\registers[527][7] ), .S0(n4264), .S1(n4493), 
        .Y(n3848) );
  MX4X1 U7443 ( .A(\registers[572][7] ), .B(\registers[573][7] ), .C(
        \registers[574][7] ), .D(\registers[575][7] ), .S0(n4263), .S1(n4492), 
        .Y(n3833) );
  MX4X1 U7444 ( .A(\registers[556][7] ), .B(\registers[557][7] ), .C(
        \registers[558][7] ), .D(\registers[559][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3838) );
  MX4X1 U7445 ( .A(\registers[716][7] ), .B(\registers[717][7] ), .C(
        \registers[718][7] ), .D(\registers[719][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3785) );
  MX4X1 U7446 ( .A(\registers[764][7] ), .B(\registers[765][7] ), .C(
        \registers[766][7] ), .D(\registers[767][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3770) );
  MX4X1 U7447 ( .A(\registers[748][7] ), .B(\registers[749][7] ), .C(
        \registers[750][7] ), .D(\registers[751][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3775) );
  MX4X1 U7448 ( .A(\registers[652][7] ), .B(\registers[653][7] ), .C(
        \registers[654][7] ), .D(\registers[655][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3806) );
  MX4X1 U7449 ( .A(\registers[700][7] ), .B(\registers[701][7] ), .C(
        \registers[702][7] ), .D(\registers[703][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3791) );
  MX4X1 U7450 ( .A(\registers[684][7] ), .B(\registers[685][7] ), .C(
        \registers[686][7] ), .D(\registers[687][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3796) );
  MX4X1 U7451 ( .A(\registers[332][0] ), .B(\registers[333][0] ), .C(
        \registers[334][0] ), .D(\registers[335][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4877) );
  MX4X1 U7452 ( .A(\registers[380][0] ), .B(\registers[381][0] ), .C(
        \registers[382][0] ), .D(\registers[383][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4862) );
  MX4X1 U7453 ( .A(\registers[364][0] ), .B(\registers[365][0] ), .C(
        \registers[366][0] ), .D(\registers[367][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4867) );
  MX4X1 U7454 ( .A(\registers[76][0] ), .B(\registers[77][0] ), .C(
        \registers[78][0] ), .D(\registers[79][0] ), .S0(n7467), .S1(n7708), 
        .Y(n4962) );
  MX4X1 U7455 ( .A(\registers[124][0] ), .B(\registers[125][0] ), .C(
        \registers[126][0] ), .D(\registers[127][0] ), .S0(n7466), .S1(n7707), 
        .Y(n4947) );
  MX4X1 U7456 ( .A(\registers[108][0] ), .B(\registers[109][0] ), .C(
        \registers[110][0] ), .D(\registers[111][0] ), .S0(n7466), .S1(n7708), 
        .Y(n4952) );
  MX4X1 U7457 ( .A(\registers[12][0] ), .B(\registers[13][0] ), .C(
        \registers[14][0] ), .D(\registers[15][0] ), .S0(n7468), .S1(n7709), 
        .Y(n4983) );
  MX4X1 U7458 ( .A(\registers[60][0] ), .B(\registers[61][0] ), .C(
        \registers[62][0] ), .D(\registers[63][0] ), .S0(n7467), .S1(n7708), 
        .Y(n4968) );
  MX4X1 U7459 ( .A(\registers[44][0] ), .B(\registers[45][0] ), .C(
        \registers[46][0] ), .D(\registers[47][0] ), .S0(n7467), .S1(n7709), 
        .Y(n4973) );
  MX4X1 U7460 ( .A(\registers[204][0] ), .B(\registers[205][0] ), .C(
        \registers[206][0] ), .D(\registers[207][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4920) );
  MX4X1 U7461 ( .A(\registers[252][0] ), .B(\registers[253][0] ), .C(
        \registers[254][0] ), .D(\registers[255][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4905) );
  MX4X1 U7462 ( .A(\registers[236][0] ), .B(\registers[237][0] ), .C(
        \registers[238][0] ), .D(\registers[239][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4910) );
  MX4X1 U7463 ( .A(\registers[140][0] ), .B(\registers[141][0] ), .C(
        \registers[142][0] ), .D(\registers[143][0] ), .S0(n7465), .S1(n7707), 
        .Y(n4941) );
  MX4X1 U7464 ( .A(\registers[188][0] ), .B(\registers[189][0] ), .C(
        \registers[190][0] ), .D(\registers[191][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4926) );
  MX4X1 U7465 ( .A(\registers[172][0] ), .B(\registers[173][0] ), .C(
        \registers[174][0] ), .D(\registers[175][0] ), .S0(n7465), .S1(n7706), 
        .Y(n4931) );
  MX4X1 U7466 ( .A(\registers[844][0] ), .B(\registers[845][0] ), .C(
        \registers[846][0] ), .D(\registers[847][0] ), .S0(n7451), .S1(n7693), 
        .Y(n4707) );
  MX4X1 U7467 ( .A(\registers[892][0] ), .B(\registers[893][0] ), .C(
        \registers[894][0] ), .D(\registers[895][0] ), .S0(n7450), .S1(n7692), 
        .Y(n4692) );
  MX4X1 U7468 ( .A(\registers[876][0] ), .B(\registers[877][0] ), .C(
        \registers[878][0] ), .D(\registers[879][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4697) );
  MX4X1 U7469 ( .A(\registers[780][0] ), .B(\registers[781][0] ), .C(
        \registers[782][0] ), .D(\registers[783][0] ), .S0(n7452), .S1(n7695), 
        .Y(n4728) );
  MX4X1 U7470 ( .A(\registers[828][0] ), .B(\registers[829][0] ), .C(
        \registers[830][0] ), .D(\registers[831][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4713) );
  MX4X1 U7471 ( .A(\registers[812][0] ), .B(\registers[813][0] ), .C(
        \registers[814][0] ), .D(\registers[815][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4718) );
  MX4X1 U7472 ( .A(\registers[972][0] ), .B(\registers[973][0] ), .C(
        \registers[974][0] ), .D(\registers[975][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4665) );
  MX4X1 U7473 ( .A(\registers[908][0] ), .B(\registers[909][0] ), .C(
        \registers[910][0] ), .D(\registers[911][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4686) );
  MX4X1 U7474 ( .A(\registers[956][0] ), .B(\registers[957][0] ), .C(
        \registers[958][0] ), .D(\registers[959][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4671) );
  MX4X1 U7475 ( .A(\registers[940][0] ), .B(\registers[941][0] ), .C(
        \registers[942][0] ), .D(\registers[943][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4676) );
  MX4X1 U7476 ( .A(\registers[588][0] ), .B(\registers[589][0] ), .C(
        \registers[590][0] ), .D(\registers[591][0] ), .S0(n7456), .S1(n7698), 
        .Y(n4792) );
  MX4X1 U7477 ( .A(\registers[636][0] ), .B(\registers[637][0] ), .C(
        \registers[638][0] ), .D(\registers[639][0] ), .S0(n7455), .S1(n7697), 
        .Y(n4777) );
  MX4X1 U7478 ( .A(\registers[620][0] ), .B(\registers[621][0] ), .C(
        \registers[622][0] ), .D(\registers[623][0] ), .S0(n7455), .S1(n7698), 
        .Y(n4782) );
  MX4X1 U7479 ( .A(\registers[524][0] ), .B(\registers[525][0] ), .C(
        \registers[526][0] ), .D(\registers[527][0] ), .S0(n7457), .S1(n7700), 
        .Y(n4813) );
  MX4X1 U7480 ( .A(\registers[572][0] ), .B(\registers[573][0] ), .C(
        \registers[574][0] ), .D(\registers[575][0] ), .S0(n7456), .S1(n7699), 
        .Y(n4798) );
  MX4X1 U7481 ( .A(\registers[556][0] ), .B(\registers[557][0] ), .C(
        \registers[558][0] ), .D(\registers[559][0] ), .S0(n7457), .S1(n7699), 
        .Y(n4803) );
  MX4X1 U7482 ( .A(\registers[716][0] ), .B(\registers[717][0] ), .C(
        \registers[718][0] ), .D(\registers[719][0] ), .S0(n7453), .S1(n7696), 
        .Y(n4750) );
  MX4X1 U7483 ( .A(\registers[764][0] ), .B(\registers[765][0] ), .C(
        \registers[766][0] ), .D(\registers[767][0] ), .S0(n7452), .S1(n7695), 
        .Y(n4735) );
  MX4X1 U7484 ( .A(\registers[748][0] ), .B(\registers[749][0] ), .C(
        \registers[750][0] ), .D(\registers[751][0] ), .S0(n7453), .S1(n7695), 
        .Y(n4740) );
  MX4X1 U7485 ( .A(\registers[652][0] ), .B(\registers[653][0] ), .C(
        \registers[654][0] ), .D(\registers[655][0] ), .S0(n7455), .S1(n7697), 
        .Y(n4771) );
  MX4X1 U7486 ( .A(\registers[700][0] ), .B(\registers[701][0] ), .C(
        \registers[702][0] ), .D(\registers[703][0] ), .S0(n7454), .S1(n7696), 
        .Y(n4756) );
  MX4X1 U7487 ( .A(\registers[684][0] ), .B(\registers[685][0] ), .C(
        \registers[686][0] ), .D(\registers[687][0] ), .S0(n7454), .S1(n7696), 
        .Y(n4761) );
  MX4X1 U7488 ( .A(\registers[332][1] ), .B(\registers[333][1] ), .C(
        \registers[334][1] ), .D(\registers[335][1] ), .S0(n7483), .S1(n7723), 
        .Y(n5217) );
  MX4X1 U7489 ( .A(\registers[380][1] ), .B(\registers[381][1] ), .C(
        \registers[382][1] ), .D(\registers[383][1] ), .S0(n7482), .S1(n7722), 
        .Y(n5202) );
  MX4X1 U7490 ( .A(\registers[364][1] ), .B(\registers[365][1] ), .C(
        \registers[366][1] ), .D(\registers[367][1] ), .S0(n7482), .S1(n7722), 
        .Y(n5207) );
  MX4X1 U7491 ( .A(\registers[76][1] ), .B(\registers[77][1] ), .C(
        \registers[78][1] ), .D(\registers[79][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5302) );
  MX4X1 U7492 ( .A(\registers[124][1] ), .B(\registers[125][1] ), .C(
        \registers[126][1] ), .D(\registers[127][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5287) );
  MX4X1 U7493 ( .A(\registers[108][1] ), .B(\registers[109][1] ), .C(
        \registers[110][1] ), .D(\registers[111][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5292) );
  MX4X1 U7494 ( .A(\registers[12][1] ), .B(\registers[13][1] ), .C(
        \registers[14][1] ), .D(\registers[15][1] ), .S0(n7489), .S1(n7729), 
        .Y(n5323) );
  MX4X1 U7495 ( .A(\registers[60][1] ), .B(\registers[61][1] ), .C(
        \registers[62][1] ), .D(\registers[63][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5308) );
  MX4X1 U7496 ( .A(\registers[44][1] ), .B(\registers[45][1] ), .C(
        \registers[46][1] ), .D(\registers[47][1] ), .S0(n7489), .S1(n7728), 
        .Y(n5313) );
  MX4X1 U7497 ( .A(\registers[204][1] ), .B(\registers[205][1] ), .C(
        \registers[206][1] ), .D(\registers[207][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5260) );
  MX4X1 U7498 ( .A(\registers[252][1] ), .B(\registers[253][1] ), .C(
        \registers[254][1] ), .D(\registers[255][1] ), .S0(n7484), .S1(n7724), 
        .Y(n5245) );
  MX4X1 U7499 ( .A(\registers[236][1] ), .B(\registers[237][1] ), .C(
        \registers[238][1] ), .D(\registers[239][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5250) );
  MX4X1 U7500 ( .A(\registers[140][1] ), .B(\registers[141][1] ), .C(
        \registers[142][1] ), .D(\registers[143][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5281) );
  MX4X1 U7501 ( .A(\registers[188][1] ), .B(\registers[189][1] ), .C(
        \registers[190][1] ), .D(\registers[191][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5266) );
  MX4X1 U7502 ( .A(\registers[172][1] ), .B(\registers[173][1] ), .C(
        \registers[174][1] ), .D(\registers[175][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5271) );
  MX4X1 U7503 ( .A(\registers[844][1] ), .B(\registers[845][1] ), .C(
        \registers[846][1] ), .D(\registers[847][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5047) );
  MX4X1 U7504 ( .A(\registers[892][1] ), .B(\registers[893][1] ), .C(
        \registers[894][1] ), .D(\registers[895][1] ), .S0(n7471), .S1(n7712), 
        .Y(n5032) );
  MX4X1 U7505 ( .A(\registers[876][1] ), .B(\registers[877][1] ), .C(
        \registers[878][1] ), .D(\registers[879][1] ), .S0(n7471), .S1(n7712), 
        .Y(n5037) );
  MX4X1 U7506 ( .A(\registers[780][1] ), .B(\registers[781][1] ), .C(
        \registers[782][1] ), .D(\registers[783][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5068) );
  MX4X1 U7507 ( .A(\registers[828][1] ), .B(\registers[829][1] ), .C(
        \registers[830][1] ), .D(\registers[831][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5053) );
  MX4X1 U7508 ( .A(\registers[812][1] ), .B(\registers[813][1] ), .C(
        \registers[814][1] ), .D(\registers[815][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5058) );
  MX4X1 U7509 ( .A(\registers[972][1] ), .B(\registers[973][1] ), .C(
        \registers[974][1] ), .D(\registers[975][1] ), .S0(n7469), .S1(n7711), 
        .Y(n5005) );
  MX4X1 U7510 ( .A(\registers[1020][1] ), .B(\registers[1021][1] ), .C(
        \registers[1022][1] ), .D(\registers[1023][1] ), .S0(n7468), .S1(n7710), .Y(n4990) );
  MX4X1 U7511 ( .A(\registers[1004][1] ), .B(\registers[1005][1] ), .C(
        \registers[1006][1] ), .D(\registers[1007][1] ), .S0(n7469), .S1(n7710), .Y(n4995) );
  MX4X1 U7512 ( .A(\registers[908][1] ), .B(\registers[909][1] ), .C(
        \registers[910][1] ), .D(\registers[911][1] ), .S0(n7471), .S1(n7712), 
        .Y(n5026) );
  MX4X1 U7513 ( .A(\registers[956][1] ), .B(\registers[957][1] ), .C(
        \registers[958][1] ), .D(\registers[959][1] ), .S0(n7470), .S1(n7711), 
        .Y(n5011) );
  MX4X1 U7514 ( .A(\registers[940][1] ), .B(\registers[941][1] ), .C(
        \registers[942][1] ), .D(\registers[943][1] ), .S0(n7470), .S1(n7711), 
        .Y(n5016) );
  MX4X1 U7515 ( .A(\registers[588][1] ), .B(\registers[589][1] ), .C(
        \registers[590][1] ), .D(\registers[591][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5132) );
  MX4X1 U7516 ( .A(\registers[636][1] ), .B(\registers[637][1] ), .C(
        \registers[638][1] ), .D(\registers[639][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5117) );
  MX4X1 U7517 ( .A(\registers[620][1] ), .B(\registers[621][1] ), .C(
        \registers[622][1] ), .D(\registers[623][1] ), .S0(n7477), .S1(n7717), 
        .Y(n5122) );
  MX4X1 U7518 ( .A(\registers[524][1] ), .B(\registers[525][1] ), .C(
        \registers[526][1] ), .D(\registers[527][1] ), .S0(n7479), .S1(n7719), 
        .Y(n5153) );
  MX4X1 U7519 ( .A(\registers[572][1] ), .B(\registers[573][1] ), .C(
        \registers[574][1] ), .D(\registers[575][1] ), .S0(n7478), .S1(n7718), 
        .Y(n5138) );
  MX4X1 U7520 ( .A(\registers[556][1] ), .B(\registers[557][1] ), .C(
        \registers[558][1] ), .D(\registers[559][1] ), .S0(n7478), .S1(n7719), 
        .Y(n5143) );
  MX4X1 U7521 ( .A(\registers[716][1] ), .B(\registers[717][1] ), .C(
        \registers[718][1] ), .D(\registers[719][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5090) );
  MX4X1 U7522 ( .A(\registers[764][1] ), .B(\registers[765][1] ), .C(
        \registers[766][1] ), .D(\registers[767][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5075) );
  MX4X1 U7523 ( .A(\registers[748][1] ), .B(\registers[749][1] ), .C(
        \registers[750][1] ), .D(\registers[751][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5080) );
  MX4X1 U7524 ( .A(\registers[652][1] ), .B(\registers[653][1] ), .C(
        \registers[654][1] ), .D(\registers[655][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5111) );
  MX4X1 U7525 ( .A(\registers[700][1] ), .B(\registers[701][1] ), .C(
        \registers[702][1] ), .D(\registers[703][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5096) );
  MX4X1 U7526 ( .A(\registers[684][1] ), .B(\registers[685][1] ), .C(
        \registers[686][1] ), .D(\registers[687][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5101) );
  MX4X1 U7527 ( .A(\registers[332][2] ), .B(\registers[333][2] ), .C(
        \registers[334][2] ), .D(\registers[335][2] ), .S0(n7504), .S1(n7743), 
        .Y(n5557) );
  MX4X1 U7528 ( .A(\registers[380][2] ), .B(\registers[381][2] ), .C(
        \registers[382][2] ), .D(\registers[383][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5542) );
  MX4X1 U7529 ( .A(\registers[364][2] ), .B(\registers[365][2] ), .C(
        \registers[366][2] ), .D(\registers[367][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5547) );
  MX4X1 U7530 ( .A(\registers[76][2] ), .B(\registers[77][2] ), .C(
        \registers[78][2] ), .D(\registers[79][2] ), .S0(n7509), .S1(n7748), 
        .Y(n5642) );
  MX4X1 U7531 ( .A(\registers[124][2] ), .B(\registers[125][2] ), .C(
        \registers[126][2] ), .D(\registers[127][2] ), .S0(n7508), .S1(n7747), 
        .Y(n5627) );
  MX4X1 U7532 ( .A(\registers[108][2] ), .B(\registers[109][2] ), .C(
        \registers[110][2] ), .D(\registers[111][2] ), .S0(n7509), .S1(n7747), 
        .Y(n5632) );
  MX4X1 U7533 ( .A(\registers[12][2] ), .B(\registers[13][2] ), .C(
        \registers[14][2] ), .D(\registers[15][2] ), .S0(n7511), .S1(n7749), 
        .Y(n5663) );
  MX4X1 U7534 ( .A(\registers[60][2] ), .B(\registers[61][2] ), .C(
        \registers[62][2] ), .D(\registers[63][2] ), .S0(n7510), .S1(n7748), 
        .Y(n5648) );
  MX4X1 U7535 ( .A(\registers[44][2] ), .B(\registers[45][2] ), .C(
        \registers[46][2] ), .D(\registers[47][2] ), .S0(n7510), .S1(n7748), 
        .Y(n5653) );
  MX4X1 U7536 ( .A(\registers[204][2] ), .B(\registers[205][2] ), .C(
        \registers[206][2] ), .D(\registers[207][2] ), .S0(n7507), .S1(n7745), 
        .Y(n5600) );
  MX4X1 U7537 ( .A(\registers[252][2] ), .B(\registers[253][2] ), .C(
        \registers[254][2] ), .D(\registers[255][2] ), .S0(n7506), .S1(n7744), 
        .Y(n5585) );
  MX4X1 U7538 ( .A(\registers[236][2] ), .B(\registers[237][2] ), .C(
        \registers[238][2] ), .D(\registers[239][2] ), .S0(n7506), .S1(n7744), 
        .Y(n5590) );
  MX4X1 U7539 ( .A(\registers[140][2] ), .B(\registers[141][2] ), .C(
        \registers[142][2] ), .D(\registers[143][2] ), .S0(n7508), .S1(n7746), 
        .Y(n5621) );
  MX4X1 U7540 ( .A(\registers[188][2] ), .B(\registers[189][2] ), .C(
        \registers[190][2] ), .D(\registers[191][2] ), .S0(n7507), .S1(n7745), 
        .Y(n5606) );
  MX4X1 U7541 ( .A(\registers[172][2] ), .B(\registers[173][2] ), .C(
        \registers[174][2] ), .D(\registers[175][2] ), .S0(n7507), .S1(n7746), 
        .Y(n5611) );
  MX4X1 U7542 ( .A(\registers[844][2] ), .B(\registers[845][2] ), .C(
        \registers[846][2] ), .D(\registers[847][2] ), .S0(n7493), .S1(n7733), 
        .Y(n5387) );
  MX4X1 U7543 ( .A(\registers[892][2] ), .B(\registers[893][2] ), .C(
        \registers[894][2] ), .D(\registers[895][2] ), .S0(n7492), .S1(n7732), 
        .Y(n5372) );
  MX4X1 U7544 ( .A(\registers[876][2] ), .B(\registers[877][2] ), .C(
        \registers[878][2] ), .D(\registers[879][2] ), .S0(n7493), .S1(n7732), 
        .Y(n5377) );
  MX4X1 U7545 ( .A(\registers[780][2] ), .B(\registers[781][2] ), .C(
        \registers[782][2] ), .D(\registers[783][2] ), .S0(n7495), .S1(n7734), 
        .Y(n5408) );
  MX4X1 U7546 ( .A(\registers[828][2] ), .B(\registers[829][2] ), .C(
        \registers[830][2] ), .D(\registers[831][2] ), .S0(n7494), .S1(n7733), 
        .Y(n5393) );
  MX4X1 U7547 ( .A(\registers[812][2] ), .B(\registers[813][2] ), .C(
        \registers[814][2] ), .D(\registers[815][2] ), .S0(n7494), .S1(n7733), 
        .Y(n5398) );
  MX4X1 U7548 ( .A(\registers[972][2] ), .B(\registers[973][2] ), .C(
        \registers[974][2] ), .D(\registers[975][2] ), .S0(n7491), .S1(n7730), 
        .Y(n5345) );
  MX4X1 U7549 ( .A(\registers[1020][2] ), .B(\registers[1021][2] ), .C(
        \registers[1022][2] ), .D(\registers[1023][2] ), .S0(n7490), .S1(n7729), .Y(n5330) );
  MX4X1 U7550 ( .A(\registers[1004][2] ), .B(\registers[1005][2] ), .C(
        \registers[1006][2] ), .D(\registers[1007][2] ), .S0(n7490), .S1(n7730), .Y(n5335) );
  MX4X1 U7551 ( .A(\registers[908][2] ), .B(\registers[909][2] ), .C(
        \registers[910][2] ), .D(\registers[911][2] ), .S0(n7492), .S1(n7732), 
        .Y(n5366) );
  MX4X1 U7552 ( .A(\registers[956][2] ), .B(\registers[957][2] ), .C(
        \registers[958][2] ), .D(\registers[959][2] ), .S0(n7491), .S1(n7731), 
        .Y(n5351) );
  MX4X1 U7553 ( .A(\registers[940][2] ), .B(\registers[941][2] ), .C(
        \registers[942][2] ), .D(\registers[943][2] ), .S0(n7491), .S1(n7731), 
        .Y(n5356) );
  MX4X1 U7554 ( .A(\registers[588][2] ), .B(\registers[589][2] ), .C(
        \registers[590][2] ), .D(\registers[591][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5472) );
  MX4X1 U7555 ( .A(\registers[636][2] ), .B(\registers[637][2] ), .C(
        \registers[638][2] ), .D(\registers[639][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5457) );
  MX4X1 U7556 ( .A(\registers[620][2] ), .B(\registers[621][2] ), .C(
        \registers[622][2] ), .D(\registers[623][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5462) );
  MX4X1 U7557 ( .A(\registers[524][2] ), .B(\registers[525][2] ), .C(
        \registers[526][2] ), .D(\registers[527][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5493) );
  MX4X1 U7558 ( .A(\registers[572][2] ), .B(\registers[573][2] ), .C(
        \registers[574][2] ), .D(\registers[575][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5478) );
  MX4X1 U7559 ( .A(\registers[556][2] ), .B(\registers[557][2] ), .C(
        \registers[558][2] ), .D(\registers[559][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5483) );
  MX4X1 U7560 ( .A(\registers[716][2] ), .B(\registers[717][2] ), .C(
        \registers[718][2] ), .D(\registers[719][2] ), .S0(n7496), .S1(n7735), 
        .Y(n5430) );
  MX4X1 U7561 ( .A(\registers[764][2] ), .B(\registers[765][2] ), .C(
        \registers[766][2] ), .D(\registers[767][2] ), .S0(n7495), .S1(n7734), 
        .Y(n5415) );
  MX4X1 U7562 ( .A(\registers[748][2] ), .B(\registers[749][2] ), .C(
        \registers[750][2] ), .D(\registers[751][2] ), .S0(n7495), .S1(n7735), 
        .Y(n5420) );
  MX4X1 U7563 ( .A(\registers[652][2] ), .B(\registers[653][2] ), .C(
        \registers[654][2] ), .D(\registers[655][2] ), .S0(n7497), .S1(n7736), 
        .Y(n5451) );
  MX4X1 U7564 ( .A(\registers[700][2] ), .B(\registers[701][2] ), .C(
        \registers[702][2] ), .D(\registers[703][2] ), .S0(n7496), .S1(n7736), 
        .Y(n5436) );
  MX4X1 U7565 ( .A(\registers[684][2] ), .B(\registers[685][2] ), .C(
        \registers[686][2] ), .D(\registers[687][2] ), .S0(n7497), .S1(n7736), 
        .Y(n5441) );
  MX4X1 U7566 ( .A(\registers[332][3] ), .B(\registers[333][3] ), .C(
        \registers[334][3] ), .D(\registers[335][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5897) );
  MX4X1 U7567 ( .A(\registers[380][3] ), .B(\registers[381][3] ), .C(
        \registers[382][3] ), .D(\registers[383][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5882) );
  MX4X1 U7568 ( .A(\registers[364][3] ), .B(\registers[365][3] ), .C(
        \registers[366][3] ), .D(\registers[367][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5887) );
  MX4X1 U7569 ( .A(\registers[76][3] ), .B(\registers[77][3] ), .C(
        \registers[78][3] ), .D(\registers[79][3] ), .S0(n7531), .S1(n7767), 
        .Y(n5982) );
  MX4X1 U7570 ( .A(\registers[124][3] ), .B(\registers[125][3] ), .C(
        \registers[126][3] ), .D(\registers[127][3] ), .S0(n7530), .S1(n7766), 
        .Y(n5967) );
  MX4X1 U7571 ( .A(\registers[108][3] ), .B(\registers[109][3] ), .C(
        \registers[110][3] ), .D(\registers[111][3] ), .S0(n7530), .S1(n7767), 
        .Y(n5972) );
  MX4X1 U7572 ( .A(\registers[12][3] ), .B(\registers[13][3] ), .C(
        \registers[14][3] ), .D(\registers[15][3] ), .S0(n7532), .S1(n7768), 
        .Y(n6003) );
  MX4X1 U7573 ( .A(\registers[60][3] ), .B(\registers[61][3] ), .C(
        \registers[62][3] ), .D(\registers[63][3] ), .S0(n7531), .S1(n7768), 
        .Y(n5988) );
  MX4X1 U7574 ( .A(\registers[44][3] ), .B(\registers[45][3] ), .C(
        \registers[46][3] ), .D(\registers[47][3] ), .S0(n7531), .S1(n7768), 
        .Y(n5993) );
  MX4X1 U7575 ( .A(\registers[204][3] ), .B(\registers[205][3] ), .C(
        \registers[206][3] ), .D(\registers[207][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5940) );
  MX4X1 U7576 ( .A(\registers[252][3] ), .B(\registers[253][3] ), .C(
        \registers[254][3] ), .D(\registers[255][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5925) );
  MX4X1 U7577 ( .A(\registers[236][3] ), .B(\registers[237][3] ), .C(
        \registers[238][3] ), .D(\registers[239][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5930) );
  MX4X1 U7578 ( .A(\registers[140][3] ), .B(\registers[141][3] ), .C(
        \registers[142][3] ), .D(\registers[143][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5961) );
  MX4X1 U7579 ( .A(\registers[188][3] ), .B(\registers[189][3] ), .C(
        \registers[190][3] ), .D(\registers[191][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5946) );
  MX4X1 U7580 ( .A(\registers[172][3] ), .B(\registers[173][3] ), .C(
        \registers[174][3] ), .D(\registers[175][3] ), .S0(n7529), .S1(n7765), 
        .Y(n5951) );
  MX4X1 U7581 ( .A(\registers[844][3] ), .B(\registers[845][3] ), .C(
        \registers[846][3] ), .D(\registers[847][3] ), .S0(n7515), .S1(n7752), 
        .Y(n5727) );
  MX4X1 U7582 ( .A(\registers[892][3] ), .B(\registers[893][3] ), .C(
        \registers[894][3] ), .D(\registers[895][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5712) );
  MX4X1 U7583 ( .A(\registers[876][3] ), .B(\registers[877][3] ), .C(
        \registers[878][3] ), .D(\registers[879][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5717) );
  MX4X1 U7584 ( .A(\registers[780][3] ), .B(\registers[781][3] ), .C(
        \registers[782][3] ), .D(\registers[783][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5748) );
  MX4X1 U7585 ( .A(\registers[828][3] ), .B(\registers[829][3] ), .C(
        \registers[830][3] ), .D(\registers[831][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5733) );
  MX4X1 U7586 ( .A(\registers[812][3] ), .B(\registers[813][3] ), .C(
        \registers[814][3] ), .D(\registers[815][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5738) );
  MX4X1 U7587 ( .A(\registers[972][3] ), .B(\registers[973][3] ), .C(
        \registers[974][3] ), .D(\registers[975][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5685) );
  MX4X1 U7588 ( .A(\registers[1020][3] ), .B(\registers[1021][3] ), .C(
        \registers[1022][3] ), .D(\registers[1023][3] ), .S0(n7511), .S1(n7749), .Y(n5670) );
  MX4X1 U7589 ( .A(\registers[1004][3] ), .B(\registers[1005][3] ), .C(
        \registers[1006][3] ), .D(\registers[1007][3] ), .S0(n7511), .S1(n7749), .Y(n5675) );
  MX4X1 U7590 ( .A(\registers[908][3] ), .B(\registers[909][3] ), .C(
        \registers[910][3] ), .D(\registers[911][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5706) );
  MX4X1 U7591 ( .A(\registers[956][3] ), .B(\registers[957][3] ), .C(
        \registers[958][3] ), .D(\registers[959][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5691) );
  MX4X1 U7592 ( .A(\registers[940][3] ), .B(\registers[941][3] ), .C(
        \registers[942][3] ), .D(\registers[943][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5696) );
  MX4X1 U7593 ( .A(\registers[588][3] ), .B(\registers[589][3] ), .C(
        \registers[590][3] ), .D(\registers[591][3] ), .S0(n7520), .S1(n7757), 
        .Y(n5812) );
  MX4X1 U7594 ( .A(\registers[636][3] ), .B(\registers[637][3] ), .C(
        \registers[638][3] ), .D(\registers[639][3] ), .S0(n7519), .S1(n7756), 
        .Y(n5797) );
  MX4X1 U7595 ( .A(\registers[620][3] ), .B(\registers[621][3] ), .C(
        \registers[622][3] ), .D(\registers[623][3] ), .S0(n7519), .S1(n7757), 
        .Y(n5802) );
  MX4X1 U7596 ( .A(\registers[524][3] ), .B(\registers[525][3] ), .C(
        \registers[526][3] ), .D(\registers[527][3] ), .S0(n7521), .S1(n7759), 
        .Y(n5833) );
  MX4X1 U7597 ( .A(\registers[572][3] ), .B(\registers[573][3] ), .C(
        \registers[574][3] ), .D(\registers[575][3] ), .S0(n7520), .S1(n7758), 
        .Y(n5818) );
  MX4X1 U7598 ( .A(\registers[556][3] ), .B(\registers[557][3] ), .C(
        \registers[558][3] ), .D(\registers[559][3] ), .S0(n7521), .S1(n7758), 
        .Y(n5823) );
  MX4X1 U7599 ( .A(\registers[716][3] ), .B(\registers[717][3] ), .C(
        \registers[718][3] ), .D(\registers[719][3] ), .S0(n7517), .S1(n7755), 
        .Y(n5770) );
  MX4X1 U7600 ( .A(\registers[764][3] ), .B(\registers[765][3] ), .C(
        \registers[766][3] ), .D(\registers[767][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5755) );
  MX4X1 U7601 ( .A(\registers[748][3] ), .B(\registers[749][3] ), .C(
        \registers[750][3] ), .D(\registers[751][3] ), .S0(n7517), .S1(n7754), 
        .Y(n5760) );
  MX4X1 U7602 ( .A(\registers[652][3] ), .B(\registers[653][3] ), .C(
        \registers[654][3] ), .D(\registers[655][3] ), .S0(n7519), .S1(n7756), 
        .Y(n5791) );
  MX4X1 U7603 ( .A(\registers[700][3] ), .B(\registers[701][3] ), .C(
        \registers[702][3] ), .D(\registers[703][3] ), .S0(n7518), .S1(n7755), 
        .Y(n5776) );
  MX4X1 U7604 ( .A(\registers[684][3] ), .B(\registers[685][3] ), .C(
        \registers[686][3] ), .D(\registers[687][3] ), .S0(n7518), .S1(n7756), 
        .Y(n5781) );
  MX4X1 U7605 ( .A(\registers[332][4] ), .B(\registers[333][4] ), .C(
        \registers[334][4] ), .D(\registers[335][4] ), .S0(n7547), .S1(n7782), 
        .Y(n6237) );
  MX4X1 U7606 ( .A(\registers[380][4] ), .B(\registers[381][4] ), .C(
        \registers[382][4] ), .D(\registers[383][4] ), .S0(n7546), .S1(n7781), 
        .Y(n6222) );
  MX4X1 U7607 ( .A(\registers[364][4] ), .B(\registers[365][4] ), .C(
        \registers[366][4] ), .D(\registers[367][4] ), .S0(n7546), .S1(n7781), 
        .Y(n6227) );
  MX4X1 U7608 ( .A(\registers[76][4] ), .B(\registers[77][4] ), .C(
        \registers[78][4] ), .D(\registers[79][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6322) );
  MX4X1 U7609 ( .A(\registers[124][4] ), .B(\registers[125][4] ), .C(
        \registers[126][4] ), .D(\registers[127][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6307) );
  MX4X1 U7610 ( .A(\registers[108][4] ), .B(\registers[109][4] ), .C(
        \registers[110][4] ), .D(\registers[111][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6312) );
  MX4X1 U7611 ( .A(\registers[12][4] ), .B(\registers[13][4] ), .C(
        \registers[14][4] ), .D(\registers[15][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6343) );
  MX4X1 U7612 ( .A(\registers[60][4] ), .B(\registers[61][4] ), .C(
        \registers[62][4] ), .D(\registers[63][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6328) );
  MX4X1 U7613 ( .A(\registers[44][4] ), .B(\registers[45][4] ), .C(
        \registers[46][4] ), .D(\registers[47][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6333) );
  MX4X1 U7614 ( .A(\registers[204][4] ), .B(\registers[205][4] ), .C(
        \registers[206][4] ), .D(\registers[207][4] ), .S0(n7549), .S1(n7784), 
        .Y(n6280) );
  MX4X1 U7615 ( .A(\registers[252][4] ), .B(\registers[253][4] ), .C(
        \registers[254][4] ), .D(\registers[255][4] ), .S0(n7548), .S1(n7784), 
        .Y(n6265) );
  MX4X1 U7616 ( .A(\registers[236][4] ), .B(\registers[237][4] ), .C(
        \registers[238][4] ), .D(\registers[239][4] ), .S0(n7549), .S1(n7784), 
        .Y(n6270) );
  MX4X1 U7617 ( .A(\registers[140][4] ), .B(\registers[141][4] ), .C(
        \registers[142][4] ), .D(\registers[143][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6301) );
  MX4X1 U7618 ( .A(\registers[188][4] ), .B(\registers[189][4] ), .C(
        \registers[190][4] ), .D(\registers[191][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6286) );
  MX4X1 U7619 ( .A(\registers[172][4] ), .B(\registers[173][4] ), .C(
        \registers[174][4] ), .D(\registers[175][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6291) );
  MX4X1 U7620 ( .A(\registers[844][4] ), .B(\registers[845][4] ), .C(
        \registers[846][4] ), .D(\registers[847][4] ), .S0(n7536), .S1(n7772), 
        .Y(n6067) );
  MX4X1 U7621 ( .A(\registers[892][4] ), .B(\registers[893][4] ), .C(
        \registers[894][4] ), .D(\registers[895][4] ), .S0(n7535), .S1(n7771), 
        .Y(n6052) );
  MX4X1 U7622 ( .A(\registers[876][4] ), .B(\registers[877][4] ), .C(
        \registers[878][4] ), .D(\registers[879][4] ), .S0(n7535), .S1(n7772), 
        .Y(n6057) );
  MX4X1 U7623 ( .A(\registers[780][4] ), .B(\registers[781][4] ), .C(
        \registers[782][4] ), .D(\registers[783][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6088) );
  MX4X1 U7624 ( .A(\registers[828][4] ), .B(\registers[829][4] ), .C(
        \registers[830][4] ), .D(\registers[831][4] ), .S0(n7536), .S1(n7772), 
        .Y(n6073) );
  MX4X1 U7625 ( .A(\registers[812][4] ), .B(\registers[813][4] ), .C(
        \registers[814][4] ), .D(\registers[815][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6078) );
  MX4X1 U7626 ( .A(\registers[972][4] ), .B(\registers[973][4] ), .C(
        \registers[974][4] ), .D(\registers[975][4] ), .S0(n7533), .S1(n7770), 
        .Y(n6025) );
  MX4X1 U7627 ( .A(\registers[1020][4] ), .B(\registers[1021][4] ), .C(
        \registers[1022][4] ), .D(\registers[1023][4] ), .S0(n7532), .S1(n7769), .Y(n6010) );
  MX4X1 U7628 ( .A(\registers[1004][4] ), .B(\registers[1005][4] ), .C(
        \registers[1006][4] ), .D(\registers[1007][4] ), .S0(n7533), .S1(n7769), .Y(n6015) );
  MX4X1 U7629 ( .A(\registers[908][4] ), .B(\registers[909][4] ), .C(
        \registers[910][4] ), .D(\registers[911][4] ), .S0(n7535), .S1(n7771), 
        .Y(n6046) );
  MX4X1 U7630 ( .A(\registers[956][4] ), .B(\registers[957][4] ), .C(
        \registers[958][4] ), .D(\registers[959][4] ), .S0(n7534), .S1(n7770), 
        .Y(n6031) );
  MX4X1 U7631 ( .A(\registers[940][4] ), .B(\registers[941][4] ), .C(
        \registers[942][4] ), .D(\registers[943][4] ), .S0(n7534), .S1(n7770), 
        .Y(n6036) );
  MX4X1 U7632 ( .A(\registers[588][4] ), .B(\registers[589][4] ), .C(
        \registers[590][4] ), .D(\registers[591][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6152) );
  MX4X1 U7633 ( .A(\registers[636][4] ), .B(\registers[637][4] ), .C(
        \registers[638][4] ), .D(\registers[639][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6137) );
  MX4X1 U7634 ( .A(\registers[620][4] ), .B(\registers[621][4] ), .C(
        \registers[622][4] ), .D(\registers[623][4] ), .S0(n7541), .S1(n7776), 
        .Y(n6142) );
  MX4X1 U7635 ( .A(\registers[524][4] ), .B(\registers[525][4] ), .C(
        \registers[526][4] ), .D(\registers[527][4] ), .S0(n7543), .S1(n7778), 
        .Y(n6173) );
  MX4X1 U7636 ( .A(\registers[572][4] ), .B(\registers[573][4] ), .C(
        \registers[574][4] ), .D(\registers[575][4] ), .S0(n7542), .S1(n7777), 
        .Y(n6158) );
  MX4X1 U7637 ( .A(\registers[556][4] ), .B(\registers[557][4] ), .C(
        \registers[558][4] ), .D(\registers[559][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6163) );
  MX4X1 U7638 ( .A(\registers[716][4] ), .B(\registers[717][4] ), .C(
        \registers[718][4] ), .D(\registers[719][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6110) );
  MX4X1 U7639 ( .A(\registers[764][4] ), .B(\registers[765][4] ), .C(
        \registers[766][4] ), .D(\registers[767][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6095) );
  MX4X1 U7640 ( .A(\registers[748][4] ), .B(\registers[749][4] ), .C(
        \registers[750][4] ), .D(\registers[751][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6100) );
  MX4X1 U7641 ( .A(\registers[652][4] ), .B(\registers[653][4] ), .C(
        \registers[654][4] ), .D(\registers[655][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6131) );
  MX4X1 U7642 ( .A(\registers[700][4] ), .B(\registers[701][4] ), .C(
        \registers[702][4] ), .D(\registers[703][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6116) );
  MX4X1 U7643 ( .A(\registers[684][4] ), .B(\registers[685][4] ), .C(
        \registers[686][4] ), .D(\registers[687][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6121) );
  MX4X1 U7644 ( .A(\registers[332][5] ), .B(\registers[333][5] ), .C(
        \registers[334][5] ), .D(\registers[335][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6577) );
  MX4X1 U7645 ( .A(\registers[380][5] ), .B(\registers[381][5] ), .C(
        \registers[382][5] ), .D(\registers[383][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6562) );
  MX4X1 U7646 ( .A(\registers[364][5] ), .B(\registers[365][5] ), .C(
        \registers[366][5] ), .D(\registers[367][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6567) );
  MX4X1 U7647 ( .A(\registers[76][5] ), .B(\registers[77][5] ), .C(
        \registers[78][5] ), .D(\registers[79][5] ), .S0(n7573), .S1(n7806), 
        .Y(n6662) );
  MX4X1 U7648 ( .A(\registers[124][5] ), .B(\registers[125][5] ), .C(
        \registers[126][5] ), .D(\registers[127][5] ), .S0(n7572), .S1(n7805), 
        .Y(n6647) );
  MX4X1 U7649 ( .A(\registers[108][5] ), .B(\registers[109][5] ), .C(
        \registers[110][5] ), .D(\registers[111][5] ), .S0(n7573), .S1(n7805), 
        .Y(n6652) );
  MX4X1 U7650 ( .A(\registers[12][5] ), .B(\registers[13][5] ), .C(
        \registers[14][5] ), .D(\registers[15][5] ), .S0(n7575), .S1(n7807), 
        .Y(n6683) );
  MX4X1 U7651 ( .A(\registers[60][5] ), .B(\registers[61][5] ), .C(
        \registers[62][5] ), .D(\registers[63][5] ), .S0(n7574), .S1(n7806), 
        .Y(n6668) );
  MX4X1 U7652 ( .A(\registers[44][5] ), .B(\registers[45][5] ), .C(
        \registers[46][5] ), .D(\registers[47][5] ), .S0(n7574), .S1(n7806), 
        .Y(n6673) );
  MX4X1 U7653 ( .A(\registers[204][5] ), .B(\registers[205][5] ), .C(
        \registers[206][5] ), .D(\registers[207][5] ), .S0(n7571), .S1(n7704), 
        .Y(n6620) );
  MX4X1 U7654 ( .A(\registers[252][5] ), .B(\registers[253][5] ), .C(
        \registers[254][5] ), .D(\registers[255][5] ), .S0(n7570), .S1(n7803), 
        .Y(n6605) );
  MX4X1 U7655 ( .A(\registers[236][5] ), .B(\registers[237][5] ), .C(
        \registers[238][5] ), .D(\registers[239][5] ), .S0(n7570), .S1(n7696), 
        .Y(n6610) );
  MX4X1 U7656 ( .A(\registers[140][5] ), .B(\registers[141][5] ), .C(
        \registers[142][5] ), .D(\registers[143][5] ), .S0(n7572), .S1(n7804), 
        .Y(n6641) );
  MX4X1 U7657 ( .A(\registers[188][5] ), .B(\registers[189][5] ), .C(
        \registers[190][5] ), .D(\registers[191][5] ), .S0(n7571), .S1(n7699), 
        .Y(n6626) );
  MX4X1 U7658 ( .A(\registers[172][5] ), .B(\registers[173][5] ), .C(
        \registers[174][5] ), .D(\registers[175][5] ), .S0(n7571), .S1(n7804), 
        .Y(n6631) );
  MX4X1 U7659 ( .A(\registers[844][5] ), .B(\registers[845][5] ), .C(
        \registers[846][5] ), .D(\registers[847][5] ), .S0(n7557), .S1(n7792), 
        .Y(n6407) );
  MX4X1 U7660 ( .A(\registers[892][5] ), .B(\registers[893][5] ), .C(
        \registers[894][5] ), .D(\registers[895][5] ), .S0(n7556), .S1(n7791), 
        .Y(n6392) );
  MX4X1 U7661 ( .A(\registers[876][5] ), .B(\registers[877][5] ), .C(
        \registers[878][5] ), .D(\registers[879][5] ), .S0(n7557), .S1(n7791), 
        .Y(n6397) );
  MX4X1 U7662 ( .A(\registers[780][5] ), .B(\registers[781][5] ), .C(
        \registers[782][5] ), .D(\registers[783][5] ), .S0(n7559), .S1(n7793), 
        .Y(n6428) );
  MX4X1 U7663 ( .A(\registers[828][5] ), .B(\registers[829][5] ), .C(
        \registers[830][5] ), .D(\registers[831][5] ), .S0(n7558), .S1(n7792), 
        .Y(n6413) );
  MX4X1 U7664 ( .A(\registers[812][5] ), .B(\registers[813][5] ), .C(
        \registers[814][5] ), .D(\registers[815][5] ), .S0(n7558), .S1(n7792), 
        .Y(n6418) );
  MX4X1 U7665 ( .A(\registers[972][5] ), .B(\registers[973][5] ), .C(
        \registers[974][5] ), .D(\registers[975][5] ), .S0(n7555), .S1(n7789), 
        .Y(n6365) );
  MX4X1 U7666 ( .A(\registers[1020][5] ), .B(\registers[1021][5] ), .C(
        \registers[1022][5] ), .D(\registers[1023][5] ), .S0(n7554), .S1(n7788), .Y(n6350) );
  MX4X1 U7667 ( .A(\registers[1004][5] ), .B(\registers[1005][5] ), .C(
        \registers[1006][5] ), .D(\registers[1007][5] ), .S0(n7554), .S1(n7789), .Y(n6355) );
  MX4X1 U7668 ( .A(\registers[908][5] ), .B(\registers[909][5] ), .C(
        \registers[910][5] ), .D(\registers[911][5] ), .S0(n7556), .S1(n7791), 
        .Y(n6386) );
  MX4X1 U7669 ( .A(\registers[956][5] ), .B(\registers[957][5] ), .C(
        \registers[958][5] ), .D(\registers[959][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6371) );
  MX4X1 U7670 ( .A(\registers[940][5] ), .B(\registers[941][5] ), .C(
        \registers[942][5] ), .D(\registers[943][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6376) );
  MX4X1 U7671 ( .A(\registers[588][5] ), .B(\registers[589][5] ), .C(
        \registers[590][5] ), .D(\registers[591][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6492) );
  MX4X1 U7672 ( .A(\registers[636][5] ), .B(\registers[637][5] ), .C(
        \registers[638][5] ), .D(\registers[639][5] ), .S0(n7562), .S1(n7796), 
        .Y(n6477) );
  MX4X1 U7673 ( .A(\registers[620][5] ), .B(\registers[621][5] ), .C(
        \registers[622][5] ), .D(\registers[623][5] ), .S0(n7562), .S1(n7796), 
        .Y(n6482) );
  MX4X1 U7674 ( .A(\registers[524][5] ), .B(\registers[525][5] ), .C(
        \registers[526][5] ), .D(\registers[527][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6513) );
  MX4X1 U7675 ( .A(\registers[572][5] ), .B(\registers[573][5] ), .C(
        \registers[574][5] ), .D(\registers[575][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6498) );
  MX4X1 U7676 ( .A(\registers[556][5] ), .B(\registers[557][5] ), .C(
        \registers[558][5] ), .D(\registers[559][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6503) );
  MX4X1 U7677 ( .A(\registers[716][5] ), .B(\registers[717][5] ), .C(
        \registers[718][5] ), .D(\registers[719][5] ), .S0(n7560), .S1(n7794), 
        .Y(n6450) );
  MX4X1 U7678 ( .A(\registers[764][5] ), .B(\registers[765][5] ), .C(
        \registers[766][5] ), .D(\registers[767][5] ), .S0(n7559), .S1(n7793), 
        .Y(n6435) );
  MX4X1 U7679 ( .A(\registers[748][5] ), .B(\registers[749][5] ), .C(
        \registers[750][5] ), .D(\registers[751][5] ), .S0(n7559), .S1(n7794), 
        .Y(n6440) );
  MX4X1 U7680 ( .A(\registers[652][5] ), .B(\registers[653][5] ), .C(
        \registers[654][5] ), .D(\registers[655][5] ), .S0(n7561), .S1(n7796), 
        .Y(n6471) );
  MX4X1 U7681 ( .A(\registers[700][5] ), .B(\registers[701][5] ), .C(
        \registers[702][5] ), .D(\registers[703][5] ), .S0(n7560), .S1(n7795), 
        .Y(n6456) );
  MX4X1 U7682 ( .A(\registers[684][5] ), .B(\registers[685][5] ), .C(
        \registers[686][5] ), .D(\registers[687][5] ), .S0(n7561), .S1(n7795), 
        .Y(n6461) );
  MX4X1 U7683 ( .A(\registers[332][6] ), .B(\registers[333][6] ), .C(
        \registers[334][6] ), .D(\registers[335][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6917) );
  MX4X1 U7684 ( .A(\registers[380][6] ), .B(\registers[381][6] ), .C(
        \registers[382][6] ), .D(\registers[383][6] ), .S0(n7588), .S1(n7819), 
        .Y(n6902) );
  MX4X1 U7685 ( .A(\registers[364][6] ), .B(\registers[365][6] ), .C(
        \registers[366][6] ), .D(\registers[367][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6907) );
  MX4X1 U7686 ( .A(\registers[76][6] ), .B(\registers[77][6] ), .C(
        \registers[78][6] ), .D(\registers[79][6] ), .S0(n7595), .S1(n7825), 
        .Y(n7002) );
  MX4X1 U7687 ( .A(\registers[124][6] ), .B(\registers[125][6] ), .C(
        \registers[126][6] ), .D(\registers[127][6] ), .S0(n7594), .S1(n7824), 
        .Y(n6987) );
  MX4X1 U7688 ( .A(\registers[108][6] ), .B(\registers[109][6] ), .C(
        \registers[110][6] ), .D(\registers[111][6] ), .S0(n7594), .S1(n7825), 
        .Y(n6992) );
  MX4X1 U7689 ( .A(\registers[12][6] ), .B(\registers[13][6] ), .C(
        \registers[14][6] ), .D(\registers[15][6] ), .S0(n7596), .S1(n7827), 
        .Y(n7023) );
  MX4X1 U7690 ( .A(\registers[60][6] ), .B(\registers[61][6] ), .C(
        \registers[62][6] ), .D(\registers[63][6] ), .S0(n7595), .S1(n7826), 
        .Y(n7008) );
  MX4X1 U7691 ( .A(\registers[44][6] ), .B(\registers[45][6] ), .C(
        \registers[46][6] ), .D(\registers[47][6] ), .S0(n7595), .S1(n7826), 
        .Y(n7013) );
  MX4X1 U7692 ( .A(\registers[204][6] ), .B(\registers[205][6] ), .C(
        \registers[206][6] ), .D(\registers[207][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6960) );
  MX4X1 U7693 ( .A(\registers[252][6] ), .B(\registers[253][6] ), .C(
        \registers[254][6] ), .D(\registers[255][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6945) );
  MX4X1 U7694 ( .A(\registers[236][6] ), .B(\registers[237][6] ), .C(
        \registers[238][6] ), .D(\registers[239][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6950) );
  MX4X1 U7695 ( .A(\registers[140][6] ), .B(\registers[141][6] ), .C(
        \registers[142][6] ), .D(\registers[143][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6981) );
  MX4X1 U7696 ( .A(\registers[188][6] ), .B(\registers[189][6] ), .C(
        \registers[190][6] ), .D(\registers[191][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6966) );
  MX4X1 U7697 ( .A(\registers[172][6] ), .B(\registers[173][6] ), .C(
        \registers[174][6] ), .D(\registers[175][6] ), .S0(n7593), .S1(n7823), 
        .Y(n6971) );
  MX4X1 U7698 ( .A(\registers[844][6] ), .B(\registers[845][6] ), .C(
        \registers[846][6] ), .D(\registers[847][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6747) );
  MX4X1 U7699 ( .A(\registers[892][6] ), .B(\registers[893][6] ), .C(
        \registers[894][6] ), .D(\registers[895][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6732) );
  MX4X1 U7700 ( .A(\registers[876][6] ), .B(\registers[877][6] ), .C(
        \registers[878][6] ), .D(\registers[879][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6737) );
  MX4X1 U7701 ( .A(\registers[780][6] ), .B(\registers[781][6] ), .C(
        \registers[782][6] ), .D(\registers[783][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6768) );
  MX4X1 U7702 ( .A(\registers[828][6] ), .B(\registers[829][6] ), .C(
        \registers[830][6] ), .D(\registers[831][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6753) );
  MX4X1 U7703 ( .A(\registers[812][6] ), .B(\registers[813][6] ), .C(
        \registers[814][6] ), .D(\registers[815][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6758) );
  MX4X1 U7704 ( .A(\registers[972][6] ), .B(\registers[973][6] ), .C(
        \registers[974][6] ), .D(\registers[975][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6705) );
  MX4X1 U7705 ( .A(\registers[1020][6] ), .B(\registers[1021][6] ), .C(
        \registers[1022][6] ), .D(\registers[1023][6] ), .S0(n7575), .S1(n7807), .Y(n6690) );
  MX4X1 U7706 ( .A(\registers[1004][6] ), .B(\registers[1005][6] ), .C(
        \registers[1006][6] ), .D(\registers[1007][6] ), .S0(n7575), .S1(n7807), .Y(n6695) );
  MX4X1 U7707 ( .A(\registers[908][6] ), .B(\registers[909][6] ), .C(
        \registers[910][6] ), .D(\registers[911][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6726) );
  MX4X1 U7708 ( .A(\registers[956][6] ), .B(\registers[957][6] ), .C(
        \registers[958][6] ), .D(\registers[959][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6711) );
  MX4X1 U7709 ( .A(\registers[940][6] ), .B(\registers[941][6] ), .C(
        \registers[942][6] ), .D(\registers[943][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6716) );
  MX4X1 U7710 ( .A(\registers[588][6] ), .B(\registers[589][6] ), .C(
        \registers[590][6] ), .D(\registers[591][6] ), .S0(n7584), .S1(n7815), 
        .Y(n6832) );
  MX4X1 U7711 ( .A(\registers[636][6] ), .B(\registers[637][6] ), .C(
        \registers[638][6] ), .D(\registers[639][6] ), .S0(n7583), .S1(n7815), 
        .Y(n6817) );
  MX4X1 U7712 ( .A(\registers[620][6] ), .B(\registers[621][6] ), .C(
        \registers[622][6] ), .D(\registers[623][6] ), .S0(n7583), .S1(n7815), 
        .Y(n6822) );
  MX4X1 U7713 ( .A(\registers[524][6] ), .B(\registers[525][6] ), .C(
        \registers[526][6] ), .D(\registers[527][6] ), .S0(n7585), .S1(n7817), 
        .Y(n6853) );
  MX4X1 U7714 ( .A(\registers[572][6] ), .B(\registers[573][6] ), .C(
        \registers[574][6] ), .D(\registers[575][6] ), .S0(n7584), .S1(n7816), 
        .Y(n6838) );
  MX4X1 U7715 ( .A(\registers[556][6] ), .B(\registers[557][6] ), .C(
        \registers[558][6] ), .D(\registers[559][6] ), .S0(n7585), .S1(n7816), 
        .Y(n6843) );
  MX4X1 U7716 ( .A(\registers[716][6] ), .B(\registers[717][6] ), .C(
        \registers[718][6] ), .D(\registers[719][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6790) );
  MX4X1 U7717 ( .A(\registers[764][6] ), .B(\registers[765][6] ), .C(
        \registers[766][6] ), .D(\registers[767][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6775) );
  MX4X1 U7718 ( .A(\registers[748][6] ), .B(\registers[749][6] ), .C(
        \registers[750][6] ), .D(\registers[751][6] ), .S0(n7581), .S1(n7812), 
        .Y(n6780) );
  MX4X1 U7719 ( .A(\registers[652][6] ), .B(\registers[653][6] ), .C(
        \registers[654][6] ), .D(\registers[655][6] ), .S0(n7583), .S1(n7814), 
        .Y(n6811) );
  MX4X1 U7720 ( .A(\registers[700][6] ), .B(\registers[701][6] ), .C(
        \registers[702][6] ), .D(\registers[703][6] ), .S0(n7582), .S1(n7813), 
        .Y(n6796) );
  MX4X1 U7721 ( .A(\registers[684][6] ), .B(\registers[685][6] ), .C(
        \registers[686][6] ), .D(\registers[687][6] ), .S0(n7582), .S1(n7814), 
        .Y(n6801) );
  MX4X1 U7722 ( .A(\registers[332][7] ), .B(\registers[333][7] ), .C(
        \registers[334][7] ), .D(\registers[335][7] ), .S0(n7611), .S1(n7840), 
        .Y(n7257) );
  MX4X1 U7723 ( .A(\registers[380][7] ), .B(\registers[381][7] ), .C(
        \registers[382][7] ), .D(\registers[383][7] ), .S0(n7610), .S1(n7839), 
        .Y(n7242) );
  MX4X1 U7724 ( .A(\registers[364][7] ), .B(\registers[365][7] ), .C(
        \registers[366][7] ), .D(\registers[367][7] ), .S0(n7610), .S1(n7839), 
        .Y(n7247) );
  MX4X1 U7725 ( .A(\registers[204][7] ), .B(\registers[205][7] ), .C(
        \registers[206][7] ), .D(\registers[207][7] ), .S0(n7613), .S1(n7843), 
        .Y(n7300) );
  MX4X1 U7726 ( .A(\registers[252][7] ), .B(\registers[253][7] ), .C(
        \registers[254][7] ), .D(\registers[255][7] ), .S0(n7612), .S1(n7842), 
        .Y(n7285) );
  MX4X1 U7727 ( .A(\registers[236][7] ), .B(\registers[237][7] ), .C(
        \registers[238][7] ), .D(\registers[239][7] ), .S0(n7613), .S1(n7842), 
        .Y(n7290) );
  MX4X1 U7728 ( .A(\registers[76][7] ), .B(\registers[77][7] ), .C(
        \registers[78][7] ), .D(\registers[79][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7342) );
  MX4X1 U7729 ( .A(\registers[124][7] ), .B(\registers[125][7] ), .C(
        \registers[126][7] ), .D(\registers[127][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7327) );
  MX4X1 U7730 ( .A(\registers[108][7] ), .B(\registers[109][7] ), .C(
        \registers[110][7] ), .D(\registers[111][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7332) );
  MX4X1 U7731 ( .A(\registers[12][7] ), .B(\registers[13][7] ), .C(
        \registers[14][7] ), .D(\registers[15][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7363) );
  MX4X1 U7732 ( .A(\registers[60][7] ), .B(\registers[61][7] ), .C(
        \registers[62][7] ), .D(\registers[63][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7348) );
  MX4X1 U7733 ( .A(\registers[44][7] ), .B(\registers[45][7] ), .C(
        \registers[46][7] ), .D(\registers[47][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7353) );
  MX4X1 U7734 ( .A(\registers[140][7] ), .B(\registers[141][7] ), .C(
        \registers[142][7] ), .D(\registers[143][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7321) );
  MX4X1 U7735 ( .A(\registers[188][7] ), .B(\registers[189][7] ), .C(
        \registers[190][7] ), .D(\registers[191][7] ), .S0(n7614), .S1(n7843), 
        .Y(n7306) );
  MX4X1 U7736 ( .A(\registers[172][7] ), .B(\registers[173][7] ), .C(
        \registers[174][7] ), .D(\registers[175][7] ), .S0(n7614), .S1(n7843), 
        .Y(n7311) );
  MX4X1 U7737 ( .A(\registers[844][7] ), .B(\registers[845][7] ), .C(
        \registers[846][7] ), .D(\registers[847][7] ), .S0(n7600), .S1(n7830), 
        .Y(n7087) );
  MX4X1 U7738 ( .A(\registers[892][7] ), .B(\registers[893][7] ), .C(
        \registers[894][7] ), .D(\registers[895][7] ), .S0(n7599), .S1(n7829), 
        .Y(n7072) );
  MX4X1 U7739 ( .A(\registers[876][7] ), .B(\registers[877][7] ), .C(
        \registers[878][7] ), .D(\registers[879][7] ), .S0(n7599), .S1(n7830), 
        .Y(n7077) );
  MX4X1 U7740 ( .A(\registers[780][7] ), .B(\registers[781][7] ), .C(
        \registers[782][7] ), .D(\registers[783][7] ), .S0(n7601), .S1(n7831), 
        .Y(n7108) );
  MX4X1 U7741 ( .A(\registers[828][7] ), .B(\registers[829][7] ), .C(
        \registers[830][7] ), .D(\registers[831][7] ), .S0(n7600), .S1(n7831), 
        .Y(n7093) );
  MX4X1 U7742 ( .A(\registers[812][7] ), .B(\registers[813][7] ), .C(
        \registers[814][7] ), .D(\registers[815][7] ), .S0(n7601), .S1(n7831), 
        .Y(n7098) );
  MX4X1 U7743 ( .A(\registers[972][7] ), .B(\registers[973][7] ), .C(
        \registers[974][7] ), .D(\registers[975][7] ), .S0(n7597), .S1(n7828), 
        .Y(n7045) );
  MX4X1 U7744 ( .A(\registers[1020][7] ), .B(\registers[1021][7] ), .C(
        \registers[1022][7] ), .D(\registers[1023][7] ), .S0(n7596), .S1(n7827), .Y(n7030) );
  MX4X1 U7745 ( .A(\registers[1004][7] ), .B(\registers[1005][7] ), .C(
        \registers[1006][7] ), .D(\registers[1007][7] ), .S0(n7597), .S1(n7827), .Y(n7035) );
  MX4X1 U7746 ( .A(\registers[908][7] ), .B(\registers[909][7] ), .C(
        \registers[910][7] ), .D(\registers[911][7] ), .S0(n7599), .S1(n7829), 
        .Y(n7066) );
  MX4X1 U7747 ( .A(\registers[956][7] ), .B(\registers[957][7] ), .C(
        \registers[958][7] ), .D(\registers[959][7] ), .S0(n7598), .S1(n7828), 
        .Y(n7051) );
  MX4X1 U7748 ( .A(\registers[940][7] ), .B(\registers[941][7] ), .C(
        \registers[942][7] ), .D(\registers[943][7] ), .S0(n7598), .S1(n7828), 
        .Y(n7056) );
  MX4X1 U7749 ( .A(\registers[588][7] ), .B(\registers[589][7] ), .C(
        \registers[590][7] ), .D(\registers[591][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7172) );
  MX4X1 U7750 ( .A(\registers[636][7] ), .B(\registers[637][7] ), .C(
        \registers[638][7] ), .D(\registers[639][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7157) );
  MX4X1 U7751 ( .A(\registers[620][7] ), .B(\registers[621][7] ), .C(
        \registers[622][7] ), .D(\registers[623][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7162) );
  MX4X1 U7752 ( .A(\registers[524][7] ), .B(\registers[525][7] ), .C(
        \registers[526][7] ), .D(\registers[527][7] ), .S0(n7607), .S1(n7836), 
        .Y(n7193) );
  MX4X1 U7753 ( .A(\registers[572][7] ), .B(\registers[573][7] ), .C(
        \registers[574][7] ), .D(\registers[575][7] ), .S0(n7606), .S1(n7835), 
        .Y(n7178) );
  MX4X1 U7754 ( .A(\registers[556][7] ), .B(\registers[557][7] ), .C(
        \registers[558][7] ), .D(\registers[559][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7183) );
  MX4X1 U7755 ( .A(\registers[716][7] ), .B(\registers[717][7] ), .C(
        \registers[718][7] ), .D(\registers[719][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7130) );
  MX4X1 U7756 ( .A(\registers[764][7] ), .B(\registers[765][7] ), .C(
        \registers[766][7] ), .D(\registers[767][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7115) );
  MX4X1 U7757 ( .A(\registers[748][7] ), .B(\registers[749][7] ), .C(
        \registers[750][7] ), .D(\registers[751][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7120) );
  MX4X1 U7758 ( .A(\registers[652][7] ), .B(\registers[653][7] ), .C(
        \registers[654][7] ), .D(\registers[655][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7151) );
  MX4X1 U7759 ( .A(\registers[700][7] ), .B(\registers[701][7] ), .C(
        \registers[702][7] ), .D(\registers[703][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7136) );
  MX4X1 U7760 ( .A(\registers[684][7] ), .B(\registers[685][7] ), .C(
        \registers[686][7] ), .D(\registers[687][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7141) );
  MX4X1 U7761 ( .A(n1454), .B(n1452), .C(n1453), .D(n1451), .S0(n4587), .S1(
        n4529), .Y(n1455) );
  MX4X1 U7762 ( .A(\registers[264][0] ), .B(\registers[265][0] ), .C(
        \registers[266][0] ), .D(\registers[267][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1452) );
  MX4X1 U7763 ( .A(\registers[268][0] ), .B(\registers[269][0] ), .C(
        \registers[270][0] ), .D(\registers[271][0] ), .S0(n4120), .S1(n4360), 
        .Y(n1451) );
  MX4X1 U7764 ( .A(\registers[256][0] ), .B(\registers[257][0] ), .C(
        \registers[258][0] ), .D(\registers[259][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1454) );
  MX4X1 U7765 ( .A(n1439), .B(n1436), .C(n1438), .D(n1434), .S0(n4587), .S1(
        n4529), .Y(n1440) );
  MX4X1 U7766 ( .A(\registers[312][0] ), .B(\registers[313][0] ), .C(
        \registers[314][0] ), .D(\registers[315][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1436) );
  MX4X1 U7767 ( .A(\registers[316][0] ), .B(\registers[317][0] ), .C(
        \registers[318][0] ), .D(\registers[319][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1434) );
  MX4X1 U7768 ( .A(\registers[304][0] ), .B(\registers[305][0] ), .C(
        \registers[306][0] ), .D(\registers[307][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1439) );
  MX4X1 U7769 ( .A(n1387), .B(n1385), .C(n1386), .D(n1384), .S0(n4612), .S1(
        n4528), .Y(n1388) );
  MX4X1 U7770 ( .A(\registers[456][0] ), .B(\registers[457][0] ), .C(
        \registers[458][0] ), .D(\registers[459][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1385) );
  MX4X1 U7771 ( .A(\registers[460][0] ), .B(\registers[461][0] ), .C(
        \registers[462][0] ), .D(\registers[463][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1384) );
  MX4X1 U7772 ( .A(\registers[448][0] ), .B(\registers[449][0] ), .C(
        \registers[450][0] ), .D(\registers[451][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1387) );
  MX4X1 U7773 ( .A(n1372), .B(n1370), .C(n1371), .D(n1368), .S0(n4599), .S1(
        n4528), .Y(n1373) );
  MX4X1 U7774 ( .A(\registers[504][0] ), .B(\registers[505][0] ), .C(
        \registers[506][0] ), .D(\registers[507][0] ), .S0(n4115), .S1(n4356), 
        .Y(n1370) );
  MX4X1 U7775 ( .A(\registers[508][0] ), .B(\registers[509][0] ), .C(
        \registers[510][0] ), .D(\registers[511][0] ), .S0(n4115), .S1(n4356), 
        .Y(n1368) );
  MX4X1 U7776 ( .A(\registers[496][0] ), .B(\registers[497][0] ), .C(
        \registers[498][0] ), .D(\registers[499][0] ), .S0(n4115), .S1(n4356), 
        .Y(n1372) );
  MX4X1 U7777 ( .A(n1410), .B(n1408), .C(n1409), .D(n1407), .S0(n4591), .S1(
        n4528), .Y(n1411) );
  MX4X1 U7778 ( .A(\registers[392][0] ), .B(\registers[393][0] ), .C(
        \registers[394][0] ), .D(\registers[395][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1408) );
  MX4X1 U7779 ( .A(\registers[396][0] ), .B(\registers[397][0] ), .C(
        \registers[398][0] ), .D(\registers[399][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1407) );
  MX4X1 U7780 ( .A(\registers[384][0] ), .B(\registers[385][0] ), .C(
        \registers[386][0] ), .D(\registers[387][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1410) );
  MX4X1 U7781 ( .A(n1393), .B(n1391), .C(n1392), .D(n1390), .S0(n4594), .S1(
        n4528), .Y(n1394) );
  MX4X1 U7782 ( .A(\registers[440][0] ), .B(\registers[441][0] ), .C(
        \registers[442][0] ), .D(\registers[443][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1391) );
  MX4X1 U7783 ( .A(\registers[444][0] ), .B(\registers[445][0] ), .C(
        \registers[446][0] ), .D(\registers[447][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1390) );
  MX4X1 U7784 ( .A(\registers[432][0] ), .B(\registers[433][0] ), .C(
        \registers[434][0] ), .D(\registers[435][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1393) );
  MX4X1 U7785 ( .A(n1811), .B(n1809), .C(n1810), .D(n1808), .S0(n4592), .S1(
        n4534), .Y(n1812) );
  MX4X1 U7786 ( .A(\registers[264][1] ), .B(\registers[265][1] ), .C(
        \registers[266][1] ), .D(\registers[267][1] ), .S0(n4141), .S1(n4380), 
        .Y(n1809) );
  MX4X1 U7787 ( .A(\registers[268][1] ), .B(\registers[269][1] ), .C(
        \registers[270][1] ), .D(\registers[271][1] ), .S0(n4141), .S1(n4380), 
        .Y(n1808) );
  MX4X1 U7788 ( .A(\registers[256][1] ), .B(\registers[257][1] ), .C(
        \registers[258][1] ), .D(\registers[259][1] ), .S0(n4141), .S1(n4380), 
        .Y(n1811) );
  MX4X1 U7789 ( .A(n1795), .B(n1793), .C(n1794), .D(n1792), .S0(n4592), .S1(
        n4533), .Y(n1796) );
  MX4X1 U7790 ( .A(\registers[312][1] ), .B(\registers[313][1] ), .C(
        \registers[314][1] ), .D(\registers[315][1] ), .S0(n4140), .S1(n4379), 
        .Y(n1793) );
  MX4X1 U7791 ( .A(\registers[316][1] ), .B(\registers[317][1] ), .C(
        \registers[318][1] ), .D(\registers[319][1] ), .S0(n4140), .S1(n4379), 
        .Y(n1792) );
  MX4X1 U7792 ( .A(\registers[304][1] ), .B(\registers[305][1] ), .C(
        \registers[306][1] ), .D(\registers[307][1] ), .S0(n4140), .S1(n4379), 
        .Y(n1795) );
  MX4X1 U7793 ( .A(n1746), .B(n1744), .C(n1745), .D(n1743), .S0(n4591), .S1(
        n4533), .Y(n1747) );
  MX4X1 U7794 ( .A(\registers[456][1] ), .B(\registers[457][1] ), .C(
        \registers[458][1] ), .D(\registers[459][1] ), .S0(n4137), .S1(n4377), 
        .Y(n1744) );
  MX4X1 U7795 ( .A(\registers[460][1] ), .B(\registers[461][1] ), .C(
        \registers[462][1] ), .D(\registers[463][1] ), .S0(n4137), .S1(n4376), 
        .Y(n1743) );
  MX4X1 U7796 ( .A(\registers[448][1] ), .B(\registers[449][1] ), .C(
        \registers[450][1] ), .D(\registers[451][1] ), .S0(n4137), .S1(n4377), 
        .Y(n1746) );
  MX4X1 U7797 ( .A(n1730), .B(n1728), .C(n1729), .D(n1727), .S0(n4591), .S1(
        n4533), .Y(n1731) );
  MX4X1 U7798 ( .A(\registers[504][1] ), .B(\registers[505][1] ), .C(
        \registers[506][1] ), .D(\registers[507][1] ), .S0(n4136), .S1(n4376), 
        .Y(n1728) );
  MX4X1 U7799 ( .A(\registers[508][1] ), .B(\registers[509][1] ), .C(
        \registers[510][1] ), .D(\registers[511][1] ), .S0(n4136), .S1(n4376), 
        .Y(n1727) );
  MX4X1 U7800 ( .A(\registers[496][1] ), .B(\registers[497][1] ), .C(
        \registers[498][1] ), .D(\registers[499][1] ), .S0(n4136), .S1(n4376), 
        .Y(n1730) );
  MX4X1 U7801 ( .A(n1767), .B(n1765), .C(n1766), .D(n1764), .S0(n4591), .S1(
        n4533), .Y(n1768) );
  MX4X1 U7802 ( .A(\registers[392][1] ), .B(\registers[393][1] ), .C(
        \registers[394][1] ), .D(\registers[395][1] ), .S0(n4138), .S1(n4378), 
        .Y(n1765) );
  MX4X1 U7803 ( .A(\registers[396][1] ), .B(\registers[397][1] ), .C(
        \registers[398][1] ), .D(\registers[399][1] ), .S0(n4138), .S1(n4378), 
        .Y(n1764) );
  MX4X1 U7804 ( .A(\registers[384][1] ), .B(\registers[385][1] ), .C(
        \registers[386][1] ), .D(\registers[387][1] ), .S0(n4138), .S1(n4378), 
        .Y(n1767) );
  MX4X1 U7805 ( .A(n1752), .B(n1750), .C(n1751), .D(n1749), .S0(n4591), .S1(
        n4533), .Y(n1753) );
  MX4X1 U7806 ( .A(\registers[440][1] ), .B(\registers[441][1] ), .C(
        \registers[442][1] ), .D(\registers[443][1] ), .S0(n4137), .S1(n4377), 
        .Y(n1750) );
  MX4X1 U7807 ( .A(\registers[444][1] ), .B(\registers[445][1] ), .C(
        \registers[446][1] ), .D(\registers[447][1] ), .S0(n4137), .S1(n4377), 
        .Y(n1749) );
  MX4X1 U7808 ( .A(\registers[432][1] ), .B(\registers[433][1] ), .C(
        \registers[434][1] ), .D(\registers[435][1] ), .S0(n4137), .S1(n4377), 
        .Y(n1752) );
  MX4X1 U7809 ( .A(n2163), .B(n2161), .C(n2162), .D(n2160), .S0(n4597), .S1(
        n4539), .Y(n2164) );
  MX4X1 U7810 ( .A(\registers[264][2] ), .B(\registers[265][2] ), .C(
        \registers[266][2] ), .D(\registers[267][2] ), .S0(n4162), .S1(n4400), 
        .Y(n2161) );
  MX4X1 U7811 ( .A(\registers[268][2] ), .B(\registers[269][2] ), .C(
        \registers[270][2] ), .D(\registers[271][2] ), .S0(n4162), .S1(n4400), 
        .Y(n2160) );
  MX4X1 U7812 ( .A(\registers[256][2] ), .B(\registers[257][2] ), .C(
        \registers[258][2] ), .D(\registers[259][2] ), .S0(n4162), .S1(n4400), 
        .Y(n2163) );
  MX4X1 U7813 ( .A(n2148), .B(n2146), .C(n2147), .D(n2145), .S0(n4597), .S1(
        n4538), .Y(n2149) );
  MX4X1 U7814 ( .A(\registers[312][2] ), .B(\registers[313][2] ), .C(
        \registers[314][2] ), .D(\registers[315][2] ), .S0(n4161), .S1(n4399), 
        .Y(n2146) );
  MX4X1 U7815 ( .A(\registers[316][2] ), .B(\registers[317][2] ), .C(
        \registers[318][2] ), .D(\registers[319][2] ), .S0(n4161), .S1(n4399), 
        .Y(n2145) );
  MX4X1 U7816 ( .A(\registers[304][2] ), .B(\registers[305][2] ), .C(
        \registers[306][2] ), .D(\registers[307][2] ), .S0(n4161), .S1(n4399), 
        .Y(n2148) );
  MX4X1 U7817 ( .A(n2097), .B(n2095), .C(n2096), .D(n2094), .S0(n4596), .S1(
        n4538), .Y(n2098) );
  MX4X1 U7818 ( .A(\registers[456][2] ), .B(\registers[457][2] ), .C(
        \registers[458][2] ), .D(\registers[459][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2095) );
  MX4X1 U7819 ( .A(\registers[460][2] ), .B(\registers[461][2] ), .C(
        \registers[462][2] ), .D(\registers[463][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2094) );
  MX4X1 U7820 ( .A(\registers[448][2] ), .B(\registers[449][2] ), .C(
        \registers[450][2] ), .D(\registers[451][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2097) );
  MX4X1 U7821 ( .A(n2082), .B(n2080), .C(n2081), .D(n2079), .S0(n4596), .S1(
        n4537), .Y(n2083) );
  MX4X1 U7822 ( .A(\registers[504][2] ), .B(\registers[505][2] ), .C(
        \registers[506][2] ), .D(\registers[507][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2080) );
  MX4X1 U7823 ( .A(\registers[508][2] ), .B(\registers[509][2] ), .C(
        \registers[510][2] ), .D(\registers[511][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2079) );
  MX4X1 U7824 ( .A(\registers[496][2] ), .B(\registers[497][2] ), .C(
        \registers[498][2] ), .D(\registers[499][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2082) );
  MX4X1 U7825 ( .A(n2119), .B(n2117), .C(n2118), .D(n2116), .S0(n4597), .S1(
        n4538), .Y(n2120) );
  MX4X1 U7826 ( .A(\registers[392][2] ), .B(\registers[393][2] ), .C(
        \registers[394][2] ), .D(\registers[395][2] ), .S0(n4160), .S1(n4397), 
        .Y(n2117) );
  MX4X1 U7827 ( .A(\registers[396][2] ), .B(\registers[397][2] ), .C(
        \registers[398][2] ), .D(\registers[399][2] ), .S0(n4160), .S1(n4397), 
        .Y(n2116) );
  MX4X1 U7828 ( .A(\registers[384][2] ), .B(\registers[385][2] ), .C(
        \registers[386][2] ), .D(\registers[387][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2119) );
  MX4X1 U7829 ( .A(n2103), .B(n2101), .C(n2102), .D(n2100), .S0(n4597), .S1(
        n4538), .Y(n2105) );
  MX4X1 U7830 ( .A(\registers[440][2] ), .B(\registers[441][2] ), .C(
        \registers[442][2] ), .D(\registers[443][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2101) );
  MX4X1 U7831 ( .A(\registers[444][2] ), .B(\registers[445][2] ), .C(
        \registers[446][2] ), .D(\registers[447][2] ), .S0(n4159), .S1(n4396), 
        .Y(n2100) );
  MX4X1 U7832 ( .A(\registers[432][2] ), .B(\registers[433][2] ), .C(
        \registers[434][2] ), .D(\registers[435][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2103) );
  MX4X1 U7833 ( .A(n2576), .B(n2574), .C(n2575), .D(n2573), .S0(n4603), .S1(
        n4542), .Y(n2577) );
  MX4X1 U7834 ( .A(\registers[264][3] ), .B(\registers[265][3] ), .C(
        \registers[266][3] ), .D(\registers[267][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2574) );
  MX4X1 U7835 ( .A(\registers[268][3] ), .B(\registers[269][3] ), .C(
        \registers[270][3] ), .D(\registers[271][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2573) );
  MX4X1 U7836 ( .A(\registers[256][3] ), .B(\registers[257][3] ), .C(
        \registers[258][3] ), .D(\registers[259][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2576) );
  MX4X1 U7837 ( .A(n2561), .B(n2559), .C(n2560), .D(n2558), .S0(n4603), .S1(
        n4543), .Y(n2562) );
  MX4X1 U7838 ( .A(\registers[312][3] ), .B(\registers[313][3] ), .C(
        \registers[314][3] ), .D(\registers[315][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2559) );
  MX4X1 U7839 ( .A(\registers[316][3] ), .B(\registers[317][3] ), .C(
        \registers[318][3] ), .D(\registers[319][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2558) );
  MX4X1 U7840 ( .A(\registers[304][3] ), .B(\registers[305][3] ), .C(
        \registers[306][3] ), .D(\registers[307][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2561) );
  MX4X1 U7841 ( .A(n2513), .B(n2511), .C(n2512), .D(n2510), .S0(n4602), .S1(
        n4543), .Y(n2514) );
  MX4X1 U7842 ( .A(\registers[456][3] ), .B(\registers[457][3] ), .C(
        \registers[458][3] ), .D(\registers[459][3] ), .S0(n4180), .S1(n4416), 
        .Y(n2511) );
  MX4X1 U7843 ( .A(\registers[460][3] ), .B(\registers[461][3] ), .C(
        \registers[462][3] ), .D(\registers[463][3] ), .S0(n4180), .S1(n4416), 
        .Y(n2510) );
  MX4X1 U7844 ( .A(\registers[448][3] ), .B(\registers[449][3] ), .C(
        \registers[450][3] ), .D(\registers[451][3] ), .S0(n4180), .S1(n4416), 
        .Y(n2513) );
  MX4X1 U7845 ( .A(n2498), .B(n2496), .C(n2497), .D(n2495), .S0(n4602), .S1(
        n4542), .Y(n2499) );
  MX4X1 U7846 ( .A(\registers[504][3] ), .B(\registers[505][3] ), .C(
        \registers[506][3] ), .D(\registers[507][3] ), .S0(n4179), .S1(n4415), 
        .Y(n2496) );
  MX4X1 U7847 ( .A(\registers[508][3] ), .B(\registers[509][3] ), .C(
        \registers[510][3] ), .D(\registers[511][3] ), .S0(n4179), .S1(n4415), 
        .Y(n2495) );
  MX4X1 U7848 ( .A(\registers[496][3] ), .B(\registers[497][3] ), .C(
        \registers[498][3] ), .D(\registers[499][3] ), .S0(n4179), .S1(n4415), 
        .Y(n2498) );
  MX4X1 U7849 ( .A(n2534), .B(n2532), .C(n2533), .D(n2531), .S0(n4602), .S1(
        n4543), .Y(n2535) );
  MX4X1 U7850 ( .A(\registers[392][3] ), .B(\registers[393][3] ), .C(
        \registers[394][3] ), .D(\registers[395][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2532) );
  MX4X1 U7851 ( .A(\registers[396][3] ), .B(\registers[397][3] ), .C(
        \registers[398][3] ), .D(\registers[399][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2531) );
  MX4X1 U7852 ( .A(\registers[384][3] ), .B(\registers[385][3] ), .C(
        \registers[386][3] ), .D(\registers[387][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2534) );
  MX4X1 U7853 ( .A(n2519), .B(n2517), .C(n2518), .D(n2516), .S0(n4602), .S1(
        n4543), .Y(n2520) );
  MX4X1 U7854 ( .A(\registers[440][3] ), .B(\registers[441][3] ), .C(
        \registers[442][3] ), .D(\registers[443][3] ), .S0(n4180), .S1(n4416), 
        .Y(n2517) );
  MX4X1 U7855 ( .A(\registers[444][3] ), .B(\registers[445][3] ), .C(
        \registers[446][3] ), .D(\registers[447][3] ), .S0(n4180), .S1(n4416), 
        .Y(n2516) );
  MX4X1 U7856 ( .A(\registers[432][3] ), .B(\registers[433][3] ), .C(
        \registers[434][3] ), .D(\registers[435][3] ), .S0(n4180), .S1(n4416), 
        .Y(n2519) );
  MX4X1 U7857 ( .A(n2916), .B(n2914), .C(n2915), .D(n2913), .S0(n4608), .S1(
        n4547), .Y(n2917) );
  MX4X1 U7858 ( .A(\registers[264][4] ), .B(\registers[265][4] ), .C(
        \registers[266][4] ), .D(\registers[267][4] ), .S0(n4205), .S1(n4439), 
        .Y(n2914) );
  MX4X1 U7859 ( .A(\registers[268][4] ), .B(\registers[269][4] ), .C(
        \registers[270][4] ), .D(\registers[271][4] ), .S0(n4205), .S1(n4439), 
        .Y(n2913) );
  MX4X1 U7860 ( .A(\registers[256][4] ), .B(\registers[257][4] ), .C(
        \registers[258][4] ), .D(\registers[259][4] ), .S0(n4205), .S1(n4439), 
        .Y(n2916) );
  MX4X1 U7861 ( .A(n2901), .B(n2899), .C(n2900), .D(n2898), .S0(n4608), .S1(
        n4547), .Y(n2902) );
  MX4X1 U7862 ( .A(\registers[312][4] ), .B(\registers[313][4] ), .C(
        \registers[314][4] ), .D(\registers[315][4] ), .S0(n4204), .S1(n4438), 
        .Y(n2899) );
  MX4X1 U7863 ( .A(\registers[316][4] ), .B(\registers[317][4] ), .C(
        \registers[318][4] ), .D(\registers[319][4] ), .S0(n4204), .S1(n4438), 
        .Y(n2898) );
  MX4X1 U7864 ( .A(\registers[304][4] ), .B(\registers[305][4] ), .C(
        \registers[306][4] ), .D(\registers[307][4] ), .S0(n4204), .S1(n4439), 
        .Y(n2901) );
  MX4X1 U7865 ( .A(n2853), .B(n2851), .C(n2852), .D(n2850), .S0(n4607), .S1(
        n4547), .Y(n2854) );
  MX4X1 U7866 ( .A(\registers[456][4] ), .B(\registers[457][4] ), .C(
        \registers[458][4] ), .D(\registers[459][4] ), .S0(n4201), .S1(n4436), 
        .Y(n2851) );
  MX4X1 U7867 ( .A(\registers[460][4] ), .B(\registers[461][4] ), .C(
        \registers[462][4] ), .D(\registers[463][4] ), .S0(n4201), .S1(n4436), 
        .Y(n2850) );
  MX4X1 U7868 ( .A(\registers[448][4] ), .B(\registers[449][4] ), .C(
        \registers[450][4] ), .D(\registers[451][4] ), .S0(n4201), .S1(n4436), 
        .Y(n2853) );
  MX4X1 U7869 ( .A(n2838), .B(n2836), .C(n2837), .D(n2835), .S0(n4607), .S1(
        n4546), .Y(n2839) );
  MX4X1 U7870 ( .A(\registers[504][4] ), .B(\registers[505][4] ), .C(
        \registers[506][4] ), .D(\registers[507][4] ), .S0(n4200), .S1(n4435), 
        .Y(n2836) );
  MX4X1 U7871 ( .A(\registers[508][4] ), .B(\registers[509][4] ), .C(
        \registers[510][4] ), .D(\registers[511][4] ), .S0(n4200), .S1(n4435), 
        .Y(n2835) );
  MX4X1 U7872 ( .A(\registers[496][4] ), .B(\registers[497][4] ), .C(
        \registers[498][4] ), .D(\registers[499][4] ), .S0(n4200), .S1(n4435), 
        .Y(n2838) );
  MX4X1 U7873 ( .A(n2874), .B(n2872), .C(n2873), .D(n2871), .S0(n4607), .S1(
        n4547), .Y(n2875) );
  MX4X1 U7874 ( .A(\registers[392][4] ), .B(\registers[393][4] ), .C(
        \registers[394][4] ), .D(\registers[395][4] ), .S0(n4202), .S1(n4437), 
        .Y(n2872) );
  MX4X1 U7875 ( .A(\registers[396][4] ), .B(\registers[397][4] ), .C(
        \registers[398][4] ), .D(\registers[399][4] ), .S0(n4202), .S1(n4437), 
        .Y(n2871) );
  MX4X1 U7876 ( .A(\registers[384][4] ), .B(\registers[385][4] ), .C(
        \registers[386][4] ), .D(\registers[387][4] ), .S0(n4202), .S1(n4437), 
        .Y(n2874) );
  MX4X1 U7877 ( .A(n2859), .B(n2857), .C(n2858), .D(n2856), .S0(n4607), .S1(
        n4547), .Y(n2860) );
  MX4X1 U7878 ( .A(\registers[440][4] ), .B(\registers[441][4] ), .C(
        \registers[442][4] ), .D(\registers[443][4] ), .S0(n4201), .S1(n4436), 
        .Y(n2857) );
  MX4X1 U7879 ( .A(\registers[444][4] ), .B(\registers[445][4] ), .C(
        \registers[446][4] ), .D(\registers[447][4] ), .S0(n4201), .S1(n4436), 
        .Y(n2856) );
  MX4X1 U7880 ( .A(\registers[432][4] ), .B(\registers[433][4] ), .C(
        \registers[434][4] ), .D(\registers[435][4] ), .S0(n4201), .S1(n4436), 
        .Y(n2859) );
  MX4X1 U7881 ( .A(n3241), .B(n3239), .C(n3240), .D(n3238), .S0(n4613), .S1(
        n4552), .Y(n3242) );
  MX4X1 U7882 ( .A(\registers[312][5] ), .B(\registers[313][5] ), .C(
        \registers[314][5] ), .D(\registers[315][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3239) );
  MX4X1 U7883 ( .A(\registers[316][5] ), .B(\registers[317][5] ), .C(
        \registers[318][5] ), .D(\registers[319][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3238) );
  MX4X1 U7884 ( .A(\registers[304][5] ), .B(\registers[305][5] ), .C(
        \registers[306][5] ), .D(\registers[307][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3241) );
  MX4X1 U7885 ( .A(n3178), .B(n3176), .C(n3177), .D(n3175), .S0(n4612), .S1(
        n4551), .Y(n3179) );
  MX4X1 U7886 ( .A(\registers[504][5] ), .B(\registers[505][5] ), .C(
        \registers[506][5] ), .D(\registers[507][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3176) );
  MX4X1 U7887 ( .A(\registers[508][5] ), .B(\registers[509][5] ), .C(
        \registers[510][5] ), .D(\registers[511][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3175) );
  MX4X1 U7888 ( .A(\registers[496][5] ), .B(\registers[497][5] ), .C(
        \registers[498][5] ), .D(\registers[499][5] ), .S0(n4221), .S1(n4455), 
        .Y(n3178) );
  MX4X1 U7889 ( .A(n3199), .B(n3197), .C(n3198), .D(n3196), .S0(n4613), .S1(
        n4552), .Y(n3200) );
  MX4X1 U7890 ( .A(\registers[440][5] ), .B(\registers[441][5] ), .C(
        \registers[442][5] ), .D(\registers[443][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3197) );
  MX4X1 U7891 ( .A(\registers[444][5] ), .B(\registers[445][5] ), .C(
        \registers[446][5] ), .D(\registers[447][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3196) );
  MX4X1 U7892 ( .A(\registers[432][5] ), .B(\registers[433][5] ), .C(
        \registers[434][5] ), .D(\registers[435][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3199) );
  MX4X1 U7893 ( .A(n3581), .B(n3579), .C(n3580), .D(n3578), .S0(n4619), .S1(
        n4557), .Y(n3582) );
  MX4X1 U7894 ( .A(\registers[312][6] ), .B(\registers[313][6] ), .C(
        \registers[314][6] ), .D(\registers[315][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3579) );
  MX4X1 U7895 ( .A(\registers[316][6] ), .B(\registers[317][6] ), .C(
        \registers[318][6] ), .D(\registers[319][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3578) );
  MX4X1 U7896 ( .A(\registers[304][6] ), .B(\registers[305][6] ), .C(
        \registers[306][6] ), .D(\registers[307][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3581) );
  MX4X1 U7897 ( .A(n3518), .B(n3516), .C(n3517), .D(n3515), .S0(n4618), .S1(
        n4556), .Y(n3519) );
  MX4X1 U7898 ( .A(\registers[504][6] ), .B(\registers[505][6] ), .C(
        \registers[506][6] ), .D(\registers[507][6] ), .S0(n4243), .S1(n4474), 
        .Y(n3516) );
  MX4X1 U7899 ( .A(\registers[508][6] ), .B(\registers[509][6] ), .C(
        \registers[510][6] ), .D(\registers[511][6] ), .S0(n4243), .S1(n4474), 
        .Y(n3515) );
  MX4X1 U7900 ( .A(\registers[496][6] ), .B(\registers[497][6] ), .C(
        \registers[498][6] ), .D(\registers[499][6] ), .S0(n4243), .S1(n4474), 
        .Y(n3518) );
  MX4X1 U7901 ( .A(n3539), .B(n3537), .C(n3538), .D(n3536), .S0(n4618), .S1(
        n4556), .Y(n3540) );
  MX4X1 U7902 ( .A(\registers[440][6] ), .B(\registers[441][6] ), .C(
        \registers[442][6] ), .D(\registers[443][6] ), .S0(n4244), .S1(n4475), 
        .Y(n3537) );
  MX4X1 U7903 ( .A(\registers[444][6] ), .B(\registers[445][6] ), .C(
        \registers[446][6] ), .D(\registers[447][6] ), .S0(n4244), .S1(n4475), 
        .Y(n3536) );
  MX4X1 U7904 ( .A(\registers[432][6] ), .B(\registers[433][6] ), .C(
        \registers[434][6] ), .D(\registers[435][6] ), .S0(n4244), .S1(n4475), 
        .Y(n3539) );
  MX4X1 U7905 ( .A(n3921), .B(n3919), .C(n3920), .D(n3918), .S0(n4624), .S1(
        n4558), .Y(n3922) );
  MX4X1 U7906 ( .A(\registers[312][7] ), .B(\registers[313][7] ), .C(
        \registers[314][7] ), .D(\registers[315][7] ), .S0(n4268), .S1(n4470), 
        .Y(n3919) );
  MX4X1 U7907 ( .A(\registers[316][7] ), .B(\registers[317][7] ), .C(
        \registers[318][7] ), .D(\registers[319][7] ), .S0(n4268), .S1(n4482), 
        .Y(n3918) );
  MX4X1 U7908 ( .A(\registers[304][7] ), .B(\registers[305][7] ), .C(
        \registers[306][7] ), .D(\registers[307][7] ), .S0(n4268), .S1(n4497), 
        .Y(n3921) );
  MX4X1 U7909 ( .A(n3858), .B(n3856), .C(n3857), .D(n3855), .S0(n4623), .S1(
        n4559), .Y(n3859) );
  MX4X1 U7910 ( .A(\registers[504][7] ), .B(\registers[505][7] ), .C(
        \registers[506][7] ), .D(\registers[507][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3856) );
  MX4X1 U7911 ( .A(\registers[508][7] ), .B(\registers[509][7] ), .C(
        \registers[510][7] ), .D(\registers[511][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3855) );
  MX4X1 U7912 ( .A(\registers[496][7] ), .B(\registers[497][7] ), .C(
        \registers[498][7] ), .D(\registers[499][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3858) );
  MX4X1 U7913 ( .A(n3879), .B(n3877), .C(n3878), .D(n3876), .S0(n4623), .S1(
        n4543), .Y(n3880) );
  MX4X1 U7914 ( .A(\registers[440][7] ), .B(\registers[441][7] ), .C(
        \registers[442][7] ), .D(\registers[443][7] ), .S0(n4265), .S1(n4495), 
        .Y(n3877) );
  MX4X1 U7915 ( .A(\registers[444][7] ), .B(\registers[445][7] ), .C(
        \registers[446][7] ), .D(\registers[447][7] ), .S0(n4265), .S1(n4495), 
        .Y(n3876) );
  MX4X1 U7916 ( .A(\registers[432][7] ), .B(\registers[433][7] ), .C(
        \registers[434][7] ), .D(\registers[435][7] ), .S0(n4265), .S1(n4495), 
        .Y(n3879) );
  MX4X1 U7917 ( .A(n4886), .B(n4884), .C(n4885), .D(n4883), .S0(n7930), .S1(
        n7870), .Y(n4887) );
  MX4X1 U7918 ( .A(\registers[312][0] ), .B(\registers[313][0] ), .C(
        \registers[314][0] ), .D(\registers[315][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4884) );
  MX4X1 U7919 ( .A(\registers[316][0] ), .B(\registers[317][0] ), .C(
        \registers[318][0] ), .D(\registers[319][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4883) );
  MX4X1 U7920 ( .A(\registers[304][0] ), .B(\registers[305][0] ), .C(
        \registers[306][0] ), .D(\registers[307][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4886) );
  MX4X1 U7921 ( .A(n4823), .B(n4821), .C(n4822), .D(n4820), .S0(n7942), .S1(
        n7869), .Y(n4824) );
  MX4X1 U7922 ( .A(\registers[504][0] ), .B(\registers[505][0] ), .C(
        \registers[506][0] ), .D(\registers[507][0] ), .S0(n7458), .S1(n7700), 
        .Y(n4821) );
  MX4X1 U7923 ( .A(\registers[508][0] ), .B(\registers[509][0] ), .C(
        \registers[510][0] ), .D(\registers[511][0] ), .S0(n7458), .S1(n7700), 
        .Y(n4820) );
  MX4X1 U7924 ( .A(\registers[496][0] ), .B(\registers[497][0] ), .C(
        \registers[498][0] ), .D(\registers[499][0] ), .S0(n7458), .S1(n7700), 
        .Y(n4823) );
  MX4X1 U7925 ( .A(n4844), .B(n4842), .C(n4843), .D(n4841), .S0(n7937), .S1(
        n7869), .Y(n4845) );
  MX4X1 U7926 ( .A(\registers[440][0] ), .B(\registers[441][0] ), .C(
        \registers[442][0] ), .D(\registers[443][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4842) );
  MX4X1 U7927 ( .A(\registers[444][0] ), .B(\registers[445][0] ), .C(
        \registers[446][0] ), .D(\registers[447][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4841) );
  MX4X1 U7928 ( .A(\registers[432][0] ), .B(\registers[433][0] ), .C(
        \registers[434][0] ), .D(\registers[435][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4844) );
  MX4X1 U7929 ( .A(n5226), .B(n5224), .C(n5225), .D(n5223), .S0(n7935), .S1(
        n7874), .Y(n5227) );
  MX4X1 U7930 ( .A(\registers[312][1] ), .B(\registers[313][1] ), .C(
        \registers[314][1] ), .D(\registers[315][1] ), .S0(n7483), .S1(n7723), 
        .Y(n5224) );
  MX4X1 U7931 ( .A(\registers[316][1] ), .B(\registers[317][1] ), .C(
        \registers[318][1] ), .D(\registers[319][1] ), .S0(n7483), .S1(n7723), 
        .Y(n5223) );
  MX4X1 U7932 ( .A(\registers[304][1] ), .B(\registers[305][1] ), .C(
        \registers[306][1] ), .D(\registers[307][1] ), .S0(n7483), .S1(n7723), 
        .Y(n5226) );
  MX4X1 U7933 ( .A(n5163), .B(n5161), .C(n5162), .D(n5160), .S0(n7934), .S1(
        n7874), .Y(n5164) );
  MX4X1 U7934 ( .A(\registers[504][1] ), .B(\registers[505][1] ), .C(
        \registers[506][1] ), .D(\registers[507][1] ), .S0(n7479), .S1(n7720), 
        .Y(n5161) );
  MX4X1 U7935 ( .A(\registers[508][1] ), .B(\registers[509][1] ), .C(
        \registers[510][1] ), .D(\registers[511][1] ), .S0(n7479), .S1(n7720), 
        .Y(n5160) );
  MX4X1 U7936 ( .A(\registers[496][1] ), .B(\registers[497][1] ), .C(
        \registers[498][1] ), .D(\registers[499][1] ), .S0(n7479), .S1(n7720), 
        .Y(n5163) );
  MX4X1 U7937 ( .A(n5184), .B(n5182), .C(n5183), .D(n5181), .S0(n7934), .S1(
        n7874), .Y(n5185) );
  MX4X1 U7938 ( .A(\registers[440][1] ), .B(\registers[441][1] ), .C(
        \registers[442][1] ), .D(\registers[443][1] ), .S0(n7480), .S1(n7721), 
        .Y(n5182) );
  MX4X1 U7939 ( .A(\registers[444][1] ), .B(\registers[445][1] ), .C(
        \registers[446][1] ), .D(\registers[447][1] ), .S0(n7480), .S1(n7721), 
        .Y(n5181) );
  MX4X1 U7940 ( .A(\registers[432][1] ), .B(\registers[433][1] ), .C(
        \registers[434][1] ), .D(\registers[435][1] ), .S0(n7480), .S1(n7721), 
        .Y(n5184) );
  MX4X1 U7941 ( .A(n5566), .B(n5564), .C(n5565), .D(n5563), .S0(n7940), .S1(
        n7879), .Y(n5567) );
  MX4X1 U7942 ( .A(\registers[312][2] ), .B(\registers[313][2] ), .C(
        \registers[314][2] ), .D(\registers[315][2] ), .S0(n7504), .S1(n7743), 
        .Y(n5564) );
  MX4X1 U7943 ( .A(\registers[316][2] ), .B(\registers[317][2] ), .C(
        \registers[318][2] ), .D(\registers[319][2] ), .S0(n7504), .S1(n7743), 
        .Y(n5563) );
  MX4X1 U7944 ( .A(\registers[304][2] ), .B(\registers[305][2] ), .C(
        \registers[306][2] ), .D(\registers[307][2] ), .S0(n7504), .S1(n7743), 
        .Y(n5566) );
  MX4X1 U7945 ( .A(n5503), .B(n5501), .C(n5502), .D(n5500), .S0(n7939), .S1(
        n7878), .Y(n5504) );
  MX4X1 U7946 ( .A(\registers[504][2] ), .B(\registers[505][2] ), .C(
        \registers[506][2] ), .D(\registers[507][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5501) );
  MX4X1 U7947 ( .A(\registers[508][2] ), .B(\registers[509][2] ), .C(
        \registers[510][2] ), .D(\registers[511][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5500) );
  MX4X1 U7948 ( .A(\registers[496][2] ), .B(\registers[497][2] ), .C(
        \registers[498][2] ), .D(\registers[499][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5503) );
  MX4X1 U7949 ( .A(n5524), .B(n5522), .C(n5523), .D(n5521), .S0(n7940), .S1(
        n7879), .Y(n5525) );
  MX4X1 U7950 ( .A(\registers[440][2] ), .B(\registers[441][2] ), .C(
        \registers[442][2] ), .D(\registers[443][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5522) );
  MX4X1 U7951 ( .A(\registers[444][2] ), .B(\registers[445][2] ), .C(
        \registers[446][2] ), .D(\registers[447][2] ), .S0(n7502), .S1(n7740), 
        .Y(n5521) );
  MX4X1 U7952 ( .A(\registers[432][2] ), .B(\registers[433][2] ), .C(
        \registers[434][2] ), .D(\registers[435][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5524) );
  MX4X1 U7953 ( .A(n5906), .B(n5904), .C(n5905), .D(n5903), .S0(n7946), .S1(
        n7884), .Y(n5907) );
  MX4X1 U7954 ( .A(\registers[312][3] ), .B(\registers[313][3] ), .C(
        \registers[314][3] ), .D(\registers[315][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5904) );
  MX4X1 U7955 ( .A(\registers[316][3] ), .B(\registers[317][3] ), .C(
        \registers[318][3] ), .D(\registers[319][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5903) );
  MX4X1 U7956 ( .A(\registers[304][3] ), .B(\registers[305][3] ), .C(
        \registers[306][3] ), .D(\registers[307][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5906) );
  MX4X1 U7957 ( .A(n5843), .B(n5841), .C(n5842), .D(n5840), .S0(n7945), .S1(
        n7883), .Y(n5844) );
  MX4X1 U7958 ( .A(\registers[504][3] ), .B(\registers[505][3] ), .C(
        \registers[506][3] ), .D(\registers[507][3] ), .S0(n7522), .S1(n7759), 
        .Y(n5841) );
  MX4X1 U7959 ( .A(\registers[508][3] ), .B(\registers[509][3] ), .C(
        \registers[510][3] ), .D(\registers[511][3] ), .S0(n7522), .S1(n7759), 
        .Y(n5840) );
  MX4X1 U7960 ( .A(\registers[496][3] ), .B(\registers[497][3] ), .C(
        \registers[498][3] ), .D(\registers[499][3] ), .S0(n7522), .S1(n7759), 
        .Y(n5843) );
  MX4X1 U7961 ( .A(n5864), .B(n5862), .C(n5863), .D(n5861), .S0(n7945), .S1(
        n7884), .Y(n5865) );
  MX4X1 U7962 ( .A(\registers[440][3] ), .B(\registers[441][3] ), .C(
        \registers[442][3] ), .D(\registers[443][3] ), .S0(n7523), .S1(n7760), 
        .Y(n5862) );
  MX4X1 U7963 ( .A(\registers[444][3] ), .B(\registers[445][3] ), .C(
        \registers[446][3] ), .D(\registers[447][3] ), .S0(n7523), .S1(n7760), 
        .Y(n5861) );
  MX4X1 U7964 ( .A(\registers[432][3] ), .B(\registers[433][3] ), .C(
        \registers[434][3] ), .D(\registers[435][3] ), .S0(n7523), .S1(n7760), 
        .Y(n5864) );
  MX4X1 U7965 ( .A(n6246), .B(n6244), .C(n6245), .D(n6243), .S0(n7951), .S1(
        n7889), .Y(n6247) );
  MX4X1 U7966 ( .A(\registers[312][4] ), .B(\registers[313][4] ), .C(
        \registers[314][4] ), .D(\registers[315][4] ), .S0(n7547), .S1(n7782), 
        .Y(n6244) );
  MX4X1 U7967 ( .A(\registers[316][4] ), .B(\registers[317][4] ), .C(
        \registers[318][4] ), .D(\registers[319][4] ), .S0(n7547), .S1(n7782), 
        .Y(n6243) );
  MX4X1 U7968 ( .A(\registers[304][4] ), .B(\registers[305][4] ), .C(
        \registers[306][4] ), .D(\registers[307][4] ), .S0(n7547), .S1(n7783), 
        .Y(n6246) );
  MX4X1 U7969 ( .A(n6183), .B(n6181), .C(n6182), .D(n6180), .S0(n7950), .S1(
        n7888), .Y(n6184) );
  MX4X1 U7970 ( .A(\registers[504][4] ), .B(\registers[505][4] ), .C(
        \registers[506][4] ), .D(\registers[507][4] ), .S0(n7543), .S1(n7779), 
        .Y(n6181) );
  MX4X1 U7971 ( .A(\registers[508][4] ), .B(\registers[509][4] ), .C(
        \registers[510][4] ), .D(\registers[511][4] ), .S0(n7543), .S1(n7779), 
        .Y(n6180) );
  MX4X1 U7972 ( .A(\registers[496][4] ), .B(\registers[497][4] ), .C(
        \registers[498][4] ), .D(\registers[499][4] ), .S0(n7543), .S1(n7779), 
        .Y(n6183) );
  MX4X1 U7973 ( .A(n6204), .B(n6202), .C(n6203), .D(n6201), .S0(n7950), .S1(
        n7889), .Y(n6205) );
  MX4X1 U7974 ( .A(\registers[440][4] ), .B(\registers[441][4] ), .C(
        \registers[442][4] ), .D(\registers[443][4] ), .S0(n7544), .S1(n7780), 
        .Y(n6202) );
  MX4X1 U7975 ( .A(\registers[444][4] ), .B(\registers[445][4] ), .C(
        \registers[446][4] ), .D(\registers[447][4] ), .S0(n7544), .S1(n7780), 
        .Y(n6201) );
  MX4X1 U7976 ( .A(\registers[432][4] ), .B(\registers[433][4] ), .C(
        \registers[434][4] ), .D(\registers[435][4] ), .S0(n7544), .S1(n7780), 
        .Y(n6204) );
  MX4X1 U7977 ( .A(n6586), .B(n6584), .C(n6585), .D(n6583), .S0(n7956), .S1(
        n7894), .Y(n6587) );
  MX4X1 U7978 ( .A(\registers[312][5] ), .B(\registers[313][5] ), .C(
        \registers[314][5] ), .D(\registers[315][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6584) );
  MX4X1 U7979 ( .A(\registers[316][5] ), .B(\registers[317][5] ), .C(
        \registers[318][5] ), .D(\registers[319][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6583) );
  MX4X1 U7980 ( .A(\registers[304][5] ), .B(\registers[305][5] ), .C(
        \registers[306][5] ), .D(\registers[307][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6586) );
  MX4X1 U7981 ( .A(n6523), .B(n6521), .C(n6522), .D(n6520), .S0(n7955), .S1(
        n7893), .Y(n6524) );
  MX4X1 U7982 ( .A(\registers[504][5] ), .B(\registers[505][5] ), .C(
        \registers[506][5] ), .D(\registers[507][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6521) );
  MX4X1 U7983 ( .A(\registers[508][5] ), .B(\registers[509][5] ), .C(
        \registers[510][5] ), .D(\registers[511][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6520) );
  MX4X1 U7984 ( .A(\registers[496][5] ), .B(\registers[497][5] ), .C(
        \registers[498][5] ), .D(\registers[499][5] ), .S0(n7564), .S1(n7799), 
        .Y(n6523) );
  MX4X1 U7985 ( .A(n6544), .B(n6542), .C(n6543), .D(n6541), .S0(n7956), .S1(
        n7894), .Y(n6545) );
  MX4X1 U7986 ( .A(\registers[440][5] ), .B(\registers[441][5] ), .C(
        \registers[442][5] ), .D(\registers[443][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6542) );
  MX4X1 U7987 ( .A(\registers[444][5] ), .B(\registers[445][5] ), .C(
        \registers[446][5] ), .D(\registers[447][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6541) );
  MX4X1 U7988 ( .A(\registers[432][5] ), .B(\registers[433][5] ), .C(
        \registers[434][5] ), .D(\registers[435][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6544) );
  MX4X1 U7989 ( .A(n6926), .B(n6924), .C(n6925), .D(n6923), .S0(n7962), .S1(
        n7897), .Y(n6927) );
  MX4X1 U7990 ( .A(\registers[312][6] ), .B(\registers[313][6] ), .C(
        \registers[314][6] ), .D(\registers[315][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6924) );
  MX4X1 U7991 ( .A(\registers[316][6] ), .B(\registers[317][6] ), .C(
        \registers[318][6] ), .D(\registers[319][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6923) );
  MX4X1 U7992 ( .A(\registers[304][6] ), .B(\registers[305][6] ), .C(
        \registers[306][6] ), .D(\registers[307][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6926) );
  MX4X1 U7993 ( .A(n6863), .B(n6861), .C(n6862), .D(n6860), .S0(n7961), .S1(
        n7891), .Y(n6864) );
  MX4X1 U7994 ( .A(\registers[504][6] ), .B(\registers[505][6] ), .C(
        \registers[506][6] ), .D(\registers[507][6] ), .S0(n7586), .S1(n7817), 
        .Y(n6861) );
  MX4X1 U7995 ( .A(\registers[508][6] ), .B(\registers[509][6] ), .C(
        \registers[510][6] ), .D(\registers[511][6] ), .S0(n7586), .S1(n7817), 
        .Y(n6860) );
  MX4X1 U7996 ( .A(\registers[496][6] ), .B(\registers[497][6] ), .C(
        \registers[498][6] ), .D(\registers[499][6] ), .S0(n7586), .S1(n7817), 
        .Y(n6863) );
  MX4X1 U7997 ( .A(n6884), .B(n6882), .C(n6883), .D(n6881), .S0(n7961), .S1(
        n7890), .Y(n6885) );
  MX4X1 U7998 ( .A(\registers[440][6] ), .B(\registers[441][6] ), .C(
        \registers[442][6] ), .D(\registers[443][6] ), .S0(n7587), .S1(n7818), 
        .Y(n6882) );
  MX4X1 U7999 ( .A(\registers[444][6] ), .B(\registers[445][6] ), .C(
        \registers[446][6] ), .D(\registers[447][6] ), .S0(n7587), .S1(n7818), 
        .Y(n6881) );
  MX4X1 U8000 ( .A(\registers[432][6] ), .B(\registers[433][6] ), .C(
        \registers[434][6] ), .D(\registers[435][6] ), .S0(n7587), .S1(n7818), 
        .Y(n6884) );
  MX4X1 U8001 ( .A(n7203), .B(n7201), .C(n7202), .D(n7200), .S0(n7966), .S1(
        n7901), .Y(n7204) );
  MX4X1 U8002 ( .A(\registers[504][7] ), .B(\registers[505][7] ), .C(
        \registers[506][7] ), .D(\registers[507][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7201) );
  MX4X1 U8003 ( .A(\registers[508][7] ), .B(\registers[509][7] ), .C(
        \registers[510][7] ), .D(\registers[511][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7200) );
  MX4X1 U8004 ( .A(\registers[496][7] ), .B(\registers[497][7] ), .C(
        \registers[498][7] ), .D(\registers[499][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7203) );
  MX4X1 U8005 ( .A(n7224), .B(n7222), .C(n7223), .D(n7221), .S0(n7966), .S1(
        n7901), .Y(n7225) );
  MX4X1 U8006 ( .A(\registers[440][7] ), .B(\registers[441][7] ), .C(
        \registers[442][7] ), .D(\registers[443][7] ), .S0(n7608), .S1(n7838), 
        .Y(n7222) );
  MX4X1 U8007 ( .A(\registers[444][7] ), .B(\registers[445][7] ), .C(
        \registers[446][7] ), .D(\registers[447][7] ), .S0(n7608), .S1(n7838), 
        .Y(n7221) );
  MX4X1 U8008 ( .A(\registers[432][7] ), .B(\registers[433][7] ), .C(
        \registers[434][7] ), .D(\registers[435][7] ), .S0(n7608), .S1(n7838), 
        .Y(n7224) );
  MX4X1 U8009 ( .A(n7266), .B(n7264), .C(n7265), .D(n7263), .S0(n7967), .S1(
        n7901), .Y(n7267) );
  MX4X1 U8010 ( .A(\registers[312][7] ), .B(\registers[313][7] ), .C(
        \registers[314][7] ), .D(\registers[315][7] ), .S0(n7611), .S1(n7840), 
        .Y(n7264) );
  MX4X1 U8011 ( .A(\registers[316][7] ), .B(\registers[317][7] ), .C(
        \registers[318][7] ), .D(\registers[319][7] ), .S0(n7611), .S1(n7840), 
        .Y(n7263) );
  MX4X1 U8012 ( .A(\registers[304][7] ), .B(\registers[305][7] ), .C(
        \registers[306][7] ), .D(\registers[307][7] ), .S0(n7611), .S1(n7841), 
        .Y(n7266) );
  MX4X1 U8013 ( .A(n1079), .B(n1077), .C(n1078), .D(n1076), .S0(n4624), .S1(
        n4526), .Y(n1080) );
  MX4X1 U8014 ( .A(\registers[920][0] ), .B(\registers[921][0] ), .C(
        \registers[922][0] ), .D(\registers[923][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1077) );
  MX4X1 U8015 ( .A(\registers[924][0] ), .B(\registers[925][0] ), .C(
        \registers[926][0] ), .D(\registers[927][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1076) );
  MX4X1 U8016 ( .A(\registers[912][0] ), .B(\registers[913][0] ), .C(
        \registers[914][0] ), .D(\registers[915][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1079) );
  MX4X1 U8017 ( .A(n4684), .B(n4682), .C(n4683), .D(n4681), .S0(n7967), .S1(
        n7867), .Y(n4685) );
  MX4X1 U8018 ( .A(\registers[920][0] ), .B(\registers[921][0] ), .C(
        \registers[922][0] ), .D(\registers[923][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4682) );
  MX4X1 U8019 ( .A(\registers[924][0] ), .B(\registers[925][0] ), .C(
        \registers[926][0] ), .D(\registers[927][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4681) );
  MX4X1 U8020 ( .A(\registers[912][0] ), .B(\registers[913][0] ), .C(
        \registers[914][0] ), .D(\registers[915][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4684) );
  MX4X1 U8021 ( .A(n1058), .B(n1056), .C(n1057), .D(n1055), .S0(n4624), .S1(
        n4525), .Y(n1059) );
  MX4X1 U8022 ( .A(\registers[984][0] ), .B(\registers[985][0] ), .C(
        \registers[986][0] ), .D(\registers[987][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1056) );
  MX4X1 U8023 ( .A(\registers[988][0] ), .B(\registers[989][0] ), .C(
        \registers[990][0] ), .D(\registers[991][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1055) );
  MX4X1 U8024 ( .A(\registers[976][0] ), .B(\registers[977][0] ), .C(
        \registers[978][0] ), .D(\registers[979][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1058) );
  MX4X1 U8025 ( .A(n4663), .B(n4661), .C(n4662), .D(n4660), .S0(n7967), .S1(
        n7866), .Y(n4664) );
  MX4X1 U8026 ( .A(\registers[984][0] ), .B(\registers[985][0] ), .C(
        \registers[986][0] ), .D(\registers[987][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4661) );
  MX4X1 U8027 ( .A(\registers[988][0] ), .B(\registers[989][0] ), .C(
        \registers[990][0] ), .D(\registers[991][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4660) );
  MX4X1 U8028 ( .A(\registers[976][0] ), .B(\registers[977][0] ), .C(
        \registers[978][0] ), .D(\registers[979][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4663) );
  MX4X1 U8029 ( .A(\registers[1016][0] ), .B(\registers[1017][0] ), .C(
        \registers[1018][0] ), .D(\registers[1019][0] ), .S0(n4252), .S1(n4350), .Y(n1046) );
  MX4X1 U8030 ( .A(\registers[1000][0] ), .B(\registers[1001][0] ), .C(
        \registers[1002][0] ), .D(\registers[1003][0] ), .S0(n4106), .S1(n4471), .Y(n1051) );
  MX4X1 U8031 ( .A(\registers[1016][0] ), .B(\registers[1017][0] ), .C(
        \registers[1018][0] ), .D(\registers[1019][0] ), .S0(n7576), .S1(n7700), .Y(n4651) );
  MX4X1 U8032 ( .A(\registers[1000][0] ), .B(\registers[1001][0] ), .C(
        \registers[1002][0] ), .D(\registers[1003][0] ), .S0(n7608), .S1(n7809), .Y(n4656) );
  MX4X1 U8033 ( .A(\registers[328][0] ), .B(\registers[329][0] ), .C(
        \registers[330][0] ), .D(\registers[331][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1429) );
  MX4X1 U8034 ( .A(\registers[376][0] ), .B(\registers[377][0] ), .C(
        \registers[378][0] ), .D(\registers[379][0] ), .S0(n4117), .S1(n4358), 
        .Y(n1414) );
  MX4X1 U8035 ( .A(\registers[360][0] ), .B(\registers[361][0] ), .C(
        \registers[362][0] ), .D(\registers[363][0] ), .S0(n4118), .S1(n4359), 
        .Y(n1419) );
  MX4X1 U8036 ( .A(\registers[72][0] ), .B(\registers[73][0] ), .C(
        \registers[74][0] ), .D(\registers[75][0] ), .S0(n4124), .S1(n4364), 
        .Y(n1520) );
  MX4X1 U8037 ( .A(\registers[120][0] ), .B(\registers[121][0] ), .C(
        \registers[122][0] ), .D(\registers[123][0] ), .S0(n4123), .S1(n4363), 
        .Y(n1504) );
  MX4X1 U8038 ( .A(\registers[104][0] ), .B(\registers[105][0] ), .C(
        \registers[106][0] ), .D(\registers[107][0] ), .S0(n4123), .S1(n4364), 
        .Y(n1510) );
  MX4X1 U8039 ( .A(\registers[8][0] ), .B(\registers[9][0] ), .C(
        \registers[10][0] ), .D(\registers[11][0] ), .S0(n4125), .S1(n4365), 
        .Y(n1543) );
  MX4X1 U8040 ( .A(\registers[56][0] ), .B(\registers[57][0] ), .C(
        \registers[58][0] ), .D(\registers[59][0] ), .S0(n4124), .S1(n4365), 
        .Y(n1526) );
  MX4X1 U8041 ( .A(\registers[40][0] ), .B(\registers[41][0] ), .C(
        \registers[42][0] ), .D(\registers[43][0] ), .S0(n4124), .S1(n4365), 
        .Y(n1531) );
  MX4X1 U8042 ( .A(\registers[200][0] ), .B(\registers[201][0] ), .C(
        \registers[202][0] ), .D(\registers[203][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1476) );
  MX4X1 U8043 ( .A(\registers[248][0] ), .B(\registers[249][0] ), .C(
        \registers[250][0] ), .D(\registers[251][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1459) );
  MX4X1 U8044 ( .A(\registers[232][0] ), .B(\registers[233][0] ), .C(
        \registers[234][0] ), .D(\registers[235][0] ), .S0(n4120), .S1(n4361), 
        .Y(n1464) );
  MX4X1 U8045 ( .A(\registers[136][0] ), .B(\registers[137][0] ), .C(
        \registers[138][0] ), .D(\registers[139][0] ), .S0(n4122), .S1(n4363), 
        .Y(n1497) );
  MX4X1 U8046 ( .A(\registers[184][0] ), .B(\registers[185][0] ), .C(
        \registers[186][0] ), .D(\registers[187][0] ), .S0(n4121), .S1(n4362), 
        .Y(n1482) );
  MX4X1 U8047 ( .A(\registers[168][0] ), .B(\registers[169][0] ), .C(
        \registers[170][0] ), .D(\registers[171][0] ), .S0(n4122), .S1(n4362), 
        .Y(n1487) );
  MX4X1 U8048 ( .A(\registers[840][0] ), .B(\registers[841][0] ), .C(
        \registers[842][0] ), .D(\registers[843][0] ), .S0(n4108), .S1(n4487), 
        .Y(n1103) );
  MX4X1 U8049 ( .A(\registers[888][0] ), .B(\registers[889][0] ), .C(
        \registers[890][0] ), .D(\registers[891][0] ), .S0(n4107), .S1(n4491), 
        .Y(n1088) );
  MX4X1 U8050 ( .A(\registers[872][0] ), .B(\registers[873][0] ), .C(
        \registers[874][0] ), .D(\registers[875][0] ), .S0(n4107), .S1(n4475), 
        .Y(n1093) );
  MX4X1 U8051 ( .A(\registers[776][0] ), .B(\registers[777][0] ), .C(
        \registers[778][0] ), .D(\registers[779][0] ), .S0(n4109), .S1(n4351), 
        .Y(n1166) );
  MX4X1 U8052 ( .A(\registers[824][0] ), .B(\registers[825][0] ), .C(
        \registers[826][0] ), .D(\registers[827][0] ), .S0(n4108), .S1(n4484), 
        .Y(n1151) );
  MX4X1 U8053 ( .A(\registers[808][0] ), .B(\registers[809][0] ), .C(
        \registers[810][0] ), .D(\registers[811][0] ), .S0(n4108), .S1(n4378), 
        .Y(n1156) );
  MX4X1 U8054 ( .A(\registers[968][0] ), .B(\registers[969][0] ), .C(
        \registers[970][0] ), .D(\registers[971][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1061) );
  MX4X1 U8055 ( .A(\registers[904][0] ), .B(\registers[905][0] ), .C(
        \registers[906][0] ), .D(\registers[907][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1082) );
  MX4X1 U8056 ( .A(\registers[952][0] ), .B(\registers[953][0] ), .C(
        \registers[954][0] ), .D(\registers[955][0] ), .S0(n4105), .S1(n4349), 
        .Y(n1067) );
  MX4X1 U8057 ( .A(\registers[936][0] ), .B(\registers[937][0] ), .C(
        \registers[938][0] ), .D(\registers[939][0] ), .S0(n4106), .S1(n4350), 
        .Y(n1072) );
  MX4X1 U8058 ( .A(\registers[584][0] ), .B(\registers[585][0] ), .C(
        \registers[586][0] ), .D(\registers[587][0] ), .S0(n4113), .S1(n4354), 
        .Y(n1339) );
  MX4X1 U8059 ( .A(\registers[632][0] ), .B(\registers[633][0] ), .C(
        \registers[634][0] ), .D(\registers[635][0] ), .S0(n4112), .S1(n4353), 
        .Y(n1313) );
  MX4X1 U8060 ( .A(\registers[616][0] ), .B(\registers[617][0] ), .C(
        \registers[618][0] ), .D(\registers[619][0] ), .S0(n4112), .S1(n4354), 
        .Y(n1323) );
  MX4X1 U8061 ( .A(\registers[520][0] ), .B(\registers[521][0] ), .C(
        \registers[522][0] ), .D(\registers[523][0] ), .S0(n4114), .S1(n4356), 
        .Y(n1360) );
  MX4X1 U8062 ( .A(\registers[568][0] ), .B(\registers[569][0] ), .C(
        \registers[570][0] ), .D(\registers[571][0] ), .S0(n4113), .S1(n4355), 
        .Y(n1345) );
  MX4X1 U8063 ( .A(\registers[552][0] ), .B(\registers[553][0] ), .C(
        \registers[554][0] ), .D(\registers[555][0] ), .S0(n4114), .S1(n4355), 
        .Y(n1350) );
  MX4X1 U8064 ( .A(\registers[712][0] ), .B(\registers[713][0] ), .C(
        \registers[714][0] ), .D(\registers[715][0] ), .S0(n4110), .S1(n4352), 
        .Y(n1202) );
  MX4X1 U8065 ( .A(\registers[760][0] ), .B(\registers[761][0] ), .C(
        \registers[762][0] ), .D(\registers[763][0] ), .S0(n4109), .S1(n4351), 
        .Y(n1173) );
  MX4X1 U8066 ( .A(\registers[744][0] ), .B(\registers[745][0] ), .C(
        \registers[746][0] ), .D(\registers[747][0] ), .S0(n4110), .S1(n4351), 
        .Y(n1178) );
  MX4X1 U8067 ( .A(\registers[648][0] ), .B(\registers[649][0] ), .C(
        \registers[650][0] ), .D(\registers[651][0] ), .S0(n4112), .S1(n4353), 
        .Y(n1301) );
  MX4X1 U8068 ( .A(\registers[696][0] ), .B(\registers[697][0] ), .C(
        \registers[698][0] ), .D(\registers[699][0] ), .S0(n4111), .S1(n4352), 
        .Y(n1270) );
  MX4X1 U8069 ( .A(\registers[680][0] ), .B(\registers[681][0] ), .C(
        \registers[682][0] ), .D(\registers[683][0] ), .S0(n4111), .S1(n4353), 
        .Y(n1281) );
  MX4X1 U8070 ( .A(\registers[328][1] ), .B(\registers[329][1] ), .C(
        \registers[330][1] ), .D(\registers[331][1] ), .S0(n4140), .S1(n4379), 
        .Y(n1787) );
  MX4X1 U8071 ( .A(\registers[376][1] ), .B(\registers[377][1] ), .C(
        \registers[378][1] ), .D(\registers[379][1] ), .S0(n4139), .S1(n4378), 
        .Y(n1771) );
  MX4X1 U8072 ( .A(\registers[360][1] ), .B(\registers[361][1] ), .C(
        \registers[362][1] ), .D(\registers[363][1] ), .S0(n4139), .S1(n4378), 
        .Y(n1777) );
  MX4X1 U8073 ( .A(\registers[72][1] ), .B(\registers[73][1] ), .C(
        \registers[74][1] ), .D(\registers[75][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1876) );
  MX4X1 U8074 ( .A(\registers[120][1] ), .B(\registers[121][1] ), .C(
        \registers[122][1] ), .D(\registers[123][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1859) );
  MX4X1 U8075 ( .A(\registers[104][1] ), .B(\registers[105][1] ), .C(
        \registers[106][1] ), .D(\registers[107][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1864) );
  MX4X1 U8076 ( .A(\registers[8][1] ), .B(\registers[9][1] ), .C(
        \registers[10][1] ), .D(\registers[11][1] ), .S0(n4146), .S1(n4385), 
        .Y(n1897) );
  MX4X1 U8077 ( .A(\registers[56][1] ), .B(\registers[57][1] ), .C(
        \registers[58][1] ), .D(\registers[59][1] ), .S0(n4145), .S1(n4384), 
        .Y(n1882) );
  MX4X1 U8078 ( .A(\registers[40][1] ), .B(\registers[41][1] ), .C(
        \registers[42][1] ), .D(\registers[43][1] ), .S0(n4146), .S1(n4385), 
        .Y(n1887) );
  MX4X1 U8079 ( .A(\registers[200][1] ), .B(\registers[201][1] ), .C(
        \registers[202][1] ), .D(\registers[203][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1831) );
  MX4X1 U8080 ( .A(\registers[248][1] ), .B(\registers[249][1] ), .C(
        \registers[250][1] ), .D(\registers[251][1] ), .S0(n4141), .S1(n4381), 
        .Y(n1816) );
  MX4X1 U8081 ( .A(\registers[232][1] ), .B(\registers[233][1] ), .C(
        \registers[234][1] ), .D(\registers[235][1] ), .S0(n4142), .S1(n4381), 
        .Y(n1821) );
  MX4X1 U8082 ( .A(\registers[136][1] ), .B(\registers[137][1] ), .C(
        \registers[138][1] ), .D(\registers[139][1] ), .S0(n4144), .S1(n4383), 
        .Y(n1853) );
  MX4X1 U8083 ( .A(\registers[184][1] ), .B(\registers[185][1] ), .C(
        \registers[186][1] ), .D(\registers[187][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1837) );
  MX4X1 U8084 ( .A(\registers[168][1] ), .B(\registers[169][1] ), .C(
        \registers[170][1] ), .D(\registers[171][1] ), .S0(n4143), .S1(n4382), 
        .Y(n1843) );
  MX4X1 U8085 ( .A(\registers[840][1] ), .B(\registers[841][1] ), .C(
        \registers[842][1] ), .D(\registers[843][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1612) );
  MX4X1 U8086 ( .A(\registers[888][1] ), .B(\registers[889][1] ), .C(
        \registers[890][1] ), .D(\registers[891][1] ), .S0(n4128), .S1(n4368), 
        .Y(n1594) );
  MX4X1 U8087 ( .A(\registers[872][1] ), .B(\registers[873][1] ), .C(
        \registers[874][1] ), .D(\registers[875][1] ), .S0(n4128), .S1(n4369), 
        .Y(n1599) );
  MX4X1 U8088 ( .A(\registers[776][1] ), .B(\registers[777][1] ), .C(
        \registers[778][1] ), .D(\registers[779][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1633) );
  MX4X1 U8089 ( .A(\registers[824][1] ), .B(\registers[825][1] ), .C(
        \registers[826][1] ), .D(\registers[827][1] ), .S0(n4129), .S1(n4369), 
        .Y(n1618) );
  MX4X1 U8090 ( .A(\registers[808][1] ), .B(\registers[809][1] ), .C(
        \registers[810][1] ), .D(\registers[811][1] ), .S0(n4130), .S1(n4370), 
        .Y(n1623) );
  MX4X1 U8091 ( .A(\registers[968][1] ), .B(\registers[969][1] ), .C(
        \registers[970][1] ), .D(\registers[971][1] ), .S0(n4126), .S1(n4367), 
        .Y(n1565) );
  MX4X1 U8092 ( .A(\registers[1016][1] ), .B(\registers[1017][1] ), .C(
        \registers[1018][1] ), .D(\registers[1019][1] ), .S0(n4125), .S1(n4366), .Y(n1550) );
  MX4X1 U8093 ( .A(\registers[1000][1] ), .B(\registers[1001][1] ), .C(
        \registers[1002][1] ), .D(\registers[1003][1] ), .S0(n4126), .S1(n4366), .Y(n1555) );
  MX4X1 U8094 ( .A(\registers[904][1] ), .B(\registers[905][1] ), .C(
        \registers[906][1] ), .D(\registers[907][1] ), .S0(n4128), .S1(n4368), 
        .Y(n1588) );
  MX4X1 U8095 ( .A(\registers[952][1] ), .B(\registers[953][1] ), .C(
        \registers[954][1] ), .D(\registers[955][1] ), .S0(n4127), .S1(n4367), 
        .Y(n1572) );
  MX4X1 U8096 ( .A(\registers[936][1] ), .B(\registers[937][1] ), .C(
        \registers[938][1] ), .D(\registers[939][1] ), .S0(n4127), .S1(n4367), 
        .Y(n1578) );
  MX4X1 U8097 ( .A(\registers[584][1] ), .B(\registers[585][1] ), .C(
        \registers[586][1] ), .D(\registers[587][1] ), .S0(n4134), .S1(n4374), 
        .Y(n1699) );
  MX4X1 U8098 ( .A(\registers[632][1] ), .B(\registers[633][1] ), .C(
        \registers[634][1] ), .D(\registers[635][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1684) );
  MX4X1 U8099 ( .A(\registers[616][1] ), .B(\registers[617][1] ), .C(
        \registers[618][1] ), .D(\registers[619][1] ), .S0(n4134), .S1(n4373), 
        .Y(n1689) );
  MX4X1 U8100 ( .A(\registers[520][1] ), .B(\registers[521][1] ), .C(
        \registers[522][1] ), .D(\registers[523][1] ), .S0(n4136), .S1(n4375), 
        .Y(n1721) );
  MX4X1 U8101 ( .A(\registers[568][1] ), .B(\registers[569][1] ), .C(
        \registers[570][1] ), .D(\registers[571][1] ), .S0(n4135), .S1(n4374), 
        .Y(n1705) );
  MX4X1 U8102 ( .A(\registers[552][1] ), .B(\registers[553][1] ), .C(
        \registers[554][1] ), .D(\registers[555][1] ), .S0(n4135), .S1(n4375), 
        .Y(n1711) );
  MX4X1 U8103 ( .A(\registers[712][1] ), .B(\registers[713][1] ), .C(
        \registers[714][1] ), .D(\registers[715][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1656) );
  MX4X1 U8104 ( .A(\registers[760][1] ), .B(\registers[761][1] ), .C(
        \registers[762][1] ), .D(\registers[763][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1640) );
  MX4X1 U8105 ( .A(\registers[744][1] ), .B(\registers[745][1] ), .C(
        \registers[746][1] ), .D(\registers[747][1] ), .S0(n4131), .S1(n4371), 
        .Y(n1646) );
  MX4X1 U8106 ( .A(\registers[648][1] ), .B(\registers[649][1] ), .C(
        \registers[650][1] ), .D(\registers[651][1] ), .S0(n4133), .S1(n4373), 
        .Y(n1678) );
  MX4X1 U8107 ( .A(\registers[696][1] ), .B(\registers[697][1] ), .C(
        \registers[698][1] ), .D(\registers[699][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1662) );
  MX4X1 U8108 ( .A(\registers[680][1] ), .B(\registers[681][1] ), .C(
        \registers[682][1] ), .D(\registers[683][1] ), .S0(n4132), .S1(n4372), 
        .Y(n1667) );
  MX4X1 U8109 ( .A(\registers[328][2] ), .B(\registers[329][2] ), .C(
        \registers[330][2] ), .D(\registers[331][2] ), .S0(n4161), .S1(n4399), 
        .Y(n2140) );
  MX4X1 U8110 ( .A(\registers[376][2] ), .B(\registers[377][2] ), .C(
        \registers[378][2] ), .D(\registers[379][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2123) );
  MX4X1 U8111 ( .A(\registers[360][2] ), .B(\registers[361][2] ), .C(
        \registers[362][2] ), .D(\registers[363][2] ), .S0(n4160), .S1(n4398), 
        .Y(n2128) );
  MX4X1 U8112 ( .A(\registers[72][2] ), .B(\registers[73][2] ), .C(
        \registers[74][2] ), .D(\registers[75][2] ), .S0(n4166), .S1(n4404), 
        .Y(n2227) );
  MX4X1 U8113 ( .A(\registers[120][2] ), .B(\registers[121][2] ), .C(
        \registers[122][2] ), .D(\registers[123][2] ), .S0(n4165), .S1(n4403), 
        .Y(n2212) );
  MX4X1 U8114 ( .A(\registers[104][2] ), .B(\registers[105][2] ), .C(
        \registers[106][2] ), .D(\registers[107][2] ), .S0(n4166), .S1(n4403), 
        .Y(n2217) );
  MX4X1 U8115 ( .A(\registers[8][2] ), .B(\registers[9][2] ), .C(
        \registers[10][2] ), .D(\registers[11][2] ), .S0(n4168), .S1(n4405), 
        .Y(n2249) );
  MX4X1 U8116 ( .A(\registers[56][2] ), .B(\registers[57][2] ), .C(
        \registers[58][2] ), .D(\registers[59][2] ), .S0(n4167), .S1(n4404), 
        .Y(n2233) );
  MX4X1 U8117 ( .A(\registers[40][2] ), .B(\registers[41][2] ), .C(
        \registers[42][2] ), .D(\registers[43][2] ), .S0(n4167), .S1(n4404), 
        .Y(n2239) );
  MX4X1 U8118 ( .A(\registers[200][2] ), .B(\registers[201][2] ), .C(
        \registers[202][2] ), .D(\registers[203][2] ), .S0(n4164), .S1(n4401), 
        .Y(n2184) );
  MX4X1 U8119 ( .A(\registers[248][2] ), .B(\registers[249][2] ), .C(
        \registers[250][2] ), .D(\registers[251][2] ), .S0(n4163), .S1(n4400), 
        .Y(n2168) );
  MX4X1 U8120 ( .A(\registers[232][2] ), .B(\registers[233][2] ), .C(
        \registers[234][2] ), .D(\registers[235][2] ), .S0(n4163), .S1(n4401), 
        .Y(n2174) );
  MX4X1 U8121 ( .A(\registers[136][2] ), .B(\registers[137][2] ), .C(
        \registers[138][2] ), .D(\registers[139][2] ), .S0(n4165), .S1(n4402), 
        .Y(n2206) );
  MX4X1 U8122 ( .A(\registers[184][2] ), .B(\registers[185][2] ), .C(
        \registers[186][2] ), .D(\registers[187][2] ), .S0(n4164), .S1(n4401), 
        .Y(n2190) );
  MX4X1 U8123 ( .A(\registers[168][2] ), .B(\registers[169][2] ), .C(
        \registers[170][2] ), .D(\registers[171][2] ), .S0(n4164), .S1(n4402), 
        .Y(n2195) );
  MX4X1 U8124 ( .A(\registers[840][2] ), .B(\registers[841][2] ), .C(
        \registers[842][2] ), .D(\registers[843][2] ), .S0(n4150), .S1(n4389), 
        .Y(n1963) );
  MX4X1 U8125 ( .A(\registers[888][2] ), .B(\registers[889][2] ), .C(
        \registers[890][2] ), .D(\registers[891][2] ), .S0(n4149), .S1(n4388), 
        .Y(n1948) );
  MX4X1 U8126 ( .A(\registers[872][2] ), .B(\registers[873][2] ), .C(
        \registers[874][2] ), .D(\registers[875][2] ), .S0(n4150), .S1(n4388), 
        .Y(n1953) );
  MX4X1 U8127 ( .A(\registers[776][2] ), .B(\registers[777][2] ), .C(
        \registers[778][2] ), .D(\registers[779][2] ), .S0(n4152), .S1(n4390), 
        .Y(n1985) );
  MX4X1 U8128 ( .A(\registers[824][2] ), .B(\registers[825][2] ), .C(
        \registers[826][2] ), .D(\registers[827][2] ), .S0(n4151), .S1(n4389), 
        .Y(n1969) );
  MX4X1 U8129 ( .A(\registers[808][2] ), .B(\registers[809][2] ), .C(
        \registers[810][2] ), .D(\registers[811][2] ), .S0(n4151), .S1(n4389), 
        .Y(n1975) );
  MX4X1 U8130 ( .A(\registers[968][2] ), .B(\registers[969][2] ), .C(
        \registers[970][2] ), .D(\registers[971][2] ), .S0(n4148), .S1(n4386), 
        .Y(n1920) );
  MX4X1 U8131 ( .A(\registers[1016][2] ), .B(\registers[1017][2] ), .C(
        \registers[1018][2] ), .D(\registers[1019][2] ), .S0(n4147), .S1(n4385), .Y(n1904) );
  MX4X1 U8132 ( .A(\registers[1000][2] ), .B(\registers[1001][2] ), .C(
        \registers[1002][2] ), .D(\registers[1003][2] ), .S0(n4147), .S1(n4386), .Y(n1910) );
  MX4X1 U8133 ( .A(\registers[904][2] ), .B(\registers[905][2] ), .C(
        \registers[906][2] ), .D(\registers[907][2] ), .S0(n4149), .S1(n4388), 
        .Y(n1942) );
  MX4X1 U8134 ( .A(\registers[952][2] ), .B(\registers[953][2] ), .C(
        \registers[954][2] ), .D(\registers[955][2] ), .S0(n4148), .S1(n4387), 
        .Y(n1926) );
  MX4X1 U8135 ( .A(\registers[936][2] ), .B(\registers[937][2] ), .C(
        \registers[938][2] ), .D(\registers[939][2] ), .S0(n4148), .S1(n4387), 
        .Y(n1931) );
  MX4X1 U8136 ( .A(\registers[584][2] ), .B(\registers[585][2] ), .C(
        \registers[586][2] ), .D(\registers[587][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2051) );
  MX4X1 U8137 ( .A(\registers[632][2] ), .B(\registers[633][2] ), .C(
        \registers[634][2] ), .D(\registers[635][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2035) );
  MX4X1 U8138 ( .A(\registers[616][2] ), .B(\registers[617][2] ), .C(
        \registers[618][2] ), .D(\registers[619][2] ), .S0(n4155), .S1(n4393), 
        .Y(n2041) );
  MX4X1 U8139 ( .A(\registers[520][2] ), .B(\registers[521][2] ), .C(
        \registers[522][2] ), .D(\registers[523][2] ), .S0(n4157), .S1(n4395), 
        .Y(n2073) );
  MX4X1 U8140 ( .A(\registers[568][2] ), .B(\registers[569][2] ), .C(
        \registers[570][2] ), .D(\registers[571][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2057) );
  MX4X1 U8141 ( .A(\registers[552][2] ), .B(\registers[553][2] ), .C(
        \registers[554][2] ), .D(\registers[555][2] ), .S0(n4156), .S1(n4394), 
        .Y(n2062) );
  MX4X1 U8142 ( .A(\registers[712][2] ), .B(\registers[713][2] ), .C(
        \registers[714][2] ), .D(\registers[715][2] ), .S0(n4153), .S1(n4391), 
        .Y(n2008) );
  MX4X1 U8143 ( .A(\registers[760][2] ), .B(\registers[761][2] ), .C(
        \registers[762][2] ), .D(\registers[763][2] ), .S0(n4152), .S1(n4390), 
        .Y(n1992) );
  MX4X1 U8144 ( .A(\registers[744][2] ), .B(\registers[745][2] ), .C(
        \registers[746][2] ), .D(\registers[747][2] ), .S0(n4152), .S1(n4391), 
        .Y(n1997) );
  MX4X1 U8145 ( .A(\registers[648][2] ), .B(\registers[649][2] ), .C(
        \registers[650][2] ), .D(\registers[651][2] ), .S0(n4154), .S1(n4393), 
        .Y(n2029) );
  MX4X1 U8146 ( .A(\registers[696][2] ), .B(\registers[697][2] ), .C(
        \registers[698][2] ), .D(\registers[699][2] ), .S0(n4153), .S1(n4392), 
        .Y(n2014) );
  MX4X1 U8147 ( .A(\registers[680][2] ), .B(\registers[681][2] ), .C(
        \registers[682][2] ), .D(\registers[683][2] ), .S0(n4154), .S1(n4392), 
        .Y(n2019) );
  MX4X1 U8148 ( .A(\registers[328][3] ), .B(\registers[329][3] ), .C(
        \registers[330][3] ), .D(\registers[331][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2553) );
  MX4X1 U8149 ( .A(\registers[376][3] ), .B(\registers[377][3] ), .C(
        \registers[378][3] ), .D(\registers[379][3] ), .S0(n4181), .S1(n4417), 
        .Y(n2538) );
  MX4X1 U8150 ( .A(\registers[360][3] ), .B(\registers[361][3] ), .C(
        \registers[362][3] ), .D(\registers[363][3] ), .S0(n4182), .S1(n4418), 
        .Y(n2543) );
  MX4X1 U8151 ( .A(\registers[72][3] ), .B(\registers[73][3] ), .C(
        \registers[74][3] ), .D(\registers[75][3] ), .S0(n4188), .S1(n4423), 
        .Y(n2638) );
  MX4X1 U8152 ( .A(\registers[120][3] ), .B(\registers[121][3] ), .C(
        \registers[122][3] ), .D(\registers[123][3] ), .S0(n4187), .S1(n4422), 
        .Y(n2623) );
  MX4X1 U8153 ( .A(\registers[104][3] ), .B(\registers[105][3] ), .C(
        \registers[106][3] ), .D(\registers[107][3] ), .S0(n4187), .S1(n4423), 
        .Y(n2628) );
  MX4X1 U8154 ( .A(\registers[8][3] ), .B(\registers[9][3] ), .C(
        \registers[10][3] ), .D(\registers[11][3] ), .S0(n4189), .S1(n4425), 
        .Y(n2659) );
  MX4X1 U8155 ( .A(\registers[56][3] ), .B(\registers[57][3] ), .C(
        \registers[58][3] ), .D(\registers[59][3] ), .S0(n4188), .S1(n4424), 
        .Y(n2644) );
  MX4X1 U8156 ( .A(\registers[40][3] ), .B(\registers[41][3] ), .C(
        \registers[42][3] ), .D(\registers[43][3] ), .S0(n4188), .S1(n4424), 
        .Y(n2649) );
  MX4X1 U8157 ( .A(\registers[200][3] ), .B(\registers[201][3] ), .C(
        \registers[202][3] ), .D(\registers[203][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2596) );
  MX4X1 U8158 ( .A(\registers[248][3] ), .B(\registers[249][3] ), .C(
        \registers[250][3] ), .D(\registers[251][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2581) );
  MX4X1 U8159 ( .A(\registers[232][3] ), .B(\registers[233][3] ), .C(
        \registers[234][3] ), .D(\registers[235][3] ), .S0(n4184), .S1(n4420), 
        .Y(n2586) );
  MX4X1 U8160 ( .A(\registers[136][3] ), .B(\registers[137][3] ), .C(
        \registers[138][3] ), .D(\registers[139][3] ), .S0(n4186), .S1(n4422), 
        .Y(n2617) );
  MX4X1 U8161 ( .A(\registers[184][3] ), .B(\registers[185][3] ), .C(
        \registers[186][3] ), .D(\registers[187][3] ), .S0(n4185), .S1(n4421), 
        .Y(n2602) );
  MX4X1 U8162 ( .A(\registers[168][3] ), .B(\registers[169][3] ), .C(
        \registers[170][3] ), .D(\registers[171][3] ), .S0(n4186), .S1(n4421), 
        .Y(n2607) );
  MX4X1 U8163 ( .A(\registers[840][3] ), .B(\registers[841][3] ), .C(
        \registers[842][3] ), .D(\registers[843][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2315) );
  MX4X1 U8164 ( .A(\registers[888][3] ), .B(\registers[889][3] ), .C(
        \registers[890][3] ), .D(\registers[891][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2299) );
  MX4X1 U8165 ( .A(\registers[872][3] ), .B(\registers[873][3] ), .C(
        \registers[874][3] ), .D(\registers[875][3] ), .S0(n4171), .S1(n4408), 
        .Y(n2305) );
  MX4X1 U8166 ( .A(\registers[776][3] ), .B(\registers[777][3] ), .C(
        \registers[778][3] ), .D(\registers[779][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2339) );
  MX4X1 U8167 ( .A(\registers[824][3] ), .B(\registers[825][3] ), .C(
        \registers[826][3] ), .D(\registers[827][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2321) );
  MX4X1 U8168 ( .A(\registers[808][3] ), .B(\registers[809][3] ), .C(
        \registers[810][3] ), .D(\registers[811][3] ), .S0(n4172), .S1(n4409), 
        .Y(n2326) );
  MX4X1 U8169 ( .A(\registers[968][3] ), .B(\registers[969][3] ), .C(
        \registers[970][3] ), .D(\registers[971][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2272) );
  MX4X1 U8170 ( .A(\registers[1016][3] ), .B(\registers[1017][3] ), .C(
        \registers[1018][3] ), .D(\registers[1019][3] ), .S0(n4168), .S1(n4405), .Y(n2256) );
  MX4X1 U8171 ( .A(\registers[1000][3] ), .B(\registers[1001][3] ), .C(
        \registers[1002][3] ), .D(\registers[1003][3] ), .S0(n4168), .S1(n4405), .Y(n2261) );
  MX4X1 U8172 ( .A(\registers[904][3] ), .B(\registers[905][3] ), .C(
        \registers[906][3] ), .D(\registers[907][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2293) );
  MX4X1 U8173 ( .A(\registers[952][3] ), .B(\registers[953][3] ), .C(
        \registers[954][3] ), .D(\registers[955][3] ), .S0(n4169), .S1(n4406), 
        .Y(n2278) );
  MX4X1 U8174 ( .A(\registers[936][3] ), .B(\registers[937][3] ), .C(
        \registers[938][3] ), .D(\registers[939][3] ), .S0(n4170), .S1(n4407), 
        .Y(n2283) );
  MX4X1 U8175 ( .A(\registers[584][3] ), .B(\registers[585][3] ), .C(
        \registers[586][3] ), .D(\registers[587][3] ), .S0(n4177), .S1(n4413), 
        .Y(n2468) );
  MX4X1 U8176 ( .A(\registers[632][3] ), .B(\registers[633][3] ), .C(
        \registers[634][3] ), .D(\registers[635][3] ), .S0(n4176), .S1(n4413), 
        .Y(n2453) );
  MX4X1 U8177 ( .A(\registers[616][3] ), .B(\registers[617][3] ), .C(
        \registers[618][3] ), .D(\registers[619][3] ), .S0(n4176), .S1(n4413), 
        .Y(n2458) );
  MX4X1 U8178 ( .A(\registers[520][3] ), .B(\registers[521][3] ), .C(
        \registers[522][3] ), .D(\registers[523][3] ), .S0(n4178), .S1(n4415), 
        .Y(n2489) );
  MX4X1 U8179 ( .A(\registers[568][3] ), .B(\registers[569][3] ), .C(
        \registers[570][3] ), .D(\registers[571][3] ), .S0(n4177), .S1(n4414), 
        .Y(n2474) );
  MX4X1 U8180 ( .A(\registers[552][3] ), .B(\registers[553][3] ), .C(
        \registers[554][3] ), .D(\registers[555][3] ), .S0(n4178), .S1(n4414), 
        .Y(n2479) );
  MX4X1 U8181 ( .A(\registers[712][3] ), .B(\registers[713][3] ), .C(
        \registers[714][3] ), .D(\registers[715][3] ), .S0(n4174), .S1(n4411), 
        .Y(n2370) );
  MX4X1 U8182 ( .A(\registers[760][3] ), .B(\registers[761][3] ), .C(
        \registers[762][3] ), .D(\registers[763][3] ), .S0(n4173), .S1(n4410), 
        .Y(n2353) );
  MX4X1 U8183 ( .A(\registers[744][3] ), .B(\registers[745][3] ), .C(
        \registers[746][3] ), .D(\registers[747][3] ), .S0(n4174), .S1(n4410), 
        .Y(n2359) );
  MX4X1 U8184 ( .A(\registers[648][3] ), .B(\registers[649][3] ), .C(
        \registers[650][3] ), .D(\registers[651][3] ), .S0(n4176), .S1(n4412), 
        .Y(n2447) );
  MX4X1 U8185 ( .A(\registers[696][3] ), .B(\registers[697][3] ), .C(
        \registers[698][3] ), .D(\registers[699][3] ), .S0(n4175), .S1(n4411), 
        .Y(n2377) );
  MX4X1 U8186 ( .A(\registers[680][3] ), .B(\registers[681][3] ), .C(
        \registers[682][3] ), .D(\registers[683][3] ), .S0(n4175), .S1(n4412), 
        .Y(n2437) );
  MX4X1 U8187 ( .A(\registers[328][4] ), .B(\registers[329][4] ), .C(
        \registers[330][4] ), .D(\registers[331][4] ), .S0(n4204), .S1(n4438), 
        .Y(n2893) );
  MX4X1 U8188 ( .A(\registers[376][4] ), .B(\registers[377][4] ), .C(
        \registers[378][4] ), .D(\registers[379][4] ), .S0(n4203), .S1(n4437), 
        .Y(n2878) );
  MX4X1 U8189 ( .A(\registers[360][4] ), .B(\registers[361][4] ), .C(
        \registers[362][4] ), .D(\registers[363][4] ), .S0(n4203), .S1(n4437), 
        .Y(n2883) );
  MX4X1 U8190 ( .A(\registers[72][4] ), .B(\registers[73][4] ), .C(
        \registers[74][4] ), .D(\registers[75][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2978) );
  MX4X1 U8191 ( .A(\registers[120][4] ), .B(\registers[121][4] ), .C(
        \registers[122][4] ), .D(\registers[123][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2963) );
  MX4X1 U8192 ( .A(\registers[104][4] ), .B(\registers[105][4] ), .C(
        \registers[106][4] ), .D(\registers[107][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2968) );
  MX4X1 U8193 ( .A(\registers[8][4] ), .B(\registers[9][4] ), .C(
        \registers[10][4] ), .D(\registers[11][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2999) );
  MX4X1 U8194 ( .A(\registers[56][4] ), .B(\registers[57][4] ), .C(
        \registers[58][4] ), .D(\registers[59][4] ), .S0(n4209), .S1(n4443), 
        .Y(n2984) );
  MX4X1 U8195 ( .A(\registers[40][4] ), .B(\registers[41][4] ), .C(
        \registers[42][4] ), .D(\registers[43][4] ), .S0(n4210), .S1(n4444), 
        .Y(n2989) );
  MX4X1 U8196 ( .A(\registers[200][4] ), .B(\registers[201][4] ), .C(
        \registers[202][4] ), .D(\registers[203][4] ), .S0(n4206), .S1(n4441), 
        .Y(n2936) );
  MX4X1 U8197 ( .A(\registers[248][4] ), .B(\registers[249][4] ), .C(
        \registers[250][4] ), .D(\registers[251][4] ), .S0(n4205), .S1(n4440), 
        .Y(n2921) );
  MX4X1 U8198 ( .A(\registers[232][4] ), .B(\registers[233][4] ), .C(
        \registers[234][4] ), .D(\registers[235][4] ), .S0(n4206), .S1(n4440), 
        .Y(n2926) );
  MX4X1 U8199 ( .A(\registers[136][4] ), .B(\registers[137][4] ), .C(
        \registers[138][4] ), .D(\registers[139][4] ), .S0(n4208), .S1(n4442), 
        .Y(n2957) );
  MX4X1 U8200 ( .A(\registers[184][4] ), .B(\registers[185][4] ), .C(
        \registers[186][4] ), .D(\registers[187][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2942) );
  MX4X1 U8201 ( .A(\registers[168][4] ), .B(\registers[169][4] ), .C(
        \registers[170][4] ), .D(\registers[171][4] ), .S0(n4207), .S1(n4441), 
        .Y(n2947) );
  MX4X1 U8202 ( .A(\registers[840][4] ), .B(\registers[841][4] ), .C(
        \registers[842][4] ), .D(\registers[843][4] ), .S0(n4193), .S1(n4428), 
        .Y(n2723) );
  MX4X1 U8203 ( .A(\registers[888][4] ), .B(\registers[889][4] ), .C(
        \registers[890][4] ), .D(\registers[891][4] ), .S0(n4192), .S1(n4427), 
        .Y(n2708) );
  MX4X1 U8204 ( .A(\registers[872][4] ), .B(\registers[873][4] ), .C(
        \registers[874][4] ), .D(\registers[875][4] ), .S0(n4192), .S1(n4428), 
        .Y(n2713) );
  MX4X1 U8205 ( .A(\registers[776][4] ), .B(\registers[777][4] ), .C(
        \registers[778][4] ), .D(\registers[779][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2744) );
  MX4X1 U8206 ( .A(\registers[824][4] ), .B(\registers[825][4] ), .C(
        \registers[826][4] ), .D(\registers[827][4] ), .S0(n4193), .S1(n4429), 
        .Y(n2729) );
  MX4X1 U8207 ( .A(\registers[808][4] ), .B(\registers[809][4] ), .C(
        \registers[810][4] ), .D(\registers[811][4] ), .S0(n4194), .S1(n4429), 
        .Y(n2734) );
  MX4X1 U8208 ( .A(\registers[968][4] ), .B(\registers[969][4] ), .C(
        \registers[970][4] ), .D(\registers[971][4] ), .S0(n4190), .S1(n4426), 
        .Y(n2681) );
  MX4X1 U8209 ( .A(\registers[1016][4] ), .B(\registers[1017][4] ), .C(
        \registers[1018][4] ), .D(\registers[1019][4] ), .S0(n4189), .S1(n4425), .Y(n2666) );
  MX4X1 U8210 ( .A(\registers[1000][4] ), .B(\registers[1001][4] ), .C(
        \registers[1002][4] ), .D(\registers[1003][4] ), .S0(n4190), .S1(n4425), .Y(n2671) );
  MX4X1 U8211 ( .A(\registers[904][4] ), .B(\registers[905][4] ), .C(
        \registers[906][4] ), .D(\registers[907][4] ), .S0(n4192), .S1(n4427), 
        .Y(n2702) );
  MX4X1 U8212 ( .A(\registers[952][4] ), .B(\registers[953][4] ), .C(
        \registers[954][4] ), .D(\registers[955][4] ), .S0(n4191), .S1(n4426), 
        .Y(n2687) );
  MX4X1 U8213 ( .A(\registers[936][4] ), .B(\registers[937][4] ), .C(
        \registers[938][4] ), .D(\registers[939][4] ), .S0(n4191), .S1(n4426), 
        .Y(n2692) );
  MX4X1 U8214 ( .A(\registers[584][4] ), .B(\registers[585][4] ), .C(
        \registers[586][4] ), .D(\registers[587][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2808) );
  MX4X1 U8215 ( .A(\registers[632][4] ), .B(\registers[633][4] ), .C(
        \registers[634][4] ), .D(\registers[635][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2793) );
  MX4X1 U8216 ( .A(\registers[616][4] ), .B(\registers[617][4] ), .C(
        \registers[618][4] ), .D(\registers[619][4] ), .S0(n4198), .S1(n4433), 
        .Y(n2798) );
  MX4X1 U8217 ( .A(\registers[520][4] ), .B(\registers[521][4] ), .C(
        \registers[522][4] ), .D(\registers[523][4] ), .S0(n4200), .S1(n4434), 
        .Y(n2829) );
  MX4X1 U8218 ( .A(\registers[568][4] ), .B(\registers[569][4] ), .C(
        \registers[570][4] ), .D(\registers[571][4] ), .S0(n4199), .S1(n4433), 
        .Y(n2814) );
  MX4X1 U8219 ( .A(\registers[552][4] ), .B(\registers[553][4] ), .C(
        \registers[554][4] ), .D(\registers[555][4] ), .S0(n4199), .S1(n4434), 
        .Y(n2819) );
  MX4X1 U8220 ( .A(\registers[712][4] ), .B(\registers[713][4] ), .C(
        \registers[714][4] ), .D(\registers[715][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2766) );
  MX4X1 U8221 ( .A(\registers[760][4] ), .B(\registers[761][4] ), .C(
        \registers[762][4] ), .D(\registers[763][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2751) );
  MX4X1 U8222 ( .A(\registers[744][4] ), .B(\registers[745][4] ), .C(
        \registers[746][4] ), .D(\registers[747][4] ), .S0(n4195), .S1(n4430), 
        .Y(n2756) );
  MX4X1 U8223 ( .A(\registers[648][4] ), .B(\registers[649][4] ), .C(
        \registers[650][4] ), .D(\registers[651][4] ), .S0(n4197), .S1(n4432), 
        .Y(n2787) );
  MX4X1 U8224 ( .A(\registers[696][4] ), .B(\registers[697][4] ), .C(
        \registers[698][4] ), .D(\registers[699][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2772) );
  MX4X1 U8225 ( .A(\registers[680][4] ), .B(\registers[681][4] ), .C(
        \registers[682][4] ), .D(\registers[683][4] ), .S0(n4196), .S1(n4431), 
        .Y(n2777) );
  MX4X1 U8226 ( .A(\registers[328][5] ), .B(\registers[329][5] ), .C(
        \registers[330][5] ), .D(\registers[331][5] ), .S0(n4225), .S1(n4458), 
        .Y(n3233) );
  MX4X1 U8227 ( .A(\registers[376][5] ), .B(\registers[377][5] ), .C(
        \registers[378][5] ), .D(\registers[379][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3218) );
  MX4X1 U8228 ( .A(\registers[360][5] ), .B(\registers[361][5] ), .C(
        \registers[362][5] ), .D(\registers[363][5] ), .S0(n4224), .S1(n4457), 
        .Y(n3223) );
  MX4X1 U8229 ( .A(\registers[72][5] ), .B(\registers[73][5] ), .C(
        \registers[74][5] ), .D(\registers[75][5] ), .S0(n4230), .S1(n4463), 
        .Y(n3318) );
  MX4X1 U8230 ( .A(\registers[120][5] ), .B(\registers[121][5] ), .C(
        \registers[122][5] ), .D(\registers[123][5] ), .S0(n4229), .S1(n4462), 
        .Y(n3303) );
  MX4X1 U8231 ( .A(\registers[104][5] ), .B(\registers[105][5] ), .C(
        \registers[106][5] ), .D(\registers[107][5] ), .S0(n4230), .S1(n4462), 
        .Y(n3308) );
  MX4X1 U8232 ( .A(\registers[8][5] ), .B(\registers[9][5] ), .C(
        \registers[10][5] ), .D(\registers[11][5] ), .S0(n4232), .S1(n4464), 
        .Y(n3339) );
  MX4X1 U8233 ( .A(\registers[56][5] ), .B(\registers[57][5] ), .C(
        \registers[58][5] ), .D(\registers[59][5] ), .S0(n4231), .S1(n4463), 
        .Y(n3324) );
  MX4X1 U8234 ( .A(\registers[40][5] ), .B(\registers[41][5] ), .C(
        \registers[42][5] ), .D(\registers[43][5] ), .S0(n4231), .S1(n4463), 
        .Y(n3329) );
  MX4X1 U8235 ( .A(\registers[200][5] ), .B(\registers[201][5] ), .C(
        \registers[202][5] ), .D(\registers[203][5] ), .S0(n4228), .S1(n4460), 
        .Y(n3276) );
  MX4X1 U8236 ( .A(\registers[248][5] ), .B(\registers[249][5] ), .C(
        \registers[250][5] ), .D(\registers[251][5] ), .S0(n4227), .S1(n4459), 
        .Y(n3261) );
  MX4X1 U8237 ( .A(\registers[232][5] ), .B(\registers[233][5] ), .C(
        \registers[234][5] ), .D(\registers[235][5] ), .S0(n4227), .S1(n4460), 
        .Y(n3266) );
  MX4X1 U8238 ( .A(\registers[136][5] ), .B(\registers[137][5] ), .C(
        \registers[138][5] ), .D(\registers[139][5] ), .S0(n4229), .S1(n4461), 
        .Y(n3297) );
  MX4X1 U8239 ( .A(\registers[184][5] ), .B(\registers[185][5] ), .C(
        \registers[186][5] ), .D(\registers[187][5] ), .S0(n4228), .S1(n4461), 
        .Y(n3282) );
  MX4X1 U8240 ( .A(\registers[168][5] ), .B(\registers[169][5] ), .C(
        \registers[170][5] ), .D(\registers[171][5] ), .S0(n4228), .S1(n4461), 
        .Y(n3287) );
  MX4X1 U8241 ( .A(\registers[840][5] ), .B(\registers[841][5] ), .C(
        \registers[842][5] ), .D(\registers[843][5] ), .S0(n4214), .S1(n4448), 
        .Y(n3063) );
  MX4X1 U8242 ( .A(\registers[888][5] ), .B(\registers[889][5] ), .C(
        \registers[890][5] ), .D(\registers[891][5] ), .S0(n4213), .S1(n4447), 
        .Y(n3048) );
  MX4X1 U8243 ( .A(\registers[872][5] ), .B(\registers[873][5] ), .C(
        \registers[874][5] ), .D(\registers[875][5] ), .S0(n4214), .S1(n4447), 
        .Y(n3053) );
  MX4X1 U8244 ( .A(\registers[776][5] ), .B(\registers[777][5] ), .C(
        \registers[778][5] ), .D(\registers[779][5] ), .S0(n4216), .S1(n4449), 
        .Y(n3084) );
  MX4X1 U8245 ( .A(\registers[824][5] ), .B(\registers[825][5] ), .C(
        \registers[826][5] ), .D(\registers[827][5] ), .S0(n4215), .S1(n4448), 
        .Y(n3069) );
  MX4X1 U8246 ( .A(\registers[808][5] ), .B(\registers[809][5] ), .C(
        \registers[810][5] ), .D(\registers[811][5] ), .S0(n4215), .S1(n4449), 
        .Y(n3074) );
  MX4X1 U8247 ( .A(\registers[968][5] ), .B(\registers[969][5] ), .C(
        \registers[970][5] ), .D(\registers[971][5] ), .S0(n4212), .S1(n4445), 
        .Y(n3021) );
  MX4X1 U8248 ( .A(\registers[1016][5] ), .B(\registers[1017][5] ), .C(
        \registers[1018][5] ), .D(\registers[1019][5] ), .S0(n4211), .S1(n4445), .Y(n3006) );
  MX4X1 U8249 ( .A(\registers[1000][5] ), .B(\registers[1001][5] ), .C(
        \registers[1002][5] ), .D(\registers[1003][5] ), .S0(n4211), .S1(n4445), .Y(n3011) );
  MX4X1 U8250 ( .A(\registers[904][5] ), .B(\registers[905][5] ), .C(
        \registers[906][5] ), .D(\registers[907][5] ), .S0(n4213), .S1(n4447), 
        .Y(n3042) );
  MX4X1 U8251 ( .A(\registers[952][5] ), .B(\registers[953][5] ), .C(
        \registers[954][5] ), .D(\registers[955][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3027) );
  MX4X1 U8252 ( .A(\registers[936][5] ), .B(\registers[937][5] ), .C(
        \registers[938][5] ), .D(\registers[939][5] ), .S0(n4212), .S1(n4446), 
        .Y(n3032) );
  MX4X1 U8253 ( .A(\registers[584][5] ), .B(\registers[585][5] ), .C(
        \registers[586][5] ), .D(\registers[587][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3148) );
  MX4X1 U8254 ( .A(\registers[632][5] ), .B(\registers[633][5] ), .C(
        \registers[634][5] ), .D(\registers[635][5] ), .S0(n4219), .S1(n4452), 
        .Y(n3133) );
  MX4X1 U8255 ( .A(\registers[616][5] ), .B(\registers[617][5] ), .C(
        \registers[618][5] ), .D(\registers[619][5] ), .S0(n4219), .S1(n4452), 
        .Y(n3138) );
  MX4X1 U8256 ( .A(\registers[520][5] ), .B(\registers[521][5] ), .C(
        \registers[522][5] ), .D(\registers[523][5] ), .S0(n4221), .S1(n4454), 
        .Y(n3169) );
  MX4X1 U8257 ( .A(\registers[568][5] ), .B(\registers[569][5] ), .C(
        \registers[570][5] ), .D(\registers[571][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3154) );
  MX4X1 U8258 ( .A(\registers[552][5] ), .B(\registers[553][5] ), .C(
        \registers[554][5] ), .D(\registers[555][5] ), .S0(n4220), .S1(n4453), 
        .Y(n3159) );
  MX4X1 U8259 ( .A(\registers[712][5] ), .B(\registers[713][5] ), .C(
        \registers[714][5] ), .D(\registers[715][5] ), .S0(n4217), .S1(n4450), 
        .Y(n3106) );
  MX4X1 U8260 ( .A(\registers[760][5] ), .B(\registers[761][5] ), .C(
        \registers[762][5] ), .D(\registers[763][5] ), .S0(n4216), .S1(n4449), 
        .Y(n3091) );
  MX4X1 U8261 ( .A(\registers[744][5] ), .B(\registers[745][5] ), .C(
        \registers[746][5] ), .D(\registers[747][5] ), .S0(n4216), .S1(n4450), 
        .Y(n3096) );
  MX4X1 U8262 ( .A(\registers[648][5] ), .B(\registers[649][5] ), .C(
        \registers[650][5] ), .D(\registers[651][5] ), .S0(n4218), .S1(n4452), 
        .Y(n3127) );
  MX4X1 U8263 ( .A(\registers[696][5] ), .B(\registers[697][5] ), .C(
        \registers[698][5] ), .D(\registers[699][5] ), .S0(n4217), .S1(n4451), 
        .Y(n3112) );
  MX4X1 U8264 ( .A(\registers[680][5] ), .B(\registers[681][5] ), .C(
        \registers[682][5] ), .D(\registers[683][5] ), .S0(n4218), .S1(n4451), 
        .Y(n3117) );
  MX4X1 U8265 ( .A(\registers[328][6] ), .B(\registers[329][6] ), .C(
        \registers[330][6] ), .D(\registers[331][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3573) );
  MX4X1 U8266 ( .A(\registers[376][6] ), .B(\registers[377][6] ), .C(
        \registers[378][6] ), .D(\registers[379][6] ), .S0(n4245), .S1(n4477), 
        .Y(n3558) );
  MX4X1 U8267 ( .A(\registers[360][6] ), .B(\registers[361][6] ), .C(
        \registers[362][6] ), .D(\registers[363][6] ), .S0(n4246), .S1(n4477), 
        .Y(n3563) );
  MX4X1 U8268 ( .A(\registers[72][6] ), .B(\registers[73][6] ), .C(
        \registers[74][6] ), .D(\registers[75][6] ), .S0(n4252), .S1(n4482), 
        .Y(n3658) );
  MX4X1 U8269 ( .A(\registers[120][6] ), .B(\registers[121][6] ), .C(
        \registers[122][6] ), .D(\registers[123][6] ), .S0(n4251), .S1(n4481), 
        .Y(n3643) );
  MX4X1 U8270 ( .A(\registers[104][6] ), .B(\registers[105][6] ), .C(
        \registers[106][6] ), .D(\registers[107][6] ), .S0(n4251), .S1(n4482), 
        .Y(n3648) );
  MX4X1 U8271 ( .A(\registers[8][6] ), .B(\registers[9][6] ), .C(
        \registers[10][6] ), .D(\registers[11][6] ), .S0(n4253), .S1(n4484), 
        .Y(n3679) );
  MX4X1 U8272 ( .A(\registers[56][6] ), .B(\registers[57][6] ), .C(
        \registers[58][6] ), .D(\registers[59][6] ), .S0(n4252), .S1(n4483), 
        .Y(n3664) );
  MX4X1 U8273 ( .A(\registers[40][6] ), .B(\registers[41][6] ), .C(
        \registers[42][6] ), .D(\registers[43][6] ), .S0(n4252), .S1(n4483), 
        .Y(n3669) );
  MX4X1 U8274 ( .A(\registers[200][6] ), .B(\registers[201][6] ), .C(
        \registers[202][6] ), .D(\registers[203][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3616) );
  MX4X1 U8275 ( .A(\registers[248][6] ), .B(\registers[249][6] ), .C(
        \registers[250][6] ), .D(\registers[251][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3601) );
  MX4X1 U8276 ( .A(\registers[232][6] ), .B(\registers[233][6] ), .C(
        \registers[234][6] ), .D(\registers[235][6] ), .S0(n4248), .S1(n4479), 
        .Y(n3606) );
  MX4X1 U8277 ( .A(\registers[136][6] ), .B(\registers[137][6] ), .C(
        \registers[138][6] ), .D(\registers[139][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3637) );
  MX4X1 U8278 ( .A(\registers[184][6] ), .B(\registers[185][6] ), .C(
        \registers[186][6] ), .D(\registers[187][6] ), .S0(n4249), .S1(n4480), 
        .Y(n3622) );
  MX4X1 U8279 ( .A(\registers[168][6] ), .B(\registers[169][6] ), .C(
        \registers[170][6] ), .D(\registers[171][6] ), .S0(n4250), .S1(n4481), 
        .Y(n3627) );
  MX4X1 U8280 ( .A(\registers[840][6] ), .B(\registers[841][6] ), .C(
        \registers[842][6] ), .D(\registers[843][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3403) );
  MX4X1 U8281 ( .A(\registers[888][6] ), .B(\registers[889][6] ), .C(
        \registers[890][6] ), .D(\registers[891][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3388) );
  MX4X1 U8282 ( .A(\registers[872][6] ), .B(\registers[873][6] ), .C(
        \registers[874][6] ), .D(\registers[875][6] ), .S0(n4235), .S1(n4467), 
        .Y(n3393) );
  MX4X1 U8283 ( .A(\registers[776][6] ), .B(\registers[777][6] ), .C(
        \registers[778][6] ), .D(\registers[779][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3424) );
  MX4X1 U8284 ( .A(\registers[824][6] ), .B(\registers[825][6] ), .C(
        \registers[826][6] ), .D(\registers[827][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3409) );
  MX4X1 U8285 ( .A(\registers[808][6] ), .B(\registers[809][6] ), .C(
        \registers[810][6] ), .D(\registers[811][6] ), .S0(n4236), .S1(n4468), 
        .Y(n3414) );
  MX4X1 U8286 ( .A(\registers[968][6] ), .B(\registers[969][6] ), .C(
        \registers[970][6] ), .D(\registers[971][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3361) );
  MX4X1 U8287 ( .A(\registers[1016][6] ), .B(\registers[1017][6] ), .C(
        \registers[1018][6] ), .D(\registers[1019][6] ), .S0(n4232), .S1(n4464), .Y(n3346) );
  MX4X1 U8288 ( .A(\registers[1000][6] ), .B(\registers[1001][6] ), .C(
        \registers[1002][6] ), .D(\registers[1003][6] ), .S0(n4232), .S1(n4465), .Y(n3351) );
  MX4X1 U8289 ( .A(\registers[904][6] ), .B(\registers[905][6] ), .C(
        \registers[906][6] ), .D(\registers[907][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3382) );
  MX4X1 U8290 ( .A(\registers[952][6] ), .B(\registers[953][6] ), .C(
        \registers[954][6] ), .D(\registers[955][6] ), .S0(n4233), .S1(n4465), 
        .Y(n3367) );
  MX4X1 U8291 ( .A(\registers[936][6] ), .B(\registers[937][6] ), .C(
        \registers[938][6] ), .D(\registers[939][6] ), .S0(n4234), .S1(n4466), 
        .Y(n3372) );
  MX4X1 U8292 ( .A(\registers[584][6] ), .B(\registers[585][6] ), .C(
        \registers[586][6] ), .D(\registers[587][6] ), .S0(n4241), .S1(n4473), 
        .Y(n3488) );
  MX4X1 U8293 ( .A(\registers[632][6] ), .B(\registers[633][6] ), .C(
        \registers[634][6] ), .D(\registers[635][6] ), .S0(n4240), .S1(n4472), 
        .Y(n3473) );
  MX4X1 U8294 ( .A(\registers[616][6] ), .B(\registers[617][6] ), .C(
        \registers[618][6] ), .D(\registers[619][6] ), .S0(n4240), .S1(n4472), 
        .Y(n3478) );
  MX4X1 U8295 ( .A(\registers[520][6] ), .B(\registers[521][6] ), .C(
        \registers[522][6] ), .D(\registers[523][6] ), .S0(n4242), .S1(n4474), 
        .Y(n3509) );
  MX4X1 U8296 ( .A(\registers[568][6] ), .B(\registers[569][6] ), .C(
        \registers[570][6] ), .D(\registers[571][6] ), .S0(n4241), .S1(n4473), 
        .Y(n3494) );
  MX4X1 U8297 ( .A(\registers[552][6] ), .B(\registers[553][6] ), .C(
        \registers[554][6] ), .D(\registers[555][6] ), .S0(n4242), .S1(n4473), 
        .Y(n3499) );
  MX4X1 U8298 ( .A(\registers[712][6] ), .B(\registers[713][6] ), .C(
        \registers[714][6] ), .D(\registers[715][6] ), .S0(n4238), .S1(n4470), 
        .Y(n3446) );
  MX4X1 U8299 ( .A(\registers[760][6] ), .B(\registers[761][6] ), .C(
        \registers[762][6] ), .D(\registers[763][6] ), .S0(n4237), .S1(n4469), 
        .Y(n3431) );
  MX4X1 U8300 ( .A(\registers[744][6] ), .B(\registers[745][6] ), .C(
        \registers[746][6] ), .D(\registers[747][6] ), .S0(n4238), .S1(n4469), 
        .Y(n3436) );
  MX4X1 U8301 ( .A(\registers[648][6] ), .B(\registers[649][6] ), .C(
        \registers[650][6] ), .D(\registers[651][6] ), .S0(n4240), .S1(n4471), 
        .Y(n3467) );
  MX4X1 U8302 ( .A(\registers[696][6] ), .B(\registers[697][6] ), .C(
        \registers[698][6] ), .D(\registers[699][6] ), .S0(n4239), .S1(n4470), 
        .Y(n3452) );
  MX4X1 U8303 ( .A(\registers[680][6] ), .B(\registers[681][6] ), .C(
        \registers[682][6] ), .D(\registers[683][6] ), .S0(n4239), .S1(n4471), 
        .Y(n3457) );
  MX4X1 U8304 ( .A(\registers[328][7] ), .B(\registers[329][7] ), .C(
        \registers[330][7] ), .D(\registers[331][7] ), .S0(n4268), .S1(n4483), 
        .Y(n3913) );
  MX4X1 U8305 ( .A(\registers[376][7] ), .B(\registers[377][7] ), .C(
        \registers[378][7] ), .D(\registers[379][7] ), .S0(n4267), .S1(n4496), 
        .Y(n3898) );
  MX4X1 U8306 ( .A(\registers[360][7] ), .B(\registers[361][7] ), .C(
        \registers[362][7] ), .D(\registers[363][7] ), .S0(n4267), .S1(n4473), 
        .Y(n3903) );
  MX4X1 U8307 ( .A(\registers[72][7] ), .B(\registers[73][7] ), .C(
        \registers[74][7] ), .D(\registers[75][7] ), .S0(n4273), .S1(n4297), 
        .Y(n3998) );
  MX4X1 U8308 ( .A(\registers[120][7] ), .B(\registers[121][7] ), .C(
        \registers[122][7] ), .D(\registers[123][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3983) );
  MX4X1 U8309 ( .A(\registers[104][7] ), .B(\registers[105][7] ), .C(
        \registers[106][7] ), .D(\registers[107][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3988) );
  MX4X1 U8310 ( .A(\registers[8][7] ), .B(\registers[9][7] ), .C(
        \registers[10][7] ), .D(\registers[11][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4019) );
  MX4X1 U8311 ( .A(\registers[56][7] ), .B(\registers[57][7] ), .C(
        \registers[58][7] ), .D(\registers[59][7] ), .S0(n4273), .S1(n4492), 
        .Y(n4004) );
  MX4X1 U8312 ( .A(\registers[40][7] ), .B(\registers[41][7] ), .C(
        \registers[42][7] ), .D(\registers[43][7] ), .S0(n4274), .S1(n4501), 
        .Y(n4009) );
  MX4X1 U8313 ( .A(\registers[200][7] ), .B(\registers[201][7] ), .C(
        \registers[202][7] ), .D(\registers[203][7] ), .S0(n4270), .S1(n4499), 
        .Y(n3956) );
  MX4X1 U8314 ( .A(\registers[248][7] ), .B(\registers[249][7] ), .C(
        \registers[250][7] ), .D(\registers[251][7] ), .S0(n4269), .S1(n4498), 
        .Y(n3941) );
  MX4X1 U8315 ( .A(\registers[232][7] ), .B(\registers[233][7] ), .C(
        \registers[234][7] ), .D(\registers[235][7] ), .S0(n4270), .S1(n4498), 
        .Y(n3946) );
  MX4X1 U8316 ( .A(\registers[136][7] ), .B(\registers[137][7] ), .C(
        \registers[138][7] ), .D(\registers[139][7] ), .S0(n4272), .S1(n4500), 
        .Y(n3977) );
  MX4X1 U8317 ( .A(\registers[184][7] ), .B(\registers[185][7] ), .C(
        \registers[186][7] ), .D(\registers[187][7] ), .S0(n4271), .S1(n4499), 
        .Y(n3962) );
  MX4X1 U8318 ( .A(\registers[168][7] ), .B(\registers[169][7] ), .C(
        \registers[170][7] ), .D(\registers[171][7] ), .S0(n4271), .S1(n4499), 
        .Y(n3967) );
  MX4X1 U8319 ( .A(\registers[840][7] ), .B(\registers[841][7] ), .C(
        \registers[842][7] ), .D(\registers[843][7] ), .S0(n4257), .S1(n4487), 
        .Y(n3743) );
  MX4X1 U8320 ( .A(\registers[888][7] ), .B(\registers[889][7] ), .C(
        \registers[890][7] ), .D(\registers[891][7] ), .S0(n4256), .S1(n4486), 
        .Y(n3728) );
  MX4X1 U8321 ( .A(\registers[872][7] ), .B(\registers[873][7] ), .C(
        \registers[874][7] ), .D(\registers[875][7] ), .S0(n4256), .S1(n4487), 
        .Y(n3733) );
  MX4X1 U8322 ( .A(\registers[776][7] ), .B(\registers[777][7] ), .C(
        \registers[778][7] ), .D(\registers[779][7] ), .S0(n4258), .S1(n4489), 
        .Y(n3764) );
  MX4X1 U8323 ( .A(\registers[824][7] ), .B(\registers[825][7] ), .C(
        \registers[826][7] ), .D(\registers[827][7] ), .S0(n4257), .S1(n4488), 
        .Y(n3749) );
  MX4X1 U8324 ( .A(\registers[808][7] ), .B(\registers[809][7] ), .C(
        \registers[810][7] ), .D(\registers[811][7] ), .S0(n4258), .S1(n4488), 
        .Y(n3754) );
  MX4X1 U8325 ( .A(\registers[968][7] ), .B(\registers[969][7] ), .C(
        \registers[970][7] ), .D(\registers[971][7] ), .S0(n4254), .S1(n4485), 
        .Y(n3701) );
  MX4X1 U8326 ( .A(\registers[1016][7] ), .B(\registers[1017][7] ), .C(
        \registers[1018][7] ), .D(\registers[1019][7] ), .S0(n4253), .S1(n4484), .Y(n3686) );
  MX4X1 U8327 ( .A(\registers[1000][7] ), .B(\registers[1001][7] ), .C(
        \registers[1002][7] ), .D(\registers[1003][7] ), .S0(n4254), .S1(n4484), .Y(n3691) );
  MX4X1 U8328 ( .A(\registers[904][7] ), .B(\registers[905][7] ), .C(
        \registers[906][7] ), .D(\registers[907][7] ), .S0(n4256), .S1(n4486), 
        .Y(n3722) );
  MX4X1 U8329 ( .A(\registers[952][7] ), .B(\registers[953][7] ), .C(
        \registers[954][7] ), .D(\registers[955][7] ), .S0(n4255), .S1(n4485), 
        .Y(n3707) );
  MX4X1 U8330 ( .A(\registers[936][7] ), .B(\registers[937][7] ), .C(
        \registers[938][7] ), .D(\registers[939][7] ), .S0(n4255), .S1(n4485), 
        .Y(n3712) );
  MX4X1 U8331 ( .A(\registers[584][7] ), .B(\registers[585][7] ), .C(
        \registers[586][7] ), .D(\registers[587][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3828) );
  MX4X1 U8332 ( .A(\registers[632][7] ), .B(\registers[633][7] ), .C(
        \registers[634][7] ), .D(\registers[635][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3813) );
  MX4X1 U8333 ( .A(\registers[616][7] ), .B(\registers[617][7] ), .C(
        \registers[618][7] ), .D(\registers[619][7] ), .S0(n4262), .S1(n4492), 
        .Y(n3818) );
  MX4X1 U8334 ( .A(\registers[520][7] ), .B(\registers[521][7] ), .C(
        \registers[522][7] ), .D(\registers[523][7] ), .S0(n4264), .S1(n4493), 
        .Y(n3849) );
  MX4X1 U8335 ( .A(\registers[568][7] ), .B(\registers[569][7] ), .C(
        \registers[570][7] ), .D(\registers[571][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3834) );
  MX4X1 U8336 ( .A(\registers[552][7] ), .B(\registers[553][7] ), .C(
        \registers[554][7] ), .D(\registers[555][7] ), .S0(n4263), .S1(n4493), 
        .Y(n3839) );
  MX4X1 U8337 ( .A(\registers[712][7] ), .B(\registers[713][7] ), .C(
        \registers[714][7] ), .D(\registers[715][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3786) );
  MX4X1 U8338 ( .A(\registers[760][7] ), .B(\registers[761][7] ), .C(
        \registers[762][7] ), .D(\registers[763][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3771) );
  MX4X1 U8339 ( .A(\registers[744][7] ), .B(\registers[745][7] ), .C(
        \registers[746][7] ), .D(\registers[747][7] ), .S0(n4259), .S1(n4489), 
        .Y(n3776) );
  MX4X1 U8340 ( .A(\registers[648][7] ), .B(\registers[649][7] ), .C(
        \registers[650][7] ), .D(\registers[651][7] ), .S0(n4261), .S1(n4491), 
        .Y(n3807) );
  MX4X1 U8341 ( .A(\registers[696][7] ), .B(\registers[697][7] ), .C(
        \registers[698][7] ), .D(\registers[699][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3792) );
  MX4X1 U8342 ( .A(\registers[680][7] ), .B(\registers[681][7] ), .C(
        \registers[682][7] ), .D(\registers[683][7] ), .S0(n4260), .S1(n4490), 
        .Y(n3797) );
  MX4X1 U8343 ( .A(\registers[328][0] ), .B(\registers[329][0] ), .C(
        \registers[330][0] ), .D(\registers[331][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4878) );
  MX4X1 U8344 ( .A(\registers[376][0] ), .B(\registers[377][0] ), .C(
        \registers[378][0] ), .D(\registers[379][0] ), .S0(n7460), .S1(n7702), 
        .Y(n4863) );
  MX4X1 U8345 ( .A(\registers[360][0] ), .B(\registers[361][0] ), .C(
        \registers[362][0] ), .D(\registers[363][0] ), .S0(n7461), .S1(n7703), 
        .Y(n4868) );
  MX4X1 U8346 ( .A(\registers[72][0] ), .B(\registers[73][0] ), .C(
        \registers[74][0] ), .D(\registers[75][0] ), .S0(n7467), .S1(n7708), 
        .Y(n4963) );
  MX4X1 U8347 ( .A(\registers[120][0] ), .B(\registers[121][0] ), .C(
        \registers[122][0] ), .D(\registers[123][0] ), .S0(n7466), .S1(n7707), 
        .Y(n4948) );
  MX4X1 U8348 ( .A(\registers[104][0] ), .B(\registers[105][0] ), .C(
        \registers[106][0] ), .D(\registers[107][0] ), .S0(n7466), .S1(n7708), 
        .Y(n4953) );
  MX4X1 U8349 ( .A(\registers[8][0] ), .B(\registers[9][0] ), .C(
        \registers[10][0] ), .D(\registers[11][0] ), .S0(n7468), .S1(n7709), 
        .Y(n4984) );
  MX4X1 U8350 ( .A(\registers[56][0] ), .B(\registers[57][0] ), .C(
        \registers[58][0] ), .D(\registers[59][0] ), .S0(n7467), .S1(n7709), 
        .Y(n4969) );
  MX4X1 U8351 ( .A(\registers[40][0] ), .B(\registers[41][0] ), .C(
        \registers[42][0] ), .D(\registers[43][0] ), .S0(n7467), .S1(n7709), 
        .Y(n4974) );
  MX4X1 U8352 ( .A(\registers[200][0] ), .B(\registers[201][0] ), .C(
        \registers[202][0] ), .D(\registers[203][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4921) );
  MX4X1 U8353 ( .A(\registers[248][0] ), .B(\registers[249][0] ), .C(
        \registers[250][0] ), .D(\registers[251][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4906) );
  MX4X1 U8354 ( .A(\registers[232][0] ), .B(\registers[233][0] ), .C(
        \registers[234][0] ), .D(\registers[235][0] ), .S0(n7463), .S1(n7705), 
        .Y(n4911) );
  MX4X1 U8355 ( .A(\registers[136][0] ), .B(\registers[137][0] ), .C(
        \registers[138][0] ), .D(\registers[139][0] ), .S0(n7465), .S1(n7707), 
        .Y(n4942) );
  MX4X1 U8356 ( .A(\registers[184][0] ), .B(\registers[185][0] ), .C(
        \registers[186][0] ), .D(\registers[187][0] ), .S0(n7464), .S1(n7706), 
        .Y(n4927) );
  MX4X1 U8357 ( .A(\registers[168][0] ), .B(\registers[169][0] ), .C(
        \registers[170][0] ), .D(\registers[171][0] ), .S0(n7465), .S1(n7706), 
        .Y(n4932) );
  MX4X1 U8358 ( .A(\registers[840][0] ), .B(\registers[841][0] ), .C(
        \registers[842][0] ), .D(\registers[843][0] ), .S0(n7451), .S1(n7693), 
        .Y(n4708) );
  MX4X1 U8359 ( .A(\registers[888][0] ), .B(\registers[889][0] ), .C(
        \registers[890][0] ), .D(\registers[891][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4693) );
  MX4X1 U8360 ( .A(\registers[872][0] ), .B(\registers[873][0] ), .C(
        \registers[874][0] ), .D(\registers[875][0] ), .S0(n7450), .S1(n7693), 
        .Y(n4698) );
  MX4X1 U8361 ( .A(\registers[776][0] ), .B(\registers[777][0] ), .C(
        \registers[778][0] ), .D(\registers[779][0] ), .S0(n7452), .S1(n7695), 
        .Y(n4729) );
  MX4X1 U8362 ( .A(\registers[824][0] ), .B(\registers[825][0] ), .C(
        \registers[826][0] ), .D(\registers[827][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4714) );
  MX4X1 U8363 ( .A(\registers[808][0] ), .B(\registers[809][0] ), .C(
        \registers[810][0] ), .D(\registers[811][0] ), .S0(n7451), .S1(n7694), 
        .Y(n4719) );
  MX4X1 U8364 ( .A(\registers[968][0] ), .B(\registers[969][0] ), .C(
        \registers[970][0] ), .D(\registers[971][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4666) );
  MX4X1 U8365 ( .A(\registers[904][0] ), .B(\registers[905][0] ), .C(
        \registers[906][0] ), .D(\registers[907][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4687) );
  MX4X1 U8366 ( .A(\registers[952][0] ), .B(\registers[953][0] ), .C(
        \registers[954][0] ), .D(\registers[955][0] ), .S0(n7448), .S1(n7691), 
        .Y(n4672) );
  MX4X1 U8367 ( .A(\registers[936][0] ), .B(\registers[937][0] ), .C(
        \registers[938][0] ), .D(\registers[939][0] ), .S0(n7449), .S1(n7692), 
        .Y(n4677) );
  MX4X1 U8368 ( .A(\registers[584][0] ), .B(\registers[585][0] ), .C(
        \registers[586][0] ), .D(\registers[587][0] ), .S0(n7456), .S1(n7698), 
        .Y(n4793) );
  MX4X1 U8369 ( .A(\registers[632][0] ), .B(\registers[633][0] ), .C(
        \registers[634][0] ), .D(\registers[635][0] ), .S0(n7455), .S1(n7697), 
        .Y(n4778) );
  MX4X1 U8370 ( .A(\registers[616][0] ), .B(\registers[617][0] ), .C(
        \registers[618][0] ), .D(\registers[619][0] ), .S0(n7455), .S1(n7698), 
        .Y(n4783) );
  MX4X1 U8371 ( .A(\registers[520][0] ), .B(\registers[521][0] ), .C(
        \registers[522][0] ), .D(\registers[523][0] ), .S0(n7457), .S1(n7700), 
        .Y(n4814) );
  MX4X1 U8372 ( .A(\registers[568][0] ), .B(\registers[569][0] ), .C(
        \registers[570][0] ), .D(\registers[571][0] ), .S0(n7456), .S1(n7699), 
        .Y(n4799) );
  MX4X1 U8373 ( .A(\registers[552][0] ), .B(\registers[553][0] ), .C(
        \registers[554][0] ), .D(\registers[555][0] ), .S0(n7457), .S1(n7699), 
        .Y(n4804) );
  MX4X1 U8374 ( .A(\registers[712][0] ), .B(\registers[713][0] ), .C(
        \registers[714][0] ), .D(\registers[715][0] ), .S0(n7453), .S1(n7696), 
        .Y(n4751) );
  MX4X1 U8375 ( .A(\registers[760][0] ), .B(\registers[761][0] ), .C(
        \registers[762][0] ), .D(\registers[763][0] ), .S0(n7452), .S1(n7695), 
        .Y(n4736) );
  MX4X1 U8376 ( .A(\registers[744][0] ), .B(\registers[745][0] ), .C(
        \registers[746][0] ), .D(\registers[747][0] ), .S0(n7453), .S1(n7695), 
        .Y(n4741) );
  MX4X1 U8377 ( .A(\registers[648][0] ), .B(\registers[649][0] ), .C(
        \registers[650][0] ), .D(\registers[651][0] ), .S0(n7455), .S1(n7697), 
        .Y(n4772) );
  MX4X1 U8378 ( .A(\registers[696][0] ), .B(\registers[697][0] ), .C(
        \registers[698][0] ), .D(\registers[699][0] ), .S0(n7454), .S1(n7696), 
        .Y(n4757) );
  MX4X1 U8379 ( .A(\registers[680][0] ), .B(\registers[681][0] ), .C(
        \registers[682][0] ), .D(\registers[683][0] ), .S0(n7454), .S1(n7697), 
        .Y(n4762) );
  MX4X1 U8380 ( .A(\registers[328][1] ), .B(\registers[329][1] ), .C(
        \registers[330][1] ), .D(\registers[331][1] ), .S0(n7483), .S1(n7723), 
        .Y(n5218) );
  MX4X1 U8381 ( .A(\registers[376][1] ), .B(\registers[377][1] ), .C(
        \registers[378][1] ), .D(\registers[379][1] ), .S0(n7482), .S1(n7722), 
        .Y(n5203) );
  MX4X1 U8382 ( .A(\registers[360][1] ), .B(\registers[361][1] ), .C(
        \registers[362][1] ), .D(\registers[363][1] ), .S0(n7482), .S1(n7722), 
        .Y(n5208) );
  MX4X1 U8383 ( .A(\registers[72][1] ), .B(\registers[73][1] ), .C(
        \registers[74][1] ), .D(\registers[75][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5303) );
  MX4X1 U8384 ( .A(\registers[120][1] ), .B(\registers[121][1] ), .C(
        \registers[122][1] ), .D(\registers[123][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5288) );
  MX4X1 U8385 ( .A(\registers[104][1] ), .B(\registers[105][1] ), .C(
        \registers[106][1] ), .D(\registers[107][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5293) );
  MX4X1 U8386 ( .A(\registers[8][1] ), .B(\registers[9][1] ), .C(
        \registers[10][1] ), .D(\registers[11][1] ), .S0(n7489), .S1(n7729), 
        .Y(n5324) );
  MX4X1 U8387 ( .A(\registers[56][1] ), .B(\registers[57][1] ), .C(
        \registers[58][1] ), .D(\registers[59][1] ), .S0(n7488), .S1(n7728), 
        .Y(n5309) );
  MX4X1 U8388 ( .A(\registers[40][1] ), .B(\registers[41][1] ), .C(
        \registers[42][1] ), .D(\registers[43][1] ), .S0(n7489), .S1(n7729), 
        .Y(n5314) );
  MX4X1 U8389 ( .A(\registers[200][1] ), .B(\registers[201][1] ), .C(
        \registers[202][1] ), .D(\registers[203][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5261) );
  MX4X1 U8390 ( .A(\registers[248][1] ), .B(\registers[249][1] ), .C(
        \registers[250][1] ), .D(\registers[251][1] ), .S0(n7484), .S1(n7725), 
        .Y(n5246) );
  MX4X1 U8391 ( .A(\registers[232][1] ), .B(\registers[233][1] ), .C(
        \registers[234][1] ), .D(\registers[235][1] ), .S0(n7485), .S1(n7725), 
        .Y(n5251) );
  MX4X1 U8392 ( .A(\registers[136][1] ), .B(\registers[137][1] ), .C(
        \registers[138][1] ), .D(\registers[139][1] ), .S0(n7487), .S1(n7727), 
        .Y(n5282) );
  MX4X1 U8393 ( .A(\registers[184][1] ), .B(\registers[185][1] ), .C(
        \registers[186][1] ), .D(\registers[187][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5267) );
  MX4X1 U8394 ( .A(\registers[168][1] ), .B(\registers[169][1] ), .C(
        \registers[170][1] ), .D(\registers[171][1] ), .S0(n7486), .S1(n7726), 
        .Y(n5272) );
  MX4X1 U8395 ( .A(\registers[840][1] ), .B(\registers[841][1] ), .C(
        \registers[842][1] ), .D(\registers[843][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5048) );
  MX4X1 U8396 ( .A(\registers[888][1] ), .B(\registers[889][1] ), .C(
        \registers[890][1] ), .D(\registers[891][1] ), .S0(n7471), .S1(n7712), 
        .Y(n5033) );
  MX4X1 U8397 ( .A(\registers[872][1] ), .B(\registers[873][1] ), .C(
        \registers[874][1] ), .D(\registers[875][1] ), .S0(n7471), .S1(n7713), 
        .Y(n5038) );
  MX4X1 U8398 ( .A(\registers[776][1] ), .B(\registers[777][1] ), .C(
        \registers[778][1] ), .D(\registers[779][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5069) );
  MX4X1 U8399 ( .A(\registers[824][1] ), .B(\registers[825][1] ), .C(
        \registers[826][1] ), .D(\registers[827][1] ), .S0(n7472), .S1(n7713), 
        .Y(n5054) );
  MX4X1 U8400 ( .A(\registers[808][1] ), .B(\registers[809][1] ), .C(
        \registers[810][1] ), .D(\registers[811][1] ), .S0(n7473), .S1(n7714), 
        .Y(n5059) );
  MX4X1 U8401 ( .A(\registers[968][1] ), .B(\registers[969][1] ), .C(
        \registers[970][1] ), .D(\registers[971][1] ), .S0(n7469), .S1(n7711), 
        .Y(n5006) );
  MX4X1 U8402 ( .A(\registers[1016][1] ), .B(\registers[1017][1] ), .C(
        \registers[1018][1] ), .D(\registers[1019][1] ), .S0(n7468), .S1(n7710), .Y(n4991) );
  MX4X1 U8403 ( .A(\registers[1000][1] ), .B(\registers[1001][1] ), .C(
        \registers[1002][1] ), .D(\registers[1003][1] ), .S0(n7469), .S1(n7710), .Y(n4996) );
  MX4X1 U8404 ( .A(\registers[904][1] ), .B(\registers[905][1] ), .C(
        \registers[906][1] ), .D(\registers[907][1] ), .S0(n7471), .S1(n7712), 
        .Y(n5027) );
  MX4X1 U8405 ( .A(\registers[952][1] ), .B(\registers[953][1] ), .C(
        \registers[954][1] ), .D(\registers[955][1] ), .S0(n7470), .S1(n7711), 
        .Y(n5012) );
  MX4X1 U8406 ( .A(\registers[936][1] ), .B(\registers[937][1] ), .C(
        \registers[938][1] ), .D(\registers[939][1] ), .S0(n7470), .S1(n7711), 
        .Y(n5017) );
  MX4X1 U8407 ( .A(\registers[584][1] ), .B(\registers[585][1] ), .C(
        \registers[586][1] ), .D(\registers[587][1] ), .S0(n7477), .S1(n7718), 
        .Y(n5133) );
  MX4X1 U8408 ( .A(\registers[632][1] ), .B(\registers[633][1] ), .C(
        \registers[634][1] ), .D(\registers[635][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5118) );
  MX4X1 U8409 ( .A(\registers[616][1] ), .B(\registers[617][1] ), .C(
        \registers[618][1] ), .D(\registers[619][1] ), .S0(n7477), .S1(n7717), 
        .Y(n5123) );
  MX4X1 U8410 ( .A(\registers[520][1] ), .B(\registers[521][1] ), .C(
        \registers[522][1] ), .D(\registers[523][1] ), .S0(n7479), .S1(n7719), 
        .Y(n5154) );
  MX4X1 U8411 ( .A(\registers[568][1] ), .B(\registers[569][1] ), .C(
        \registers[570][1] ), .D(\registers[571][1] ), .S0(n7478), .S1(n7718), 
        .Y(n5139) );
  MX4X1 U8412 ( .A(\registers[552][1] ), .B(\registers[553][1] ), .C(
        \registers[554][1] ), .D(\registers[555][1] ), .S0(n7478), .S1(n7719), 
        .Y(n5144) );
  MX4X1 U8413 ( .A(\registers[712][1] ), .B(\registers[713][1] ), .C(
        \registers[714][1] ), .D(\registers[715][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5091) );
  MX4X1 U8414 ( .A(\registers[760][1] ), .B(\registers[761][1] ), .C(
        \registers[762][1] ), .D(\registers[763][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5076) );
  MX4X1 U8415 ( .A(\registers[744][1] ), .B(\registers[745][1] ), .C(
        \registers[746][1] ), .D(\registers[747][1] ), .S0(n7474), .S1(n7715), 
        .Y(n5081) );
  MX4X1 U8416 ( .A(\registers[648][1] ), .B(\registers[649][1] ), .C(
        \registers[650][1] ), .D(\registers[651][1] ), .S0(n7476), .S1(n7717), 
        .Y(n5112) );
  MX4X1 U8417 ( .A(\registers[696][1] ), .B(\registers[697][1] ), .C(
        \registers[698][1] ), .D(\registers[699][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5097) );
  MX4X1 U8418 ( .A(\registers[680][1] ), .B(\registers[681][1] ), .C(
        \registers[682][1] ), .D(\registers[683][1] ), .S0(n7475), .S1(n7716), 
        .Y(n5102) );
  MX4X1 U8419 ( .A(\registers[328][2] ), .B(\registers[329][2] ), .C(
        \registers[330][2] ), .D(\registers[331][2] ), .S0(n7504), .S1(n7743), 
        .Y(n5558) );
  MX4X1 U8420 ( .A(\registers[376][2] ), .B(\registers[377][2] ), .C(
        \registers[378][2] ), .D(\registers[379][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5543) );
  MX4X1 U8421 ( .A(\registers[360][2] ), .B(\registers[361][2] ), .C(
        \registers[362][2] ), .D(\registers[363][2] ), .S0(n7503), .S1(n7742), 
        .Y(n5548) );
  MX4X1 U8422 ( .A(\registers[72][2] ), .B(\registers[73][2] ), .C(
        \registers[74][2] ), .D(\registers[75][2] ), .S0(n7509), .S1(n7748), 
        .Y(n5643) );
  MX4X1 U8423 ( .A(\registers[120][2] ), .B(\registers[121][2] ), .C(
        \registers[122][2] ), .D(\registers[123][2] ), .S0(n7508), .S1(n7747), 
        .Y(n5628) );
  MX4X1 U8424 ( .A(\registers[104][2] ), .B(\registers[105][2] ), .C(
        \registers[106][2] ), .D(\registers[107][2] ), .S0(n7509), .S1(n7747), 
        .Y(n5633) );
  MX4X1 U8425 ( .A(\registers[8][2] ), .B(\registers[9][2] ), .C(
        \registers[10][2] ), .D(\registers[11][2] ), .S0(n7511), .S1(n7749), 
        .Y(n5664) );
  MX4X1 U8426 ( .A(\registers[56][2] ), .B(\registers[57][2] ), .C(
        \registers[58][2] ), .D(\registers[59][2] ), .S0(n7510), .S1(n7748), 
        .Y(n5649) );
  MX4X1 U8427 ( .A(\registers[40][2] ), .B(\registers[41][2] ), .C(
        \registers[42][2] ), .D(\registers[43][2] ), .S0(n7510), .S1(n7748), 
        .Y(n5654) );
  MX4X1 U8428 ( .A(\registers[200][2] ), .B(\registers[201][2] ), .C(
        \registers[202][2] ), .D(\registers[203][2] ), .S0(n7507), .S1(n7745), 
        .Y(n5601) );
  MX4X1 U8429 ( .A(\registers[248][2] ), .B(\registers[249][2] ), .C(
        \registers[250][2] ), .D(\registers[251][2] ), .S0(n7506), .S1(n7744), 
        .Y(n5586) );
  MX4X1 U8430 ( .A(\registers[232][2] ), .B(\registers[233][2] ), .C(
        \registers[234][2] ), .D(\registers[235][2] ), .S0(n7506), .S1(n7745), 
        .Y(n5591) );
  MX4X1 U8431 ( .A(\registers[136][2] ), .B(\registers[137][2] ), .C(
        \registers[138][2] ), .D(\registers[139][2] ), .S0(n7508), .S1(n7746), 
        .Y(n5622) );
  MX4X1 U8432 ( .A(\registers[184][2] ), .B(\registers[185][2] ), .C(
        \registers[186][2] ), .D(\registers[187][2] ), .S0(n7507), .S1(n7745), 
        .Y(n5607) );
  MX4X1 U8433 ( .A(\registers[168][2] ), .B(\registers[169][2] ), .C(
        \registers[170][2] ), .D(\registers[171][2] ), .S0(n7507), .S1(n7746), 
        .Y(n5612) );
  MX4X1 U8434 ( .A(\registers[840][2] ), .B(\registers[841][2] ), .C(
        \registers[842][2] ), .D(\registers[843][2] ), .S0(n7493), .S1(n7733), 
        .Y(n5388) );
  MX4X1 U8435 ( .A(\registers[888][2] ), .B(\registers[889][2] ), .C(
        \registers[890][2] ), .D(\registers[891][2] ), .S0(n7492), .S1(n7732), 
        .Y(n5373) );
  MX4X1 U8436 ( .A(\registers[872][2] ), .B(\registers[873][2] ), .C(
        \registers[874][2] ), .D(\registers[875][2] ), .S0(n7493), .S1(n7732), 
        .Y(n5378) );
  MX4X1 U8437 ( .A(\registers[776][2] ), .B(\registers[777][2] ), .C(
        \registers[778][2] ), .D(\registers[779][2] ), .S0(n7495), .S1(n7734), 
        .Y(n5409) );
  MX4X1 U8438 ( .A(\registers[824][2] ), .B(\registers[825][2] ), .C(
        \registers[826][2] ), .D(\registers[827][2] ), .S0(n7494), .S1(n7733), 
        .Y(n5394) );
  MX4X1 U8439 ( .A(\registers[808][2] ), .B(\registers[809][2] ), .C(
        \registers[810][2] ), .D(\registers[811][2] ), .S0(n7494), .S1(n7733), 
        .Y(n5399) );
  MX4X1 U8440 ( .A(\registers[968][2] ), .B(\registers[969][2] ), .C(
        \registers[970][2] ), .D(\registers[971][2] ), .S0(n7491), .S1(n7730), 
        .Y(n5346) );
  MX4X1 U8441 ( .A(\registers[1016][2] ), .B(\registers[1017][2] ), .C(
        \registers[1018][2] ), .D(\registers[1019][2] ), .S0(n7490), .S1(n7729), .Y(n5331) );
  MX4X1 U8442 ( .A(\registers[1000][2] ), .B(\registers[1001][2] ), .C(
        \registers[1002][2] ), .D(\registers[1003][2] ), .S0(n7490), .S1(n7730), .Y(n5336) );
  MX4X1 U8443 ( .A(\registers[904][2] ), .B(\registers[905][2] ), .C(
        \registers[906][2] ), .D(\registers[907][2] ), .S0(n7492), .S1(n7732), 
        .Y(n5367) );
  MX4X1 U8444 ( .A(\registers[952][2] ), .B(\registers[953][2] ), .C(
        \registers[954][2] ), .D(\registers[955][2] ), .S0(n7491), .S1(n7731), 
        .Y(n5352) );
  MX4X1 U8445 ( .A(\registers[936][2] ), .B(\registers[937][2] ), .C(
        \registers[938][2] ), .D(\registers[939][2] ), .S0(n7491), .S1(n7731), 
        .Y(n5357) );
  MX4X1 U8446 ( .A(\registers[584][2] ), .B(\registers[585][2] ), .C(
        \registers[586][2] ), .D(\registers[587][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5473) );
  MX4X1 U8447 ( .A(\registers[632][2] ), .B(\registers[633][2] ), .C(
        \registers[634][2] ), .D(\registers[635][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5458) );
  MX4X1 U8448 ( .A(\registers[616][2] ), .B(\registers[617][2] ), .C(
        \registers[618][2] ), .D(\registers[619][2] ), .S0(n7498), .S1(n7737), 
        .Y(n5463) );
  MX4X1 U8449 ( .A(\registers[520][2] ), .B(\registers[521][2] ), .C(
        \registers[522][2] ), .D(\registers[523][2] ), .S0(n7500), .S1(n7739), 
        .Y(n5494) );
  MX4X1 U8450 ( .A(\registers[568][2] ), .B(\registers[569][2] ), .C(
        \registers[570][2] ), .D(\registers[571][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5479) );
  MX4X1 U8451 ( .A(\registers[552][2] ), .B(\registers[553][2] ), .C(
        \registers[554][2] ), .D(\registers[555][2] ), .S0(n7499), .S1(n7738), 
        .Y(n5484) );
  MX4X1 U8452 ( .A(\registers[712][2] ), .B(\registers[713][2] ), .C(
        \registers[714][2] ), .D(\registers[715][2] ), .S0(n7496), .S1(n7735), 
        .Y(n5431) );
  MX4X1 U8453 ( .A(\registers[760][2] ), .B(\registers[761][2] ), .C(
        \registers[762][2] ), .D(\registers[763][2] ), .S0(n7495), .S1(n7734), 
        .Y(n5416) );
  MX4X1 U8454 ( .A(\registers[744][2] ), .B(\registers[745][2] ), .C(
        \registers[746][2] ), .D(\registers[747][2] ), .S0(n7495), .S1(n7735), 
        .Y(n5421) );
  MX4X1 U8455 ( .A(\registers[648][2] ), .B(\registers[649][2] ), .C(
        \registers[650][2] ), .D(\registers[651][2] ), .S0(n7497), .S1(n7737), 
        .Y(n5452) );
  MX4X1 U8456 ( .A(\registers[696][2] ), .B(\registers[697][2] ), .C(
        \registers[698][2] ), .D(\registers[699][2] ), .S0(n7496), .S1(n7736), 
        .Y(n5437) );
  MX4X1 U8457 ( .A(\registers[680][2] ), .B(\registers[681][2] ), .C(
        \registers[682][2] ), .D(\registers[683][2] ), .S0(n7497), .S1(n7736), 
        .Y(n5442) );
  MX4X1 U8458 ( .A(\registers[328][3] ), .B(\registers[329][3] ), .C(
        \registers[330][3] ), .D(\registers[331][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5898) );
  MX4X1 U8459 ( .A(\registers[376][3] ), .B(\registers[377][3] ), .C(
        \registers[378][3] ), .D(\registers[379][3] ), .S0(n7524), .S1(n7761), 
        .Y(n5883) );
  MX4X1 U8460 ( .A(\registers[360][3] ), .B(\registers[361][3] ), .C(
        \registers[362][3] ), .D(\registers[363][3] ), .S0(n7525), .S1(n7762), 
        .Y(n5888) );
  MX4X1 U8461 ( .A(\registers[72][3] ), .B(\registers[73][3] ), .C(
        \registers[74][3] ), .D(\registers[75][3] ), .S0(n7531), .S1(n7767), 
        .Y(n5983) );
  MX4X1 U8462 ( .A(\registers[120][3] ), .B(\registers[121][3] ), .C(
        \registers[122][3] ), .D(\registers[123][3] ), .S0(n7530), .S1(n7766), 
        .Y(n5968) );
  MX4X1 U8463 ( .A(\registers[104][3] ), .B(\registers[105][3] ), .C(
        \registers[106][3] ), .D(\registers[107][3] ), .S0(n7530), .S1(n7767), 
        .Y(n5973) );
  MX4X1 U8464 ( .A(\registers[8][3] ), .B(\registers[9][3] ), .C(
        \registers[10][3] ), .D(\registers[11][3] ), .S0(n7532), .S1(n7769), 
        .Y(n6004) );
  MX4X1 U8465 ( .A(\registers[56][3] ), .B(\registers[57][3] ), .C(
        \registers[58][3] ), .D(\registers[59][3] ), .S0(n7531), .S1(n7768), 
        .Y(n5989) );
  MX4X1 U8466 ( .A(\registers[40][3] ), .B(\registers[41][3] ), .C(
        \registers[42][3] ), .D(\registers[43][3] ), .S0(n7531), .S1(n7768), 
        .Y(n5994) );
  MX4X1 U8467 ( .A(\registers[200][3] ), .B(\registers[201][3] ), .C(
        \registers[202][3] ), .D(\registers[203][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5941) );
  MX4X1 U8468 ( .A(\registers[248][3] ), .B(\registers[249][3] ), .C(
        \registers[250][3] ), .D(\registers[251][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5926) );
  MX4X1 U8469 ( .A(\registers[232][3] ), .B(\registers[233][3] ), .C(
        \registers[234][3] ), .D(\registers[235][3] ), .S0(n7527), .S1(n7764), 
        .Y(n5931) );
  MX4X1 U8470 ( .A(\registers[136][3] ), .B(\registers[137][3] ), .C(
        \registers[138][3] ), .D(\registers[139][3] ), .S0(n7529), .S1(n7766), 
        .Y(n5962) );
  MX4X1 U8471 ( .A(\registers[184][3] ), .B(\registers[185][3] ), .C(
        \registers[186][3] ), .D(\registers[187][3] ), .S0(n7528), .S1(n7765), 
        .Y(n5947) );
  MX4X1 U8472 ( .A(\registers[168][3] ), .B(\registers[169][3] ), .C(
        \registers[170][3] ), .D(\registers[171][3] ), .S0(n7529), .S1(n7765), 
        .Y(n5952) );
  MX4X1 U8473 ( .A(\registers[840][3] ), .B(\registers[841][3] ), .C(
        \registers[842][3] ), .D(\registers[843][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5728) );
  MX4X1 U8474 ( .A(\registers[888][3] ), .B(\registers[889][3] ), .C(
        \registers[890][3] ), .D(\registers[891][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5713) );
  MX4X1 U8475 ( .A(\registers[872][3] ), .B(\registers[873][3] ), .C(
        \registers[874][3] ), .D(\registers[875][3] ), .S0(n7514), .S1(n7752), 
        .Y(n5718) );
  MX4X1 U8476 ( .A(\registers[776][3] ), .B(\registers[777][3] ), .C(
        \registers[778][3] ), .D(\registers[779][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5749) );
  MX4X1 U8477 ( .A(\registers[824][3] ), .B(\registers[825][3] ), .C(
        \registers[826][3] ), .D(\registers[827][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5734) );
  MX4X1 U8478 ( .A(\registers[808][3] ), .B(\registers[809][3] ), .C(
        \registers[810][3] ), .D(\registers[811][3] ), .S0(n7515), .S1(n7753), 
        .Y(n5739) );
  MX4X1 U8479 ( .A(\registers[968][3] ), .B(\registers[969][3] ), .C(
        \registers[970][3] ), .D(\registers[971][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5686) );
  MX4X1 U8480 ( .A(\registers[1016][3] ), .B(\registers[1017][3] ), .C(
        \registers[1018][3] ), .D(\registers[1019][3] ), .S0(n7511), .S1(n7749), .Y(n5671) );
  MX4X1 U8481 ( .A(\registers[1000][3] ), .B(\registers[1001][3] ), .C(
        \registers[1002][3] ), .D(\registers[1003][3] ), .S0(n7511), .S1(n7749), .Y(n5676) );
  MX4X1 U8482 ( .A(\registers[904][3] ), .B(\registers[905][3] ), .C(
        \registers[906][3] ), .D(\registers[907][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5707) );
  MX4X1 U8483 ( .A(\registers[952][3] ), .B(\registers[953][3] ), .C(
        \registers[954][3] ), .D(\registers[955][3] ), .S0(n7512), .S1(n7750), 
        .Y(n5692) );
  MX4X1 U8484 ( .A(\registers[936][3] ), .B(\registers[937][3] ), .C(
        \registers[938][3] ), .D(\registers[939][3] ), .S0(n7513), .S1(n7751), 
        .Y(n5697) );
  MX4X1 U8485 ( .A(\registers[584][3] ), .B(\registers[585][3] ), .C(
        \registers[586][3] ), .D(\registers[587][3] ), .S0(n7520), .S1(n7757), 
        .Y(n5813) );
  MX4X1 U8486 ( .A(\registers[632][3] ), .B(\registers[633][3] ), .C(
        \registers[634][3] ), .D(\registers[635][3] ), .S0(n7519), .S1(n7757), 
        .Y(n5798) );
  MX4X1 U8487 ( .A(\registers[616][3] ), .B(\registers[617][3] ), .C(
        \registers[618][3] ), .D(\registers[619][3] ), .S0(n7519), .S1(n7757), 
        .Y(n5803) );
  MX4X1 U8488 ( .A(\registers[520][3] ), .B(\registers[521][3] ), .C(
        \registers[522][3] ), .D(\registers[523][3] ), .S0(n7521), .S1(n7759), 
        .Y(n5834) );
  MX4X1 U8489 ( .A(\registers[568][3] ), .B(\registers[569][3] ), .C(
        \registers[570][3] ), .D(\registers[571][3] ), .S0(n7520), .S1(n7758), 
        .Y(n5819) );
  MX4X1 U8490 ( .A(\registers[552][3] ), .B(\registers[553][3] ), .C(
        \registers[554][3] ), .D(\registers[555][3] ), .S0(n7521), .S1(n7758), 
        .Y(n5824) );
  MX4X1 U8491 ( .A(\registers[712][3] ), .B(\registers[713][3] ), .C(
        \registers[714][3] ), .D(\registers[715][3] ), .S0(n7517), .S1(n7755), 
        .Y(n5771) );
  MX4X1 U8492 ( .A(\registers[760][3] ), .B(\registers[761][3] ), .C(
        \registers[762][3] ), .D(\registers[763][3] ), .S0(n7516), .S1(n7754), 
        .Y(n5756) );
  MX4X1 U8493 ( .A(\registers[744][3] ), .B(\registers[745][3] ), .C(
        \registers[746][3] ), .D(\registers[747][3] ), .S0(n7517), .S1(n7754), 
        .Y(n5761) );
  MX4X1 U8494 ( .A(\registers[648][3] ), .B(\registers[649][3] ), .C(
        \registers[650][3] ), .D(\registers[651][3] ), .S0(n7519), .S1(n7756), 
        .Y(n5792) );
  MX4X1 U8495 ( .A(\registers[696][3] ), .B(\registers[697][3] ), .C(
        \registers[698][3] ), .D(\registers[699][3] ), .S0(n7518), .S1(n7755), 
        .Y(n5777) );
  MX4X1 U8496 ( .A(\registers[680][3] ), .B(\registers[681][3] ), .C(
        \registers[682][3] ), .D(\registers[683][3] ), .S0(n7518), .S1(n7756), 
        .Y(n5782) );
  MX4X1 U8497 ( .A(\registers[328][4] ), .B(\registers[329][4] ), .C(
        \registers[330][4] ), .D(\registers[331][4] ), .S0(n7547), .S1(n7782), 
        .Y(n6238) );
  MX4X1 U8498 ( .A(\registers[376][4] ), .B(\registers[377][4] ), .C(
        \registers[378][4] ), .D(\registers[379][4] ), .S0(n7546), .S1(n7781), 
        .Y(n6223) );
  MX4X1 U8499 ( .A(\registers[360][4] ), .B(\registers[361][4] ), .C(
        \registers[362][4] ), .D(\registers[363][4] ), .S0(n7546), .S1(n7781), 
        .Y(n6228) );
  MX4X1 U8500 ( .A(\registers[72][4] ), .B(\registers[73][4] ), .C(
        \registers[74][4] ), .D(\registers[75][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6323) );
  MX4X1 U8501 ( .A(\registers[120][4] ), .B(\registers[121][4] ), .C(
        \registers[122][4] ), .D(\registers[123][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6308) );
  MX4X1 U8502 ( .A(\registers[104][4] ), .B(\registers[105][4] ), .C(
        \registers[106][4] ), .D(\registers[107][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6313) );
  MX4X1 U8503 ( .A(\registers[8][4] ), .B(\registers[9][4] ), .C(
        \registers[10][4] ), .D(\registers[11][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6344) );
  MX4X1 U8504 ( .A(\registers[56][4] ), .B(\registers[57][4] ), .C(
        \registers[58][4] ), .D(\registers[59][4] ), .S0(n7552), .S1(n7787), 
        .Y(n6329) );
  MX4X1 U8505 ( .A(\registers[40][4] ), .B(\registers[41][4] ), .C(
        \registers[42][4] ), .D(\registers[43][4] ), .S0(n7553), .S1(n7788), 
        .Y(n6334) );
  MX4X1 U8506 ( .A(\registers[200][4] ), .B(\registers[201][4] ), .C(
        \registers[202][4] ), .D(\registers[203][4] ), .S0(n7549), .S1(n7785), 
        .Y(n6281) );
  MX4X1 U8507 ( .A(\registers[248][4] ), .B(\registers[249][4] ), .C(
        \registers[250][4] ), .D(\registers[251][4] ), .S0(n7548), .S1(n7784), 
        .Y(n6266) );
  MX4X1 U8508 ( .A(\registers[232][4] ), .B(\registers[233][4] ), .C(
        \registers[234][4] ), .D(\registers[235][4] ), .S0(n7549), .S1(n7784), 
        .Y(n6271) );
  MX4X1 U8509 ( .A(\registers[136][4] ), .B(\registers[137][4] ), .C(
        \registers[138][4] ), .D(\registers[139][4] ), .S0(n7551), .S1(n7786), 
        .Y(n6302) );
  MX4X1 U8510 ( .A(\registers[184][4] ), .B(\registers[185][4] ), .C(
        \registers[186][4] ), .D(\registers[187][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6287) );
  MX4X1 U8511 ( .A(\registers[168][4] ), .B(\registers[169][4] ), .C(
        \registers[170][4] ), .D(\registers[171][4] ), .S0(n7550), .S1(n7785), 
        .Y(n6292) );
  MX4X1 U8512 ( .A(\registers[840][4] ), .B(\registers[841][4] ), .C(
        \registers[842][4] ), .D(\registers[843][4] ), .S0(n7536), .S1(n7772), 
        .Y(n6068) );
  MX4X1 U8513 ( .A(\registers[888][4] ), .B(\registers[889][4] ), .C(
        \registers[890][4] ), .D(\registers[891][4] ), .S0(n7535), .S1(n7771), 
        .Y(n6053) );
  MX4X1 U8514 ( .A(\registers[872][4] ), .B(\registers[873][4] ), .C(
        \registers[874][4] ), .D(\registers[875][4] ), .S0(n7535), .S1(n7772), 
        .Y(n6058) );
  MX4X1 U8515 ( .A(\registers[776][4] ), .B(\registers[777][4] ), .C(
        \registers[778][4] ), .D(\registers[779][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6089) );
  MX4X1 U8516 ( .A(\registers[824][4] ), .B(\registers[825][4] ), .C(
        \registers[826][4] ), .D(\registers[827][4] ), .S0(n7536), .S1(n7773), 
        .Y(n6074) );
  MX4X1 U8517 ( .A(\registers[808][4] ), .B(\registers[809][4] ), .C(
        \registers[810][4] ), .D(\registers[811][4] ), .S0(n7537), .S1(n7773), 
        .Y(n6079) );
  MX4X1 U8518 ( .A(\registers[968][4] ), .B(\registers[969][4] ), .C(
        \registers[970][4] ), .D(\registers[971][4] ), .S0(n7533), .S1(n7770), 
        .Y(n6026) );
  MX4X1 U8519 ( .A(\registers[1016][4] ), .B(\registers[1017][4] ), .C(
        \registers[1018][4] ), .D(\registers[1019][4] ), .S0(n7532), .S1(n7769), .Y(n6011) );
  MX4X1 U8520 ( .A(\registers[1000][4] ), .B(\registers[1001][4] ), .C(
        \registers[1002][4] ), .D(\registers[1003][4] ), .S0(n7533), .S1(n7769), .Y(n6016) );
  MX4X1 U8521 ( .A(\registers[904][4] ), .B(\registers[905][4] ), .C(
        \registers[906][4] ), .D(\registers[907][4] ), .S0(n7535), .S1(n7771), 
        .Y(n6047) );
  MX4X1 U8522 ( .A(\registers[952][4] ), .B(\registers[953][4] ), .C(
        \registers[954][4] ), .D(\registers[955][4] ), .S0(n7534), .S1(n7770), 
        .Y(n6032) );
  MX4X1 U8523 ( .A(\registers[936][4] ), .B(\registers[937][4] ), .C(
        \registers[938][4] ), .D(\registers[939][4] ), .S0(n7534), .S1(n7770), 
        .Y(n6037) );
  MX4X1 U8524 ( .A(\registers[584][4] ), .B(\registers[585][4] ), .C(
        \registers[586][4] ), .D(\registers[587][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6153) );
  MX4X1 U8525 ( .A(\registers[632][4] ), .B(\registers[633][4] ), .C(
        \registers[634][4] ), .D(\registers[635][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6138) );
  MX4X1 U8526 ( .A(\registers[616][4] ), .B(\registers[617][4] ), .C(
        \registers[618][4] ), .D(\registers[619][4] ), .S0(n7541), .S1(n7777), 
        .Y(n6143) );
  MX4X1 U8527 ( .A(\registers[520][4] ), .B(\registers[521][4] ), .C(
        \registers[522][4] ), .D(\registers[523][4] ), .S0(n7543), .S1(n7778), 
        .Y(n6174) );
  MX4X1 U8528 ( .A(\registers[568][4] ), .B(\registers[569][4] ), .C(
        \registers[570][4] ), .D(\registers[571][4] ), .S0(n7542), .S1(n7777), 
        .Y(n6159) );
  MX4X1 U8529 ( .A(\registers[552][4] ), .B(\registers[553][4] ), .C(
        \registers[554][4] ), .D(\registers[555][4] ), .S0(n7542), .S1(n7778), 
        .Y(n6164) );
  MX4X1 U8530 ( .A(\registers[712][4] ), .B(\registers[713][4] ), .C(
        \registers[714][4] ), .D(\registers[715][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6111) );
  MX4X1 U8531 ( .A(\registers[760][4] ), .B(\registers[761][4] ), .C(
        \registers[762][4] ), .D(\registers[763][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6096) );
  MX4X1 U8532 ( .A(\registers[744][4] ), .B(\registers[745][4] ), .C(
        \registers[746][4] ), .D(\registers[747][4] ), .S0(n7538), .S1(n7774), 
        .Y(n6101) );
  MX4X1 U8533 ( .A(\registers[648][4] ), .B(\registers[649][4] ), .C(
        \registers[650][4] ), .D(\registers[651][4] ), .S0(n7540), .S1(n7776), 
        .Y(n6132) );
  MX4X1 U8534 ( .A(\registers[696][4] ), .B(\registers[697][4] ), .C(
        \registers[698][4] ), .D(\registers[699][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6117) );
  MX4X1 U8535 ( .A(\registers[680][4] ), .B(\registers[681][4] ), .C(
        \registers[682][4] ), .D(\registers[683][4] ), .S0(n7539), .S1(n7775), 
        .Y(n6122) );
  MX4X1 U8536 ( .A(\registers[328][5] ), .B(\registers[329][5] ), .C(
        \registers[330][5] ), .D(\registers[331][5] ), .S0(n7568), .S1(n7802), 
        .Y(n6578) );
  MX4X1 U8537 ( .A(\registers[376][5] ), .B(\registers[377][5] ), .C(
        \registers[378][5] ), .D(\registers[379][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6563) );
  MX4X1 U8538 ( .A(\registers[360][5] ), .B(\registers[361][5] ), .C(
        \registers[362][5] ), .D(\registers[363][5] ), .S0(n7567), .S1(n7801), 
        .Y(n6568) );
  MX4X1 U8539 ( .A(\registers[72][5] ), .B(\registers[73][5] ), .C(
        \registers[74][5] ), .D(\registers[75][5] ), .S0(n7573), .S1(n7806), 
        .Y(n6663) );
  MX4X1 U8540 ( .A(\registers[120][5] ), .B(\registers[121][5] ), .C(
        \registers[122][5] ), .D(\registers[123][5] ), .S0(n7572), .S1(n7805), 
        .Y(n6648) );
  MX4X1 U8541 ( .A(\registers[104][5] ), .B(\registers[105][5] ), .C(
        \registers[106][5] ), .D(\registers[107][5] ), .S0(n7573), .S1(n7805), 
        .Y(n6653) );
  MX4X1 U8542 ( .A(\registers[8][5] ), .B(\registers[9][5] ), .C(
        \registers[10][5] ), .D(\registers[11][5] ), .S0(n7575), .S1(n7807), 
        .Y(n6684) );
  MX4X1 U8543 ( .A(\registers[56][5] ), .B(\registers[57][5] ), .C(
        \registers[58][5] ), .D(\registers[59][5] ), .S0(n7574), .S1(n7806), 
        .Y(n6669) );
  MX4X1 U8544 ( .A(\registers[40][5] ), .B(\registers[41][5] ), .C(
        \registers[42][5] ), .D(\registers[43][5] ), .S0(n7574), .S1(n7806), 
        .Y(n6674) );
  MX4X1 U8545 ( .A(\registers[200][5] ), .B(\registers[201][5] ), .C(
        \registers[202][5] ), .D(\registers[203][5] ), .S0(n7571), .S1(n7831), 
        .Y(n6621) );
  MX4X1 U8546 ( .A(\registers[248][5] ), .B(\registers[249][5] ), .C(
        \registers[250][5] ), .D(\registers[251][5] ), .S0(n7570), .S1(n7803), 
        .Y(n6606) );
  MX4X1 U8547 ( .A(\registers[232][5] ), .B(\registers[233][5] ), .C(
        \registers[234][5] ), .D(\registers[235][5] ), .S0(n7570), .S1(n7822), 
        .Y(n6611) );
  MX4X1 U8548 ( .A(\registers[136][5] ), .B(\registers[137][5] ), .C(
        \registers[138][5] ), .D(\registers[139][5] ), .S0(n7572), .S1(n7804), 
        .Y(n6642) );
  MX4X1 U8549 ( .A(\registers[184][5] ), .B(\registers[185][5] ), .C(
        \registers[186][5] ), .D(\registers[187][5] ), .S0(n7571), .S1(n7804), 
        .Y(n6627) );
  MX4X1 U8550 ( .A(\registers[168][5] ), .B(\registers[169][5] ), .C(
        \registers[170][5] ), .D(\registers[171][5] ), .S0(n7571), .S1(n7804), 
        .Y(n6632) );
  MX4X1 U8551 ( .A(\registers[840][5] ), .B(\registers[841][5] ), .C(
        \registers[842][5] ), .D(\registers[843][5] ), .S0(n7557), .S1(n7792), 
        .Y(n6408) );
  MX4X1 U8552 ( .A(\registers[888][5] ), .B(\registers[889][5] ), .C(
        \registers[890][5] ), .D(\registers[891][5] ), .S0(n7556), .S1(n7791), 
        .Y(n6393) );
  MX4X1 U8553 ( .A(\registers[872][5] ), .B(\registers[873][5] ), .C(
        \registers[874][5] ), .D(\registers[875][5] ), .S0(n7557), .S1(n7791), 
        .Y(n6398) );
  MX4X1 U8554 ( .A(\registers[776][5] ), .B(\registers[777][5] ), .C(
        \registers[778][5] ), .D(\registers[779][5] ), .S0(n7559), .S1(n7793), 
        .Y(n6429) );
  MX4X1 U8555 ( .A(\registers[824][5] ), .B(\registers[825][5] ), .C(
        \registers[826][5] ), .D(\registers[827][5] ), .S0(n7558), .S1(n7792), 
        .Y(n6414) );
  MX4X1 U8556 ( .A(\registers[808][5] ), .B(\registers[809][5] ), .C(
        \registers[810][5] ), .D(\registers[811][5] ), .S0(n7558), .S1(n7793), 
        .Y(n6419) );
  MX4X1 U8557 ( .A(\registers[968][5] ), .B(\registers[969][5] ), .C(
        \registers[970][5] ), .D(\registers[971][5] ), .S0(n7555), .S1(n7789), 
        .Y(n6366) );
  MX4X1 U8558 ( .A(\registers[1016][5] ), .B(\registers[1017][5] ), .C(
        \registers[1018][5] ), .D(\registers[1019][5] ), .S0(n7554), .S1(n7789), .Y(n6351) );
  MX4X1 U8559 ( .A(\registers[1000][5] ), .B(\registers[1001][5] ), .C(
        \registers[1002][5] ), .D(\registers[1003][5] ), .S0(n7554), .S1(n7789), .Y(n6356) );
  MX4X1 U8560 ( .A(\registers[904][5] ), .B(\registers[905][5] ), .C(
        \registers[906][5] ), .D(\registers[907][5] ), .S0(n7556), .S1(n7791), 
        .Y(n6387) );
  MX4X1 U8561 ( .A(\registers[952][5] ), .B(\registers[953][5] ), .C(
        \registers[954][5] ), .D(\registers[955][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6372) );
  MX4X1 U8562 ( .A(\registers[936][5] ), .B(\registers[937][5] ), .C(
        \registers[938][5] ), .D(\registers[939][5] ), .S0(n7555), .S1(n7790), 
        .Y(n6377) );
  MX4X1 U8563 ( .A(\registers[584][5] ), .B(\registers[585][5] ), .C(
        \registers[586][5] ), .D(\registers[587][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6493) );
  MX4X1 U8564 ( .A(\registers[632][5] ), .B(\registers[633][5] ), .C(
        \registers[634][5] ), .D(\registers[635][5] ), .S0(n7562), .S1(n7796), 
        .Y(n6478) );
  MX4X1 U8565 ( .A(\registers[616][5] ), .B(\registers[617][5] ), .C(
        \registers[618][5] ), .D(\registers[619][5] ), .S0(n7562), .S1(n7796), 
        .Y(n6483) );
  MX4X1 U8566 ( .A(\registers[520][5] ), .B(\registers[521][5] ), .C(
        \registers[522][5] ), .D(\registers[523][5] ), .S0(n7564), .S1(n7798), 
        .Y(n6514) );
  MX4X1 U8567 ( .A(\registers[568][5] ), .B(\registers[569][5] ), .C(
        \registers[570][5] ), .D(\registers[571][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6499) );
  MX4X1 U8568 ( .A(\registers[552][5] ), .B(\registers[553][5] ), .C(
        \registers[554][5] ), .D(\registers[555][5] ), .S0(n7563), .S1(n7797), 
        .Y(n6504) );
  MX4X1 U8569 ( .A(\registers[712][5] ), .B(\registers[713][5] ), .C(
        \registers[714][5] ), .D(\registers[715][5] ), .S0(n7560), .S1(n7794), 
        .Y(n6451) );
  MX4X1 U8570 ( .A(\registers[760][5] ), .B(\registers[761][5] ), .C(
        \registers[762][5] ), .D(\registers[763][5] ), .S0(n7559), .S1(n7793), 
        .Y(n6436) );
  MX4X1 U8571 ( .A(\registers[744][5] ), .B(\registers[745][5] ), .C(
        \registers[746][5] ), .D(\registers[747][5] ), .S0(n7559), .S1(n7794), 
        .Y(n6441) );
  MX4X1 U8572 ( .A(\registers[648][5] ), .B(\registers[649][5] ), .C(
        \registers[650][5] ), .D(\registers[651][5] ), .S0(n7561), .S1(n7796), 
        .Y(n6472) );
  MX4X1 U8573 ( .A(\registers[696][5] ), .B(\registers[697][5] ), .C(
        \registers[698][5] ), .D(\registers[699][5] ), .S0(n7560), .S1(n7795), 
        .Y(n6457) );
  MX4X1 U8574 ( .A(\registers[680][5] ), .B(\registers[681][5] ), .C(
        \registers[682][5] ), .D(\registers[683][5] ), .S0(n7561), .S1(n7795), 
        .Y(n6462) );
  MX4X1 U8575 ( .A(\registers[328][6] ), .B(\registers[329][6] ), .C(
        \registers[330][6] ), .D(\registers[331][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6918) );
  MX4X1 U8576 ( .A(\registers[376][6] ), .B(\registers[377][6] ), .C(
        \registers[378][6] ), .D(\registers[379][6] ), .S0(n7588), .S1(n7820), 
        .Y(n6903) );
  MX4X1 U8577 ( .A(\registers[360][6] ), .B(\registers[361][6] ), .C(
        \registers[362][6] ), .D(\registers[363][6] ), .S0(n7589), .S1(n7820), 
        .Y(n6908) );
  MX4X1 U8578 ( .A(\registers[72][6] ), .B(\registers[73][6] ), .C(
        \registers[74][6] ), .D(\registers[75][6] ), .S0(n7595), .S1(n7825), 
        .Y(n7003) );
  MX4X1 U8579 ( .A(\registers[120][6] ), .B(\registers[121][6] ), .C(
        \registers[122][6] ), .D(\registers[123][6] ), .S0(n7594), .S1(n7824), 
        .Y(n6988) );
  MX4X1 U8580 ( .A(\registers[104][6] ), .B(\registers[105][6] ), .C(
        \registers[106][6] ), .D(\registers[107][6] ), .S0(n7594), .S1(n7825), 
        .Y(n6993) );
  MX4X1 U8581 ( .A(\registers[8][6] ), .B(\registers[9][6] ), .C(
        \registers[10][6] ), .D(\registers[11][6] ), .S0(n7596), .S1(n7827), 
        .Y(n7024) );
  MX4X1 U8582 ( .A(\registers[56][6] ), .B(\registers[57][6] ), .C(
        \registers[58][6] ), .D(\registers[59][6] ), .S0(n7595), .S1(n7826), 
        .Y(n7009) );
  MX4X1 U8583 ( .A(\registers[40][6] ), .B(\registers[41][6] ), .C(
        \registers[42][6] ), .D(\registers[43][6] ), .S0(n7595), .S1(n7826), 
        .Y(n7014) );
  MX4X1 U8584 ( .A(\registers[200][6] ), .B(\registers[201][6] ), .C(
        \registers[202][6] ), .D(\registers[203][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6961) );
  MX4X1 U8585 ( .A(\registers[248][6] ), .B(\registers[249][6] ), .C(
        \registers[250][6] ), .D(\registers[251][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6946) );
  MX4X1 U8586 ( .A(\registers[232][6] ), .B(\registers[233][6] ), .C(
        \registers[234][6] ), .D(\registers[235][6] ), .S0(n7591), .S1(n7822), 
        .Y(n6951) );
  MX4X1 U8587 ( .A(\registers[136][6] ), .B(\registers[137][6] ), .C(
        \registers[138][6] ), .D(\registers[139][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6982) );
  MX4X1 U8588 ( .A(\registers[184][6] ), .B(\registers[185][6] ), .C(
        \registers[186][6] ), .D(\registers[187][6] ), .S0(n7592), .S1(n7823), 
        .Y(n6967) );
  MX4X1 U8589 ( .A(\registers[168][6] ), .B(\registers[169][6] ), .C(
        \registers[170][6] ), .D(\registers[171][6] ), .S0(n7593), .S1(n7824), 
        .Y(n6972) );
  MX4X1 U8590 ( .A(\registers[840][6] ), .B(\registers[841][6] ), .C(
        \registers[842][6] ), .D(\registers[843][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6748) );
  MX4X1 U8591 ( .A(\registers[888][6] ), .B(\registers[889][6] ), .C(
        \registers[890][6] ), .D(\registers[891][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6733) );
  MX4X1 U8592 ( .A(\registers[872][6] ), .B(\registers[873][6] ), .C(
        \registers[874][6] ), .D(\registers[875][6] ), .S0(n7578), .S1(n7810), 
        .Y(n6738) );
  MX4X1 U8593 ( .A(\registers[776][6] ), .B(\registers[777][6] ), .C(
        \registers[778][6] ), .D(\registers[779][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6769) );
  MX4X1 U8594 ( .A(\registers[824][6] ), .B(\registers[825][6] ), .C(
        \registers[826][6] ), .D(\registers[827][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6754) );
  MX4X1 U8595 ( .A(\registers[808][6] ), .B(\registers[809][6] ), .C(
        \registers[810][6] ), .D(\registers[811][6] ), .S0(n7579), .S1(n7811), 
        .Y(n6759) );
  MX4X1 U8596 ( .A(\registers[968][6] ), .B(\registers[969][6] ), .C(
        \registers[970][6] ), .D(\registers[971][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6706) );
  MX4X1 U8597 ( .A(\registers[1016][6] ), .B(\registers[1017][6] ), .C(
        \registers[1018][6] ), .D(\registers[1019][6] ), .S0(n7575), .S1(n7807), .Y(n6691) );
  MX4X1 U8598 ( .A(\registers[1000][6] ), .B(\registers[1001][6] ), .C(
        \registers[1002][6] ), .D(\registers[1003][6] ), .S0(n7575), .S1(n7808), .Y(n6696) );
  MX4X1 U8599 ( .A(\registers[904][6] ), .B(\registers[905][6] ), .C(
        \registers[906][6] ), .D(\registers[907][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6727) );
  MX4X1 U8600 ( .A(\registers[952][6] ), .B(\registers[953][6] ), .C(
        \registers[954][6] ), .D(\registers[955][6] ), .S0(n7576), .S1(n7808), 
        .Y(n6712) );
  MX4X1 U8601 ( .A(\registers[936][6] ), .B(\registers[937][6] ), .C(
        \registers[938][6] ), .D(\registers[939][6] ), .S0(n7577), .S1(n7809), 
        .Y(n6717) );
  MX4X1 U8602 ( .A(\registers[584][6] ), .B(\registers[585][6] ), .C(
        \registers[586][6] ), .D(\registers[587][6] ), .S0(n7584), .S1(n7816), 
        .Y(n6833) );
  MX4X1 U8603 ( .A(\registers[632][6] ), .B(\registers[633][6] ), .C(
        \registers[634][6] ), .D(\registers[635][6] ), .S0(n7583), .S1(n7815), 
        .Y(n6818) );
  MX4X1 U8604 ( .A(\registers[616][6] ), .B(\registers[617][6] ), .C(
        \registers[618][6] ), .D(\registers[619][6] ), .S0(n7583), .S1(n7815), 
        .Y(n6823) );
  MX4X1 U8605 ( .A(\registers[520][6] ), .B(\registers[521][6] ), .C(
        \registers[522][6] ), .D(\registers[523][6] ), .S0(n7585), .S1(n7817), 
        .Y(n6854) );
  MX4X1 U8606 ( .A(\registers[568][6] ), .B(\registers[569][6] ), .C(
        \registers[570][6] ), .D(\registers[571][6] ), .S0(n7584), .S1(n7816), 
        .Y(n6839) );
  MX4X1 U8607 ( .A(\registers[552][6] ), .B(\registers[553][6] ), .C(
        \registers[554][6] ), .D(\registers[555][6] ), .S0(n7585), .S1(n7816), 
        .Y(n6844) );
  MX4X1 U8608 ( .A(\registers[712][6] ), .B(\registers[713][6] ), .C(
        \registers[714][6] ), .D(\registers[715][6] ), .S0(n7581), .S1(n7813), 
        .Y(n6791) );
  MX4X1 U8609 ( .A(\registers[760][6] ), .B(\registers[761][6] ), .C(
        \registers[762][6] ), .D(\registers[763][6] ), .S0(n7580), .S1(n7812), 
        .Y(n6776) );
  MX4X1 U8610 ( .A(\registers[744][6] ), .B(\registers[745][6] ), .C(
        \registers[746][6] ), .D(\registers[747][6] ), .S0(n7581), .S1(n7812), 
        .Y(n6781) );
  MX4X1 U8611 ( .A(\registers[648][6] ), .B(\registers[649][6] ), .C(
        \registers[650][6] ), .D(\registers[651][6] ), .S0(n7583), .S1(n7814), 
        .Y(n6812) );
  MX4X1 U8612 ( .A(\registers[696][6] ), .B(\registers[697][6] ), .C(
        \registers[698][6] ), .D(\registers[699][6] ), .S0(n7582), .S1(n7813), 
        .Y(n6797) );
  MX4X1 U8613 ( .A(\registers[680][6] ), .B(\registers[681][6] ), .C(
        \registers[682][6] ), .D(\registers[683][6] ), .S0(n7582), .S1(n7814), 
        .Y(n6802) );
  MX4X1 U8614 ( .A(\registers[328][7] ), .B(\registers[329][7] ), .C(
        \registers[330][7] ), .D(\registers[331][7] ), .S0(n7611), .S1(n7840), 
        .Y(n7258) );
  MX4X1 U8615 ( .A(\registers[376][7] ), .B(\registers[377][7] ), .C(
        \registers[378][7] ), .D(\registers[379][7] ), .S0(n7610), .S1(n7839), 
        .Y(n7243) );
  MX4X1 U8616 ( .A(\registers[360][7] ), .B(\registers[361][7] ), .C(
        \registers[362][7] ), .D(\registers[363][7] ), .S0(n7610), .S1(n7840), 
        .Y(n7248) );
  MX4X1 U8617 ( .A(\registers[200][7] ), .B(\registers[201][7] ), .C(
        \registers[202][7] ), .D(\registers[203][7] ), .S0(n7613), .S1(n7843), 
        .Y(n7301) );
  MX4X1 U8618 ( .A(\registers[248][7] ), .B(\registers[249][7] ), .C(
        \registers[250][7] ), .D(\registers[251][7] ), .S0(n7612), .S1(n7842), 
        .Y(n7286) );
  MX4X1 U8619 ( .A(\registers[232][7] ), .B(\registers[233][7] ), .C(
        \registers[234][7] ), .D(\registers[235][7] ), .S0(n7613), .S1(n7842), 
        .Y(n7291) );
  MX4X1 U8620 ( .A(\registers[72][7] ), .B(\registers[73][7] ), .C(
        \registers[74][7] ), .D(\registers[75][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7343) );
  MX4X1 U8621 ( .A(\registers[120][7] ), .B(\registers[121][7] ), .C(
        \registers[122][7] ), .D(\registers[123][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7328) );
  MX4X1 U8622 ( .A(\registers[104][7] ), .B(\registers[105][7] ), .C(
        \registers[106][7] ), .D(\registers[107][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7333) );
  MX4X1 U8623 ( .A(\registers[8][7] ), .B(\registers[9][7] ), .C(
        \registers[10][7] ), .D(\registers[11][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7364) );
  MX4X1 U8624 ( .A(\registers[56][7] ), .B(\registers[57][7] ), .C(
        \registers[58][7] ), .D(\registers[59][7] ), .S0(n7616), .S1(n7845), 
        .Y(n7349) );
  MX4X1 U8625 ( .A(\registers[40][7] ), .B(\registers[41][7] ), .C(
        \registers[42][7] ), .D(\registers[43][7] ), .S0(n7617), .S1(n7846), 
        .Y(n7354) );
  MX4X1 U8626 ( .A(\registers[136][7] ), .B(\registers[137][7] ), .C(
        \registers[138][7] ), .D(\registers[139][7] ), .S0(n7615), .S1(n7844), 
        .Y(n7322) );
  MX4X1 U8627 ( .A(\registers[184][7] ), .B(\registers[185][7] ), .C(
        \registers[186][7] ), .D(\registers[187][7] ), .S0(n7614), .S1(n7843), 
        .Y(n7307) );
  MX4X1 U8628 ( .A(\registers[168][7] ), .B(\registers[169][7] ), .C(
        \registers[170][7] ), .D(\registers[171][7] ), .S0(n7614), .S1(n7843), 
        .Y(n7312) );
  MX4X1 U8629 ( .A(\registers[840][7] ), .B(\registers[841][7] ), .C(
        \registers[842][7] ), .D(\registers[843][7] ), .S0(n7600), .S1(n7830), 
        .Y(n7088) );
  MX4X1 U8630 ( .A(\registers[888][7] ), .B(\registers[889][7] ), .C(
        \registers[890][7] ), .D(\registers[891][7] ), .S0(n7599), .S1(n7829), 
        .Y(n7073) );
  MX4X1 U8631 ( .A(\registers[872][7] ), .B(\registers[873][7] ), .C(
        \registers[874][7] ), .D(\registers[875][7] ), .S0(n7599), .S1(n7830), 
        .Y(n7078) );
  MX4X1 U8632 ( .A(\registers[776][7] ), .B(\registers[777][7] ), .C(
        \registers[778][7] ), .D(\registers[779][7] ), .S0(n7601), .S1(n7832), 
        .Y(n7109) );
  MX4X1 U8633 ( .A(\registers[824][7] ), .B(\registers[825][7] ), .C(
        \registers[826][7] ), .D(\registers[827][7] ), .S0(n7600), .S1(n7831), 
        .Y(n7094) );
  MX4X1 U8634 ( .A(\registers[808][7] ), .B(\registers[809][7] ), .C(
        \registers[810][7] ), .D(\registers[811][7] ), .S0(n7601), .S1(n7831), 
        .Y(n7099) );
  MX4X1 U8635 ( .A(\registers[968][7] ), .B(\registers[969][7] ), .C(
        \registers[970][7] ), .D(\registers[971][7] ), .S0(n7597), .S1(n7828), 
        .Y(n7046) );
  MX4X1 U8636 ( .A(\registers[1016][7] ), .B(\registers[1017][7] ), .C(
        \registers[1018][7] ), .D(\registers[1019][7] ), .S0(n7596), .S1(n7827), .Y(n7031) );
  MX4X1 U8637 ( .A(\registers[1000][7] ), .B(\registers[1001][7] ), .C(
        \registers[1002][7] ), .D(\registers[1003][7] ), .S0(n7597), .S1(n7827), .Y(n7036) );
  MX4X1 U8638 ( .A(\registers[904][7] ), .B(\registers[905][7] ), .C(
        \registers[906][7] ), .D(\registers[907][7] ), .S0(n7599), .S1(n7829), 
        .Y(n7067) );
  MX4X1 U8639 ( .A(\registers[952][7] ), .B(\registers[953][7] ), .C(
        \registers[954][7] ), .D(\registers[955][7] ), .S0(n7598), .S1(n7828), 
        .Y(n7052) );
  MX4X1 U8640 ( .A(\registers[936][7] ), .B(\registers[937][7] ), .C(
        \registers[938][7] ), .D(\registers[939][7] ), .S0(n7598), .S1(n7828), 
        .Y(n7057) );
  MX4X1 U8641 ( .A(\registers[584][7] ), .B(\registers[585][7] ), .C(
        \registers[586][7] ), .D(\registers[587][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7173) );
  MX4X1 U8642 ( .A(\registers[632][7] ), .B(\registers[633][7] ), .C(
        \registers[634][7] ), .D(\registers[635][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7158) );
  MX4X1 U8643 ( .A(\registers[616][7] ), .B(\registers[617][7] ), .C(
        \registers[618][7] ), .D(\registers[619][7] ), .S0(n7605), .S1(n7835), 
        .Y(n7163) );
  MX4X1 U8644 ( .A(\registers[520][7] ), .B(\registers[521][7] ), .C(
        \registers[522][7] ), .D(\registers[523][7] ), .S0(n7607), .S1(n7836), 
        .Y(n7194) );
  MX4X1 U8645 ( .A(\registers[568][7] ), .B(\registers[569][7] ), .C(
        \registers[570][7] ), .D(\registers[571][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7179) );
  MX4X1 U8646 ( .A(\registers[552][7] ), .B(\registers[553][7] ), .C(
        \registers[554][7] ), .D(\registers[555][7] ), .S0(n7606), .S1(n7836), 
        .Y(n7184) );
  MX4X1 U8647 ( .A(\registers[712][7] ), .B(\registers[713][7] ), .C(
        \registers[714][7] ), .D(\registers[715][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7131) );
  MX4X1 U8648 ( .A(\registers[760][7] ), .B(\registers[761][7] ), .C(
        \registers[762][7] ), .D(\registers[763][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7116) );
  MX4X1 U8649 ( .A(\registers[744][7] ), .B(\registers[745][7] ), .C(
        \registers[746][7] ), .D(\registers[747][7] ), .S0(n7602), .S1(n7832), 
        .Y(n7121) );
  MX4X1 U8650 ( .A(\registers[648][7] ), .B(\registers[649][7] ), .C(
        \registers[650][7] ), .D(\registers[651][7] ), .S0(n7604), .S1(n7834), 
        .Y(n7152) );
  MX4X1 U8651 ( .A(\registers[696][7] ), .B(\registers[697][7] ), .C(
        \registers[698][7] ), .D(\registers[699][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7137) );
  MX4X1 U8652 ( .A(\registers[680][7] ), .B(\registers[681][7] ), .C(
        \registers[682][7] ), .D(\registers[683][7] ), .S0(n7603), .S1(n7833), 
        .Y(n7142) );
  MX4X1 U8653 ( .A(n1444), .B(n1442), .C(n1443), .D(n1441), .S0(n4587), .S1(
        n4529), .Y(n1445) );
  MX4X1 U8654 ( .A(\registers[296][0] ), .B(\registers[297][0] ), .C(
        \registers[298][0] ), .D(\registers[299][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1442) );
  MX4X1 U8655 ( .A(\registers[300][0] ), .B(\registers[301][0] ), .C(
        \registers[302][0] ), .D(\registers[303][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1441) );
  MX4X1 U8656 ( .A(\registers[288][0] ), .B(\registers[289][0] ), .C(
        \registers[290][0] ), .D(\registers[291][0] ), .S0(n4119), .S1(n4360), 
        .Y(n1444) );
  MX4X1 U8657 ( .A(n1377), .B(n1375), .C(n1376), .D(n1374), .S0(n4588), .S1(
        n4528), .Y(n1378) );
  MX4X1 U8658 ( .A(\registers[488][0] ), .B(\registers[489][0] ), .C(
        \registers[490][0] ), .D(\registers[491][0] ), .S0(n4115), .S1(n4356), 
        .Y(n1375) );
  MX4X1 U8659 ( .A(\registers[492][0] ), .B(\registers[493][0] ), .C(
        \registers[494][0] ), .D(\registers[495][0] ), .S0(n4115), .S1(n4356), 
        .Y(n1374) );
  MX4X1 U8660 ( .A(\registers[480][0] ), .B(\registers[481][0] ), .C(
        \registers[482][0] ), .D(\registers[483][0] ), .S0(n4115), .S1(n4356), 
        .Y(n1377) );
  MX4X1 U8661 ( .A(n1398), .B(n1396), .C(n1397), .D(n1395), .S0(n4589), .S1(
        n4528), .Y(n1399) );
  MX4X1 U8662 ( .A(\registers[424][0] ), .B(\registers[425][0] ), .C(
        \registers[426][0] ), .D(\registers[427][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1396) );
  MX4X1 U8663 ( .A(\registers[428][0] ), .B(\registers[429][0] ), .C(
        \registers[430][0] ), .D(\registers[431][0] ), .S0(n4116), .S1(n4357), 
        .Y(n1395) );
  MX4X1 U8664 ( .A(\registers[416][0] ), .B(\registers[417][0] ), .C(
        \registers[418][0] ), .D(\registers[419][0] ), .S0(n4116), .S1(n4358), 
        .Y(n1398) );
  MX4X1 U8665 ( .A(n1800), .B(n1798), .C(n1799), .D(n1797), .S0(n4592), .S1(
        n4534), .Y(n1801) );
  MX4X1 U8666 ( .A(\registers[296][1] ), .B(\registers[297][1] ), .C(
        \registers[298][1] ), .D(\registers[299][1] ), .S0(n4140), .S1(n4380), 
        .Y(n1798) );
  MX4X1 U8667 ( .A(\registers[300][1] ), .B(\registers[301][1] ), .C(
        \registers[302][1] ), .D(\registers[303][1] ), .S0(n4140), .S1(n4380), 
        .Y(n1797) );
  MX4X1 U8668 ( .A(\registers[288][1] ), .B(\registers[289][1] ), .C(
        \registers[290][1] ), .D(\registers[291][1] ), .S0(n4140), .S1(n4380), 
        .Y(n1800) );
  MX4X1 U8669 ( .A(n1735), .B(n1733), .C(n1734), .D(n1732), .S0(n4591), .S1(
        n4533), .Y(n1736) );
  MX4X1 U8670 ( .A(\registers[488][1] ), .B(\registers[489][1] ), .C(
        \registers[490][1] ), .D(\registers[491][1] ), .S0(n4136), .S1(n4376), 
        .Y(n1733) );
  MX4X1 U8671 ( .A(\registers[492][1] ), .B(\registers[493][1] ), .C(
        \registers[494][1] ), .D(\registers[495][1] ), .S0(n4136), .S1(n4376), 
        .Y(n1732) );
  MX4X1 U8672 ( .A(\registers[480][1] ), .B(\registers[481][1] ), .C(
        \registers[482][1] ), .D(\registers[483][1] ), .S0(n4136), .S1(n4376), 
        .Y(n1735) );
  MX4X1 U8673 ( .A(n1757), .B(n1755), .C(n1756), .D(n1754), .S0(n4591), .S1(
        n4533), .Y(n1758) );
  MX4X1 U8674 ( .A(\registers[424][1] ), .B(\registers[425][1] ), .C(
        \registers[426][1] ), .D(\registers[427][1] ), .S0(n4138), .S1(n4377), 
        .Y(n1755) );
  MX4X1 U8675 ( .A(\registers[428][1] ), .B(\registers[429][1] ), .C(
        \registers[430][1] ), .D(\registers[431][1] ), .S0(n4138), .S1(n4377), 
        .Y(n1754) );
  MX4X1 U8676 ( .A(\registers[416][1] ), .B(\registers[417][1] ), .C(
        \registers[418][1] ), .D(\registers[419][1] ), .S0(n4138), .S1(n4377), 
        .Y(n1757) );
  MX4X1 U8677 ( .A(n2153), .B(n2151), .C(n2152), .D(n2150), .S0(n4597), .S1(
        n4538), .Y(n2154) );
  MX4X1 U8678 ( .A(\registers[296][2] ), .B(\registers[297][2] ), .C(
        \registers[298][2] ), .D(\registers[299][2] ), .S0(n4162), .S1(n4399), 
        .Y(n2151) );
  MX4X1 U8679 ( .A(\registers[300][2] ), .B(\registers[301][2] ), .C(
        \registers[302][2] ), .D(\registers[303][2] ), .S0(n4162), .S1(n4399), 
        .Y(n2150) );
  MX4X1 U8680 ( .A(\registers[288][2] ), .B(\registers[289][2] ), .C(
        \registers[290][2] ), .D(\registers[291][2] ), .S0(n4162), .S1(n4399), 
        .Y(n2153) );
  MX4X1 U8681 ( .A(n2087), .B(n2085), .C(n2086), .D(n2084), .S0(n4596), .S1(
        n4538), .Y(n2088) );
  MX4X1 U8682 ( .A(\registers[488][2] ), .B(\registers[489][2] ), .C(
        \registers[490][2] ), .D(\registers[491][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2085) );
  MX4X1 U8683 ( .A(\registers[492][2] ), .B(\registers[493][2] ), .C(
        \registers[494][2] ), .D(\registers[495][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2084) );
  MX4X1 U8684 ( .A(\registers[480][2] ), .B(\registers[481][2] ), .C(
        \registers[482][2] ), .D(\registers[483][2] ), .S0(n4158), .S1(n4396), 
        .Y(n2087) );
  MX4X1 U8685 ( .A(n2109), .B(n2107), .C(n2108), .D(n2106), .S0(n4597), .S1(
        n4538), .Y(n2110) );
  MX4X1 U8686 ( .A(\registers[424][2] ), .B(\registers[425][2] ), .C(
        \registers[426][2] ), .D(\registers[427][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2107) );
  MX4X1 U8687 ( .A(\registers[428][2] ), .B(\registers[429][2] ), .C(
        \registers[430][2] ), .D(\registers[431][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2106) );
  MX4X1 U8688 ( .A(\registers[416][2] ), .B(\registers[417][2] ), .C(
        \registers[418][2] ), .D(\registers[419][2] ), .S0(n4159), .S1(n4397), 
        .Y(n2109) );
  MX4X1 U8689 ( .A(n2566), .B(n2564), .C(n2565), .D(n2563), .S0(n4603), .S1(
        n4543), .Y(n2567) );
  MX4X1 U8690 ( .A(\registers[296][3] ), .B(\registers[297][3] ), .C(
        \registers[298][3] ), .D(\registers[299][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2564) );
  MX4X1 U8691 ( .A(\registers[300][3] ), .B(\registers[301][3] ), .C(
        \registers[302][3] ), .D(\registers[303][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2563) );
  MX4X1 U8692 ( .A(\registers[288][3] ), .B(\registers[289][3] ), .C(
        \registers[290][3] ), .D(\registers[291][3] ), .S0(n4183), .S1(n4419), 
        .Y(n2566) );
  MX4X1 U8693 ( .A(n2503), .B(n2501), .C(n2502), .D(n2500), .S0(n4602), .S1(
        n4542), .Y(n2504) );
  MX4X1 U8694 ( .A(\registers[488][3] ), .B(\registers[489][3] ), .C(
        \registers[490][3] ), .D(\registers[491][3] ), .S0(n4179), .S1(n4415), 
        .Y(n2501) );
  MX4X1 U8695 ( .A(\registers[492][3] ), .B(\registers[493][3] ), .C(
        \registers[494][3] ), .D(\registers[495][3] ), .S0(n4179), .S1(n4415), 
        .Y(n2500) );
  MX4X1 U8696 ( .A(\registers[480][3] ), .B(\registers[481][3] ), .C(
        \registers[482][3] ), .D(\registers[483][3] ), .S0(n4179), .S1(n4415), 
        .Y(n2503) );
  MX4X1 U8697 ( .A(n2524), .B(n2522), .C(n2523), .D(n2521), .S0(n4602), .S1(
        n4543), .Y(n2525) );
  MX4X1 U8698 ( .A(\registers[424][3] ), .B(\registers[425][3] ), .C(
        \registers[426][3] ), .D(\registers[427][3] ), .S0(n4180), .S1(n4417), 
        .Y(n2522) );
  MX4X1 U8699 ( .A(\registers[428][3] ), .B(\registers[429][3] ), .C(
        \registers[430][3] ), .D(\registers[431][3] ), .S0(n4180), .S1(n4416), 
        .Y(n2521) );
  MX4X1 U8700 ( .A(\registers[416][3] ), .B(\registers[417][3] ), .C(
        \registers[418][3] ), .D(\registers[419][3] ), .S0(n4180), .S1(n4417), 
        .Y(n2524) );
  MX4X1 U8701 ( .A(n2906), .B(n2904), .C(n2905), .D(n2903), .S0(n4608), .S1(
        n4547), .Y(n2907) );
  MX4X1 U8702 ( .A(\registers[296][4] ), .B(\registers[297][4] ), .C(
        \registers[298][4] ), .D(\registers[299][4] ), .S0(n4204), .S1(n4439), 
        .Y(n2904) );
  MX4X1 U8703 ( .A(\registers[300][4] ), .B(\registers[301][4] ), .C(
        \registers[302][4] ), .D(\registers[303][4] ), .S0(n4204), .S1(n4439), 
        .Y(n2903) );
  MX4X1 U8704 ( .A(\registers[288][4] ), .B(\registers[289][4] ), .C(
        \registers[290][4] ), .D(\registers[291][4] ), .S0(n4204), .S1(n4439), 
        .Y(n2906) );
  MX4X1 U8705 ( .A(n2843), .B(n2841), .C(n2842), .D(n2840), .S0(n4607), .S1(
        n4546), .Y(n2844) );
  MX4X1 U8706 ( .A(\registers[488][4] ), .B(\registers[489][4] ), .C(
        \registers[490][4] ), .D(\registers[491][4] ), .S0(n4200), .S1(n4435), 
        .Y(n2841) );
  MX4X1 U8707 ( .A(\registers[492][4] ), .B(\registers[493][4] ), .C(
        \registers[494][4] ), .D(\registers[495][4] ), .S0(n4200), .S1(n4435), 
        .Y(n2840) );
  MX4X1 U8708 ( .A(\registers[480][4] ), .B(\registers[481][4] ), .C(
        \registers[482][4] ), .D(\registers[483][4] ), .S0(n4200), .S1(n4435), 
        .Y(n2843) );
  MX4X1 U8709 ( .A(n2864), .B(n2862), .C(n2863), .D(n2861), .S0(n4607), .S1(
        n4547), .Y(n2865) );
  MX4X1 U8710 ( .A(\registers[424][4] ), .B(\registers[425][4] ), .C(
        \registers[426][4] ), .D(\registers[427][4] ), .S0(n4202), .S1(n4436), 
        .Y(n2862) );
  MX4X1 U8711 ( .A(\registers[428][4] ), .B(\registers[429][4] ), .C(
        \registers[430][4] ), .D(\registers[431][4] ), .S0(n4202), .S1(n4436), 
        .Y(n2861) );
  MX4X1 U8712 ( .A(\registers[416][4] ), .B(\registers[417][4] ), .C(
        \registers[418][4] ), .D(\registers[419][4] ), .S0(n4202), .S1(n4436), 
        .Y(n2864) );
  MX4X1 U8713 ( .A(n3246), .B(n3244), .C(n3245), .D(n3243), .S0(n4613), .S1(
        n4552), .Y(n3247) );
  MX4X1 U8714 ( .A(\registers[296][5] ), .B(\registers[297][5] ), .C(
        \registers[298][5] ), .D(\registers[299][5] ), .S0(n4226), .S1(n4458), 
        .Y(n3244) );
  MX4X1 U8715 ( .A(\registers[300][5] ), .B(\registers[301][5] ), .C(
        \registers[302][5] ), .D(\registers[303][5] ), .S0(n4226), .S1(n4458), 
        .Y(n3243) );
  MX4X1 U8716 ( .A(\registers[288][5] ), .B(\registers[289][5] ), .C(
        \registers[290][5] ), .D(\registers[291][5] ), .S0(n4226), .S1(n4459), 
        .Y(n3246) );
  MX4X1 U8717 ( .A(n3183), .B(n3181), .C(n3182), .D(n3180), .S0(n4612), .S1(
        n4551), .Y(n3184) );
  MX4X1 U8718 ( .A(\registers[488][5] ), .B(\registers[489][5] ), .C(
        \registers[490][5] ), .D(\registers[491][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3181) );
  MX4X1 U8719 ( .A(\registers[492][5] ), .B(\registers[493][5] ), .C(
        \registers[494][5] ), .D(\registers[495][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3180) );
  MX4X1 U8720 ( .A(\registers[480][5] ), .B(\registers[481][5] ), .C(
        \registers[482][5] ), .D(\registers[483][5] ), .S0(n4222), .S1(n4455), 
        .Y(n3183) );
  MX4X1 U8721 ( .A(n3204), .B(n3202), .C(n3203), .D(n3201), .S0(n4613), .S1(
        n4552), .Y(n3205) );
  MX4X1 U8722 ( .A(\registers[424][5] ), .B(\registers[425][5] ), .C(
        \registers[426][5] ), .D(\registers[427][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3202) );
  MX4X1 U8723 ( .A(\registers[428][5] ), .B(\registers[429][5] ), .C(
        \registers[430][5] ), .D(\registers[431][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3201) );
  MX4X1 U8724 ( .A(\registers[416][5] ), .B(\registers[417][5] ), .C(
        \registers[418][5] ), .D(\registers[419][5] ), .S0(n4223), .S1(n4456), 
        .Y(n3204) );
  MX4X1 U8725 ( .A(n3586), .B(n3584), .C(n3585), .D(n3583), .S0(n4619), .S1(
        n4557), .Y(n3587) );
  MX4X1 U8726 ( .A(\registers[296][6] ), .B(\registers[297][6] ), .C(
        \registers[298][6] ), .D(\registers[299][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3584) );
  MX4X1 U8727 ( .A(\registers[300][6] ), .B(\registers[301][6] ), .C(
        \registers[302][6] ), .D(\registers[303][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3583) );
  MX4X1 U8728 ( .A(\registers[288][6] ), .B(\registers[289][6] ), .C(
        \registers[290][6] ), .D(\registers[291][6] ), .S0(n4247), .S1(n4478), 
        .Y(n3586) );
  MX4X1 U8729 ( .A(n3523), .B(n3521), .C(n3522), .D(n3520), .S0(n4618), .S1(
        n4556), .Y(n3524) );
  MX4X1 U8730 ( .A(\registers[488][6] ), .B(\registers[489][6] ), .C(
        \registers[490][6] ), .D(\registers[491][6] ), .S0(n4243), .S1(n4474), 
        .Y(n3521) );
  MX4X1 U8731 ( .A(\registers[492][6] ), .B(\registers[493][6] ), .C(
        \registers[494][6] ), .D(\registers[495][6] ), .S0(n4243), .S1(n4474), 
        .Y(n3520) );
  MX4X1 U8732 ( .A(\registers[480][6] ), .B(\registers[481][6] ), .C(
        \registers[482][6] ), .D(\registers[483][6] ), .S0(n4243), .S1(n4475), 
        .Y(n3523) );
  MX4X1 U8733 ( .A(n3544), .B(n3542), .C(n3543), .D(n3541), .S0(n4618), .S1(
        n4557), .Y(n3545) );
  MX4X1 U8734 ( .A(\registers[424][6] ), .B(\registers[425][6] ), .C(
        \registers[426][6] ), .D(\registers[427][6] ), .S0(n4244), .S1(n4476), 
        .Y(n3542) );
  MX4X1 U8735 ( .A(\registers[428][6] ), .B(\registers[429][6] ), .C(
        \registers[430][6] ), .D(\registers[431][6] ), .S0(n4244), .S1(n4476), 
        .Y(n3541) );
  MX4X1 U8736 ( .A(\registers[416][6] ), .B(\registers[417][6] ), .C(
        \registers[418][6] ), .D(\registers[419][6] ), .S0(n4244), .S1(n4476), 
        .Y(n3544) );
  MX4X1 U8737 ( .A(n3926), .B(n3924), .C(n3925), .D(n3923), .S0(n4624), .S1(
        n4558), .Y(n3927) );
  MX4X1 U8738 ( .A(\registers[296][7] ), .B(\registers[297][7] ), .C(
        \registers[298][7] ), .D(\registers[299][7] ), .S0(n4268), .S1(n4497), 
        .Y(n3924) );
  MX4X1 U8739 ( .A(\registers[300][7] ), .B(\registers[301][7] ), .C(
        \registers[302][7] ), .D(\registers[303][7] ), .S0(n4268), .S1(n4497), 
        .Y(n3923) );
  MX4X1 U8740 ( .A(\registers[288][7] ), .B(\registers[289][7] ), .C(
        \registers[290][7] ), .D(\registers[291][7] ), .S0(n4268), .S1(n4497), 
        .Y(n3926) );
  MX4X1 U8741 ( .A(n3863), .B(n3861), .C(n3862), .D(n3860), .S0(n4623), .S1(
        N70), .Y(n3864) );
  MX4X1 U8742 ( .A(\registers[488][7] ), .B(\registers[489][7] ), .C(
        \registers[490][7] ), .D(\registers[491][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3861) );
  MX4X1 U8743 ( .A(\registers[492][7] ), .B(\registers[493][7] ), .C(
        \registers[494][7] ), .D(\registers[495][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3860) );
  MX4X1 U8744 ( .A(\registers[480][7] ), .B(\registers[481][7] ), .C(
        \registers[482][7] ), .D(\registers[483][7] ), .S0(n4264), .S1(n4494), 
        .Y(n3863) );
  MX4X1 U8745 ( .A(n3884), .B(n3882), .C(n3883), .D(n3881), .S0(n4623), .S1(
        n4540), .Y(n3885) );
  MX4X1 U8746 ( .A(\registers[424][7] ), .B(\registers[425][7] ), .C(
        \registers[426][7] ), .D(\registers[427][7] ), .S0(n4266), .S1(n4495), 
        .Y(n3882) );
  MX4X1 U8747 ( .A(\registers[428][7] ), .B(\registers[429][7] ), .C(
        \registers[430][7] ), .D(\registers[431][7] ), .S0(n4266), .S1(n4495), 
        .Y(n3881) );
  MX4X1 U8748 ( .A(\registers[416][7] ), .B(\registers[417][7] ), .C(
        \registers[418][7] ), .D(\registers[419][7] ), .S0(n4266), .S1(n4495), 
        .Y(n3884) );
  MX4X1 U8749 ( .A(n4891), .B(n4889), .C(n4890), .D(n4888), .S0(n7930), .S1(
        n7870), .Y(n4892) );
  MX4X1 U8750 ( .A(\registers[296][0] ), .B(\registers[297][0] ), .C(
        \registers[298][0] ), .D(\registers[299][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4889) );
  MX4X1 U8751 ( .A(\registers[300][0] ), .B(\registers[301][0] ), .C(
        \registers[302][0] ), .D(\registers[303][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4888) );
  MX4X1 U8752 ( .A(\registers[288][0] ), .B(\registers[289][0] ), .C(
        \registers[290][0] ), .D(\registers[291][0] ), .S0(n7462), .S1(n7704), 
        .Y(n4891) );
  MX4X1 U8753 ( .A(n4828), .B(n4826), .C(n4827), .D(n4825), .S0(n7931), .S1(
        n7869), .Y(n4829) );
  MX4X1 U8754 ( .A(\registers[488][0] ), .B(\registers[489][0] ), .C(
        \registers[490][0] ), .D(\registers[491][0] ), .S0(n7458), .S1(n7700), 
        .Y(n4826) );
  MX4X1 U8755 ( .A(\registers[492][0] ), .B(\registers[493][0] ), .C(
        \registers[494][0] ), .D(\registers[495][0] ), .S0(n7458), .S1(n7700), 
        .Y(n4825) );
  MX4X1 U8756 ( .A(\registers[480][0] ), .B(\registers[481][0] ), .C(
        \registers[482][0] ), .D(\registers[483][0] ), .S0(n7458), .S1(n7700), 
        .Y(n4828) );
  MX4X1 U8757 ( .A(n4849), .B(n4847), .C(n4848), .D(n4846), .S0(n7932), .S1(
        n7869), .Y(n4850) );
  MX4X1 U8758 ( .A(\registers[424][0] ), .B(\registers[425][0] ), .C(
        \registers[426][0] ), .D(\registers[427][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4847) );
  MX4X1 U8759 ( .A(\registers[428][0] ), .B(\registers[429][0] ), .C(
        \registers[430][0] ), .D(\registers[431][0] ), .S0(n7459), .S1(n7701), 
        .Y(n4846) );
  MX4X1 U8760 ( .A(\registers[416][0] ), .B(\registers[417][0] ), .C(
        \registers[418][0] ), .D(\registers[419][0] ), .S0(n7459), .S1(n7702), 
        .Y(n4849) );
  MX4X1 U8761 ( .A(n5231), .B(n5229), .C(n5230), .D(n5228), .S0(n7935), .S1(
        n7875), .Y(n5232) );
  MX4X1 U8762 ( .A(\registers[296][1] ), .B(\registers[297][1] ), .C(
        \registers[298][1] ), .D(\registers[299][1] ), .S0(n7483), .S1(n7724), 
        .Y(n5229) );
  MX4X1 U8763 ( .A(\registers[300][1] ), .B(\registers[301][1] ), .C(
        \registers[302][1] ), .D(\registers[303][1] ), .S0(n7483), .S1(n7724), 
        .Y(n5228) );
  MX4X1 U8764 ( .A(\registers[288][1] ), .B(\registers[289][1] ), .C(
        \registers[290][1] ), .D(\registers[291][1] ), .S0(n7483), .S1(n7724), 
        .Y(n5231) );
  MX4X1 U8765 ( .A(n5168), .B(n5166), .C(n5167), .D(n5165), .S0(n7934), .S1(
        n7874), .Y(n5169) );
  MX4X1 U8766 ( .A(\registers[488][1] ), .B(\registers[489][1] ), .C(
        \registers[490][1] ), .D(\registers[491][1] ), .S0(n7479), .S1(n7720), 
        .Y(n5166) );
  MX4X1 U8767 ( .A(\registers[492][1] ), .B(\registers[493][1] ), .C(
        \registers[494][1] ), .D(\registers[495][1] ), .S0(n7479), .S1(n7720), 
        .Y(n5165) );
  MX4X1 U8768 ( .A(\registers[480][1] ), .B(\registers[481][1] ), .C(
        \registers[482][1] ), .D(\registers[483][1] ), .S0(n7479), .S1(n7720), 
        .Y(n5168) );
  MX4X1 U8769 ( .A(n5189), .B(n5187), .C(n5188), .D(n5186), .S0(n7934), .S1(
        n7874), .Y(n5190) );
  MX4X1 U8770 ( .A(\registers[424][1] ), .B(\registers[425][1] ), .C(
        \registers[426][1] ), .D(\registers[427][1] ), .S0(n7481), .S1(n7721), 
        .Y(n5187) );
  MX4X1 U8771 ( .A(\registers[428][1] ), .B(\registers[429][1] ), .C(
        \registers[430][1] ), .D(\registers[431][1] ), .S0(n7481), .S1(n7721), 
        .Y(n5186) );
  MX4X1 U8772 ( .A(\registers[416][1] ), .B(\registers[417][1] ), .C(
        \registers[418][1] ), .D(\registers[419][1] ), .S0(n7481), .S1(n7721), 
        .Y(n5189) );
  MX4X1 U8773 ( .A(n5571), .B(n5569), .C(n5570), .D(n5568), .S0(n7940), .S1(
        n7879), .Y(n5572) );
  MX4X1 U8774 ( .A(\registers[296][2] ), .B(\registers[297][2] ), .C(
        \registers[298][2] ), .D(\registers[299][2] ), .S0(n7505), .S1(n7743), 
        .Y(n5569) );
  MX4X1 U8775 ( .A(\registers[300][2] ), .B(\registers[301][2] ), .C(
        \registers[302][2] ), .D(\registers[303][2] ), .S0(n7505), .S1(n7743), 
        .Y(n5568) );
  MX4X1 U8776 ( .A(\registers[288][2] ), .B(\registers[289][2] ), .C(
        \registers[290][2] ), .D(\registers[291][2] ), .S0(n7505), .S1(n7743), 
        .Y(n5571) );
  MX4X1 U8777 ( .A(n5508), .B(n5506), .C(n5507), .D(n5505), .S0(n7939), .S1(
        n7879), .Y(n5509) );
  MX4X1 U8778 ( .A(\registers[488][2] ), .B(\registers[489][2] ), .C(
        \registers[490][2] ), .D(\registers[491][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5506) );
  MX4X1 U8779 ( .A(\registers[492][2] ), .B(\registers[493][2] ), .C(
        \registers[494][2] ), .D(\registers[495][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5505) );
  MX4X1 U8780 ( .A(\registers[480][2] ), .B(\registers[481][2] ), .C(
        \registers[482][2] ), .D(\registers[483][2] ), .S0(n7501), .S1(n7740), 
        .Y(n5508) );
  MX4X1 U8781 ( .A(n5529), .B(n5527), .C(n5528), .D(n5526), .S0(n7940), .S1(
        n7879), .Y(n5530) );
  MX4X1 U8782 ( .A(\registers[424][2] ), .B(\registers[425][2] ), .C(
        \registers[426][2] ), .D(\registers[427][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5527) );
  MX4X1 U8783 ( .A(\registers[428][2] ), .B(\registers[429][2] ), .C(
        \registers[430][2] ), .D(\registers[431][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5526) );
  MX4X1 U8784 ( .A(\registers[416][2] ), .B(\registers[417][2] ), .C(
        \registers[418][2] ), .D(\registers[419][2] ), .S0(n7502), .S1(n7741), 
        .Y(n5529) );
  MX4X1 U8785 ( .A(n5911), .B(n5909), .C(n5910), .D(n5908), .S0(n7946), .S1(
        n7884), .Y(n5912) );
  MX4X1 U8786 ( .A(\registers[296][3] ), .B(\registers[297][3] ), .C(
        \registers[298][3] ), .D(\registers[299][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5909) );
  MX4X1 U8787 ( .A(\registers[300][3] ), .B(\registers[301][3] ), .C(
        \registers[302][3] ), .D(\registers[303][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5908) );
  MX4X1 U8788 ( .A(\registers[288][3] ), .B(\registers[289][3] ), .C(
        \registers[290][3] ), .D(\registers[291][3] ), .S0(n7526), .S1(n7763), 
        .Y(n5911) );
  MX4X1 U8789 ( .A(n5848), .B(n5846), .C(n5847), .D(n5845), .S0(n7945), .S1(
        n7883), .Y(n5849) );
  MX4X1 U8790 ( .A(\registers[488][3] ), .B(\registers[489][3] ), .C(
        \registers[490][3] ), .D(\registers[491][3] ), .S0(n7522), .S1(n7759), 
        .Y(n5846) );
  MX4X1 U8791 ( .A(\registers[492][3] ), .B(\registers[493][3] ), .C(
        \registers[494][3] ), .D(\registers[495][3] ), .S0(n7522), .S1(n7759), 
        .Y(n5845) );
  MX4X1 U8792 ( .A(\registers[480][3] ), .B(\registers[481][3] ), .C(
        \registers[482][3] ), .D(\registers[483][3] ), .S0(n7522), .S1(n7759), 
        .Y(n5848) );
  MX4X1 U8793 ( .A(n5869), .B(n5867), .C(n5868), .D(n5866), .S0(n7945), .S1(
        n7884), .Y(n5870) );
  MX4X1 U8794 ( .A(\registers[424][3] ), .B(\registers[425][3] ), .C(
        \registers[426][3] ), .D(\registers[427][3] ), .S0(n7523), .S1(n7761), 
        .Y(n5867) );
  MX4X1 U8795 ( .A(\registers[428][3] ), .B(\registers[429][3] ), .C(
        \registers[430][3] ), .D(\registers[431][3] ), .S0(n7523), .S1(n7760), 
        .Y(n5866) );
  MX4X1 U8796 ( .A(\registers[416][3] ), .B(\registers[417][3] ), .C(
        \registers[418][3] ), .D(\registers[419][3] ), .S0(n7523), .S1(n7761), 
        .Y(n5869) );
  MX4X1 U8797 ( .A(n6251), .B(n6249), .C(n6250), .D(n6248), .S0(n7951), .S1(
        n7889), .Y(n6252) );
  MX4X1 U8798 ( .A(\registers[296][4] ), .B(\registers[297][4] ), .C(
        \registers[298][4] ), .D(\registers[299][4] ), .S0(n7547), .S1(n7783), 
        .Y(n6249) );
  MX4X1 U8799 ( .A(\registers[300][4] ), .B(\registers[301][4] ), .C(
        \registers[302][4] ), .D(\registers[303][4] ), .S0(n7547), .S1(n7783), 
        .Y(n6248) );
  MX4X1 U8800 ( .A(\registers[288][4] ), .B(\registers[289][4] ), .C(
        \registers[290][4] ), .D(\registers[291][4] ), .S0(n7547), .S1(n7783), 
        .Y(n6251) );
  MX4X1 U8801 ( .A(n6188), .B(n6186), .C(n6187), .D(n6185), .S0(n7950), .S1(
        n7888), .Y(n6189) );
  MX4X1 U8802 ( .A(\registers[488][4] ), .B(\registers[489][4] ), .C(
        \registers[490][4] ), .D(\registers[491][4] ), .S0(n7543), .S1(n7779), 
        .Y(n6186) );
  MX4X1 U8803 ( .A(\registers[492][4] ), .B(\registers[493][4] ), .C(
        \registers[494][4] ), .D(\registers[495][4] ), .S0(n7543), .S1(n7779), 
        .Y(n6185) );
  MX4X1 U8804 ( .A(\registers[480][4] ), .B(\registers[481][4] ), .C(
        \registers[482][4] ), .D(\registers[483][4] ), .S0(n7543), .S1(n7779), 
        .Y(n6188) );
  MX4X1 U8805 ( .A(n6209), .B(n6207), .C(n6208), .D(n6206), .S0(n7950), .S1(
        n7889), .Y(n6210) );
  MX4X1 U8806 ( .A(\registers[424][4] ), .B(\registers[425][4] ), .C(
        \registers[426][4] ), .D(\registers[427][4] ), .S0(n7545), .S1(n7780), 
        .Y(n6207) );
  MX4X1 U8807 ( .A(\registers[428][4] ), .B(\registers[429][4] ), .C(
        \registers[430][4] ), .D(\registers[431][4] ), .S0(n7545), .S1(n7780), 
        .Y(n6206) );
  MX4X1 U8808 ( .A(\registers[416][4] ), .B(\registers[417][4] ), .C(
        \registers[418][4] ), .D(\registers[419][4] ), .S0(n7545), .S1(n7780), 
        .Y(n6209) );
  MX4X1 U8809 ( .A(n6591), .B(n6589), .C(n6590), .D(n6588), .S0(n7956), .S1(
        n7894), .Y(n6592) );
  MX4X1 U8810 ( .A(\registers[296][5] ), .B(\registers[297][5] ), .C(
        \registers[298][5] ), .D(\registers[299][5] ), .S0(n7569), .S1(n7802), 
        .Y(n6589) );
  MX4X1 U8811 ( .A(\registers[300][5] ), .B(\registers[301][5] ), .C(
        \registers[302][5] ), .D(\registers[303][5] ), .S0(n7569), .S1(n7802), 
        .Y(n6588) );
  MX4X1 U8812 ( .A(\registers[288][5] ), .B(\registers[289][5] ), .C(
        \registers[290][5] ), .D(\registers[291][5] ), .S0(n7569), .S1(n7803), 
        .Y(n6591) );
  MX4X1 U8813 ( .A(n6528), .B(n6526), .C(n6527), .D(n6525), .S0(n7955), .S1(
        n7893), .Y(n6529) );
  MX4X1 U8814 ( .A(\registers[488][5] ), .B(\registers[489][5] ), .C(
        \registers[490][5] ), .D(\registers[491][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6526) );
  MX4X1 U8815 ( .A(\registers[492][5] ), .B(\registers[493][5] ), .C(
        \registers[494][5] ), .D(\registers[495][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6525) );
  MX4X1 U8816 ( .A(\registers[480][5] ), .B(\registers[481][5] ), .C(
        \registers[482][5] ), .D(\registers[483][5] ), .S0(n7565), .S1(n7799), 
        .Y(n6528) );
  MX4X1 U8817 ( .A(n6549), .B(n6547), .C(n6548), .D(n6546), .S0(n7956), .S1(
        n7894), .Y(n6550) );
  MX4X1 U8818 ( .A(\registers[424][5] ), .B(\registers[425][5] ), .C(
        \registers[426][5] ), .D(\registers[427][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6547) );
  MX4X1 U8819 ( .A(\registers[428][5] ), .B(\registers[429][5] ), .C(
        \registers[430][5] ), .D(\registers[431][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6546) );
  MX4X1 U8820 ( .A(\registers[416][5] ), .B(\registers[417][5] ), .C(
        \registers[418][5] ), .D(\registers[419][5] ), .S0(n7566), .S1(n7800), 
        .Y(n6549) );
  MX4X1 U8821 ( .A(n6931), .B(n6929), .C(n6930), .D(n6928), .S0(n7962), .S1(
        n7897), .Y(n6932) );
  MX4X1 U8822 ( .A(\registers[296][6] ), .B(\registers[297][6] ), .C(
        \registers[298][6] ), .D(\registers[299][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6929) );
  MX4X1 U8823 ( .A(\registers[300][6] ), .B(\registers[301][6] ), .C(
        \registers[302][6] ), .D(\registers[303][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6928) );
  MX4X1 U8824 ( .A(\registers[288][6] ), .B(\registers[289][6] ), .C(
        \registers[290][6] ), .D(\registers[291][6] ), .S0(n7590), .S1(n7821), 
        .Y(n6931) );
  MX4X1 U8825 ( .A(n6868), .B(n6866), .C(n6867), .D(n6865), .S0(n7961), .S1(
        n7892), .Y(n6869) );
  MX4X1 U8826 ( .A(\registers[488][6] ), .B(\registers[489][6] ), .C(
        \registers[490][6] ), .D(\registers[491][6] ), .S0(n7586), .S1(n7817), 
        .Y(n6866) );
  MX4X1 U8827 ( .A(\registers[492][6] ), .B(\registers[493][6] ), .C(
        \registers[494][6] ), .D(\registers[495][6] ), .S0(n7586), .S1(n7817), 
        .Y(n6865) );
  MX4X1 U8828 ( .A(\registers[480][6] ), .B(\registers[481][6] ), .C(
        \registers[482][6] ), .D(\registers[483][6] ), .S0(n7586), .S1(n7818), 
        .Y(n6868) );
  MX4X1 U8829 ( .A(n6889), .B(n6887), .C(n6888), .D(n6886), .S0(n7961), .S1(
        n7897), .Y(n6890) );
  MX4X1 U8830 ( .A(\registers[424][6] ), .B(\registers[425][6] ), .C(
        \registers[426][6] ), .D(\registers[427][6] ), .S0(n7587), .S1(n7819), 
        .Y(n6887) );
  MX4X1 U8831 ( .A(\registers[428][6] ), .B(\registers[429][6] ), .C(
        \registers[430][6] ), .D(\registers[431][6] ), .S0(n7587), .S1(n7819), 
        .Y(n6886) );
  MX4X1 U8832 ( .A(\registers[416][6] ), .B(\registers[417][6] ), .C(
        \registers[418][6] ), .D(\registers[419][6] ), .S0(n7587), .S1(n7819), 
        .Y(n6889) );
  MX4X1 U8833 ( .A(n7208), .B(n7206), .C(n7207), .D(n7205), .S0(n7966), .S1(
        n7901), .Y(n7209) );
  MX4X1 U8834 ( .A(\registers[488][7] ), .B(\registers[489][7] ), .C(
        \registers[490][7] ), .D(\registers[491][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7206) );
  MX4X1 U8835 ( .A(\registers[492][7] ), .B(\registers[493][7] ), .C(
        \registers[494][7] ), .D(\registers[495][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7205) );
  MX4X1 U8836 ( .A(\registers[480][7] ), .B(\registers[481][7] ), .C(
        \registers[482][7] ), .D(\registers[483][7] ), .S0(n7607), .S1(n7837), 
        .Y(n7208) );
  MX4X1 U8837 ( .A(n7229), .B(n7227), .C(n7228), .D(n7226), .S0(n7966), .S1(
        n7901), .Y(n7230) );
  MX4X1 U8838 ( .A(\registers[424][7] ), .B(\registers[425][7] ), .C(
        \registers[426][7] ), .D(\registers[427][7] ), .S0(n7609), .S1(n7838), 
        .Y(n7227) );
  MX4X1 U8839 ( .A(\registers[428][7] ), .B(\registers[429][7] ), .C(
        \registers[430][7] ), .D(\registers[431][7] ), .S0(n7609), .S1(n7838), 
        .Y(n7226) );
  MX4X1 U8840 ( .A(\registers[416][7] ), .B(\registers[417][7] ), .C(
        \registers[418][7] ), .D(\registers[419][7] ), .S0(n7609), .S1(n7838), 
        .Y(n7229) );
  MX4X1 U8841 ( .A(n7271), .B(n7269), .C(n7270), .D(n7268), .S0(n7967), .S1(
        n7889), .Y(n7272) );
  MX4X1 U8842 ( .A(\registers[296][7] ), .B(\registers[297][7] ), .C(
        \registers[298][7] ), .D(\registers[299][7] ), .S0(n7611), .S1(n7841), 
        .Y(n7269) );
  MX4X1 U8843 ( .A(\registers[300][7] ), .B(\registers[301][7] ), .C(
        \registers[302][7] ), .D(\registers[303][7] ), .S0(n7611), .S1(n7841), 
        .Y(n7268) );
  MX4X1 U8844 ( .A(\registers[288][7] ), .B(\registers[289][7] ), .C(
        \registers[290][7] ), .D(\registers[291][7] ), .S0(n7611), .S1(n7841), 
        .Y(n7271) );
  INVX1 U8845 ( .A(pixel_i[10]), .Y(n8918) );
  INVX1 U8846 ( .A(pixel_i[11]), .Y(n8919) );
  INVX1 U8847 ( .A(pixel_i[1]), .Y(N1198) );
  INVX1 U8848 ( .A(pixel_i[12]), .Y(n8920) );
  OAI2BB2X1 U8849 ( .B0(n1265), .B1(n8681), .A0N(\registers[0][0] ), .A1N(
        n1266), .Y(n2429) );
  OAI2BB2X1 U8850 ( .B0(n1265), .B1(n8711), .A0N(\registers[0][1] ), .A1N(
        n1266), .Y(n2430) );
  OAI2BB2X1 U8851 ( .B0(n1265), .B1(n8739), .A0N(\registers[0][2] ), .A1N(
        n1266), .Y(n2431) );
  OAI2BB2X1 U8852 ( .B0(n1265), .B1(n8764), .A0N(\registers[0][3] ), .A1N(
        n1266), .Y(n2432) );
  OAI2BB2X1 U8853 ( .B0(n1265), .B1(n8789), .A0N(\registers[0][4] ), .A1N(
        n1266), .Y(n2433) );
  OAI2BB2X1 U8854 ( .B0(n1265), .B1(n8818), .A0N(\registers[0][5] ), .A1N(
        n1266), .Y(n2434) );
  OAI2BB2X1 U8855 ( .B0(n1265), .B1(n8847), .A0N(\registers[0][6] ), .A1N(
        n1266), .Y(n2435) );
  OAI2BB2X1 U8856 ( .B0(n1265), .B1(n8876), .A0N(\registers[0][7] ), .A1N(
        n1266), .Y(n2436) );
  NOR3X2 U8857 ( .A(ena_out), .B(rst), .C(n1264), .Y(n1212) );
  NAND2X1 U8858 ( .A(StartBit), .B(Block_Done), .Y(n1264) );
  NOR2X2 U8859 ( .A(state[0]), .B(state[1]), .Y(n1206) );
  NOR2BX2 U8860 ( .AN(state[0]), .B(state[1]), .Y(n1200) );
  NOR2BX1 U8861 ( .AN(n1194), .B(param_i[1]), .Y(n1189) );
  OAI22X1 U8862 ( .A0(n1239), .A1(n8965), .B0(param_i[1]), .B1(n1238), .Y(
        n2427) );
  AND3X2 U8863 ( .A(param_i[0]), .B(n8966), .C(n1189), .Y(n1044) );
  AND3X2 U8864 ( .A(param_i[1]), .B(n8966), .C(n1194), .Y(n1192) );
  OAI2BB2X1 U8865 ( .B0(n8443), .B1(n1149), .A0N(params[0]), .A1N(n8443), .Y(
        n2424) );
  OAI2BB2X1 U8866 ( .B0(n8443), .B1(n1148), .A0N(params[1]), .A1N(n8443), .Y(
        n2423) );
  OAI2BB2X1 U8867 ( .B0(n8443), .B1(n1147), .A0N(params[2]), .A1N(n8443), .Y(
        n2422) );
  OAI2BB2X1 U8868 ( .B0(n8443), .B1(n1146), .A0N(params[3]), .A1N(n8443), .Y(
        n2421) );
  OAI2BB2X1 U8869 ( .B0(n8443), .B1(n1145), .A0N(params[4]), .A1N(n8443), .Y(
        n2420) );
  OAI2BB2X1 U8870 ( .B0(n8443), .B1(n1144), .A0N(params[5]), .A1N(n8443), .Y(
        n2419) );
  OAI2BB2X1 U8871 ( .B0(n8443), .B1(n1143), .A0N(params[6]), .A1N(n8443), .Y(
        n2418) );
  OAI2BB2X1 U8872 ( .B0(n8443), .B1(n1142), .A0N(params[7]), .A1N(n8443), .Y(
        n2417) );
  OAI2BB2X1 U8873 ( .B0(n8444), .B1(n1141), .A0N(params[13]), .A1N(n8444), .Y(
        n2416) );
  OAI2BB2X1 U8874 ( .B0(n8444), .B1(n1140), .A0N(params[14]), .A1N(n8444), .Y(
        n2415) );
  OAI2BB2X1 U8875 ( .B0(n8444), .B1(n1139), .A0N(params[15]), .A1N(n8444), .Y(
        n2414) );
  OAI2BB2X1 U8876 ( .B0(n8444), .B1(n1138), .A0N(params[16]), .A1N(n8444), .Y(
        n2413) );
  OAI2BB2X1 U8877 ( .B0(n8444), .B1(n1137), .A0N(params[17]), .A1N(n8444), .Y(
        n2412) );
  OAI2BB2X1 U8878 ( .B0(n8444), .B1(n1136), .A0N(params[18]), .A1N(n8444), .Y(
        n2411) );
  OAI2BB2X1 U8879 ( .B0(n8444), .B1(n1135), .A0N(params[19]), .A1N(n8444), .Y(
        n2410) );
  OAI2BB2X1 U8880 ( .B0(n8444), .B1(n1134), .A0N(params[20]), .A1N(n8444), .Y(
        n2409) );
  OAI2BB2X1 U8881 ( .B0(n8446), .B1(n1126), .A0N(params[28]), .A1N(n8446), .Y(
        n2401) );
  OAI2BB2X1 U8882 ( .B0(n8446), .B1(n1125), .A0N(params[29]), .A1N(n8446), .Y(
        n2400) );
  OAI2BB2X1 U8883 ( .B0(n8446), .B1(n1124), .A0N(params[30]), .A1N(n8446), .Y(
        n2399) );
  OAI2BB2X1 U8884 ( .B0(n8446), .B1(n1123), .A0N(params[31]), .A1N(n8446), .Y(
        n2398) );
  OAI2BB2X1 U8885 ( .B0(n8446), .B1(n1122), .A0N(params[32]), .A1N(n8446), .Y(
        n2397) );
  OAI2BB2X1 U8886 ( .B0(n8446), .B1(n1121), .A0N(params[33]), .A1N(n8446), .Y(
        n2396) );
  OAI2BB2X1 U8887 ( .B0(n8446), .B1(n1120), .A0N(params[34]), .A1N(n8446), .Y(
        n2395) );
  OAI2BB2X1 U8888 ( .B0(n8445), .B1(n1133), .A0N(params[21]), .A1N(n8445), .Y(
        n2408) );
  OAI2BB2X1 U8889 ( .B0(n8445), .B1(n1132), .A0N(params[22]), .A1N(n8445), .Y(
        n2407) );
  OAI2BB2X1 U8890 ( .B0(n8445), .B1(n1131), .A0N(params[23]), .A1N(n8445), .Y(
        n2406) );
  OAI2BB2X1 U8891 ( .B0(n8445), .B1(n1130), .A0N(params[24]), .A1N(n8445), .Y(
        n2405) );
  OAI2BB2X1 U8892 ( .B0(n8445), .B1(n1129), .A0N(params[25]), .A1N(n8445), .Y(
        n2404) );
  OAI2BB2X1 U8893 ( .B0(n8445), .B1(n1128), .A0N(params[26]), .A1N(n8445), .Y(
        n2403) );
  OAI2BB2X1 U8894 ( .B0(n8445), .B1(n1127), .A0N(params[27]), .A1N(n8445), .Y(
        n2402) );
  OAI2BB2X1 U8895 ( .B0(n8447), .B1(n1119), .A0N(params[35]), .A1N(n8447), .Y(
        n2394) );
  OAI2BB2X1 U8896 ( .B0(n8447), .B1(n1118), .A0N(params[36]), .A1N(n8447), .Y(
        n2393) );
  OAI2BB2X1 U8897 ( .B0(n8447), .B1(n1117), .A0N(params[37]), .A1N(n8447), .Y(
        n2392) );
  OAI2BB2X1 U8898 ( .B0(n8447), .B1(n1116), .A0N(params[38]), .A1N(n8447), .Y(
        n2391) );
  OAI2BB2X1 U8899 ( .B0(n8447), .B1(n1115), .A0N(params[39]), .A1N(n8447), .Y(
        n2390) );
  OAI2BB2X1 U8900 ( .B0(n8447), .B1(n1114), .A0N(params[40]), .A1N(n8447), .Y(
        n2389) );
  BUFX3 U8901 ( .A(n1190), .Y(n8446) );
  NAND3X1 U8902 ( .A(param_i[2]), .B(n8964), .C(n1189), .Y(n1190) );
  BUFX3 U8903 ( .A(n1191), .Y(n8445) );
  NAND2X1 U8904 ( .A(n1192), .B(param_i[0]), .Y(n1191) );
  BUFX3 U8905 ( .A(n1188), .Y(n8447) );
  NAND3X1 U8906 ( .A(param_i[0]), .B(param_i[2]), .C(n1189), .Y(n1188) );
  OAI32X1 U8907 ( .A0(n1197), .A1(param_i[0]), .A2(n8958), .B0(n8964), .B1(
        n1240), .Y(n2428) );
  AOI21X1 U8908 ( .A0(n1186), .A1(param_i[0]), .B0(param_i[3]), .Y(n1241) );
  NAND3X1 U8909 ( .A(param_i[0]), .B(n1240), .C(n8961), .Y(n1238) );
  INVX1 U8910 ( .A(param_i[1]), .Y(n8965) );
  OAI2BB2X1 U8911 ( .B0(n8448), .B1(n1113), .A0N(params[41]), .A1N(n8448), .Y(
        n2388) );
  OAI2BB2X1 U8912 ( .B0(n8448), .B1(n1112), .A0N(params[42]), .A1N(n8448), .Y(
        n2387) );
  OAI2BB2X1 U8913 ( .B0(n8448), .B1(n1111), .A0N(params[43]), .A1N(n8448), .Y(
        n2386) );
  OAI2BB2X1 U8914 ( .B0(n8448), .B1(n1110), .A0N(params[44]), .A1N(n8448), .Y(
        n2385) );
  OAI2BB2X1 U8915 ( .B0(n8448), .B1(n1109), .A0N(params[45]), .A1N(n8448), .Y(
        n2384) );
  OAI2BB2X1 U8916 ( .B0(n8448), .B1(n1108), .A0N(params[46]), .A1N(n8448), .Y(
        n2383) );
  INVX1 U8917 ( .A(n1262), .Y(n8957) );
  AOI32X1 U8918 ( .A0(StartBit), .A1(n8973), .A2(n1263), .B0(n8962), .B1(
        \registers[0][0] ), .Y(n1262) );
  INVX1 U8919 ( .A(n1263), .Y(n8962) );
  NAND3BX1 U8920 ( .AN(ena_out), .B(n8973), .C(n1264), .Y(n1263) );
  XOR2X1 U8921 ( .A(pixel_i[9]), .B(\r402/carry[9] ), .Y(N1206) );
  AND2X1 U8922 ( .A(\r402/carry[8] ), .B(pixel_i[8]), .Y(\r402/carry[9] ) );
  XOR2X1 U8923 ( .A(pixel_i[8]), .B(\r402/carry[8] ), .Y(N1205) );
  AND2X1 U8924 ( .A(\r402/carry[7] ), .B(pixel_i[7]), .Y(\r402/carry[8] ) );
  XOR2X1 U8925 ( .A(pixel_i[7]), .B(\r402/carry[7] ), .Y(N1204) );
  AND2X1 U8926 ( .A(\r402/carry[6] ), .B(pixel_i[6]), .Y(\r402/carry[7] ) );
  XOR2X1 U8927 ( .A(pixel_i[6]), .B(\r402/carry[6] ), .Y(N1203) );
  AND2X1 U8928 ( .A(\r402/carry[5] ), .B(n9), .Y(\r402/carry[6] ) );
  XOR2X1 U8929 ( .A(n9), .B(\r402/carry[5] ), .Y(N1202) );
  AND2X1 U8930 ( .A(\r402/carry[4] ), .B(pixel_i[4]), .Y(\r402/carry[5] ) );
  XOR2X1 U8931 ( .A(pixel_i[4]), .B(\r402/carry[4] ), .Y(N1201) );
  OR2X1 U8932 ( .A(pixel_i[3]), .B(\r402/carry[3] ), .Y(\r402/carry[4] ) );
  XNOR2X1 U8933 ( .A(\r402/carry[3] ), .B(pixel_i[3]), .Y(N1200) );
  AND2X1 U8934 ( .A(pixel_i[1]), .B(pixel_i[2]), .Y(\r402/carry[3] ) );
  XOR2X1 U8935 ( .A(pixel_i[2]), .B(pixel_i[1]), .Y(N1199) );
  NOR2X1 U8936 ( .A(M2[19]), .B(M2[18]), .Y(n8887) );
  NOR4BX1 U8937 ( .AN(n8887), .B(M2[16]), .C(M2[15]), .D(M2[17]), .Y(n8914) );
  NAND2BX1 U8938 ( .AN(M2[7]), .B(pixel_i[7]), .Y(n8888) );
  OAI222XL U8939 ( .A0(n8888), .A1(n8917), .B0(M2[8]), .B1(n8888), .C0(M2[8]), 
        .C1(n8917), .Y(n8889) );
  OAI222XL U8940 ( .A0(pixel_i[9]), .A1(n8889), .B0(n8889), .B1(n6), .C0(
        pixel_i[9]), .C1(n6), .Y(n8908) );
  NAND2BX1 U8941 ( .AN(M2[4]), .B(pixel_i[4]), .Y(n8890) );
  OAI222XL U8942 ( .A0(n8), .A1(n8890), .B0(M2[5]), .B1(n8890), .C0(M2[5]), 
        .C1(n8), .Y(n8891) );
  OAI222XL U8943 ( .A0(pixel_i[6]), .A1(n8891), .B0(n7), .B1(n8891), .C0(
        pixel_i[6]), .C1(n7), .Y(n8906) );
  NOR2BX1 U8944 ( .AN(M2[4]), .B(pixel_i[4]), .Y(n8892) );
  OAI22X1 U8945 ( .A0(n8892), .A1(n8), .B0(M2[5]), .B1(n8892), .Y(n8900) );
  NAND2BX1 U8946 ( .AN(pixel_i[2]), .B(M2[2]), .Y(n8893) );
  AOI22X1 U8947 ( .A0(n8893), .A1(n5), .B0(n8893), .B1(pixel_i[3]), .Y(n8898)
         );
  AOI22X1 U8948 ( .A0(M2[1]), .A1(N1198), .B0(M2[0]), .B1(n8915), .Y(n8894) );
  AOI2BB1X1 U8949 ( .A0N(N1198), .A1N(M2[1]), .B0(n8894), .Y(n8897) );
  NOR2BX1 U8950 ( .AN(pixel_i[2]), .B(M2[2]), .Y(n8895) );
  AOI22X1 U8951 ( .A0(n8895), .A1(n5), .B0(pixel_i[3]), .B1(n8895), .Y(n8896)
         );
  OAI221XL U8952 ( .A0(M2[3]), .A1(n8916), .B0(n8898), .B1(n8897), .C0(n8896), 
        .Y(n8899) );
  OAI211X1 U8953 ( .A0(pixel_i[6]), .A1(n7), .B0(n8900), .C0(n8899), .Y(n8905)
         );
  NOR2BX1 U8954 ( .AN(M2[7]), .B(pixel_i[7]), .Y(n8901) );
  OAI22X1 U8955 ( .A0(n8901), .A1(n8917), .B0(M2[8]), .B1(n8901), .Y(n8902) );
  OAI21XL U8956 ( .A0(pixel_i[9]), .A1(n6), .B0(n8902), .Y(n8903) );
  OAI22X1 U8957 ( .A0(n8903), .A1(M2[10]), .B0(n8903), .B1(n8918), .Y(n8904)
         );
  OAI2BB1X1 U8958 ( .A0N(n8906), .A1N(n8905), .B0(n8904), .Y(n8907) );
  OAI221XL U8959 ( .A0(n8918), .A1(M2[10]), .B0(n8918), .B1(n8908), .C0(n8907), 
        .Y(n8912) );
  OAI222XL U8960 ( .A0(n8908), .A1(M2[10]), .B0(n8919), .B1(M2[11]), .C0(n8920), .C1(M2[12]), .Y(n8911) );
  AND2X1 U8961 ( .A(M2[11]), .B(n8919), .Y(n8909) );
  OAI222XL U8962 ( .A0(M2[12]), .A1(n8920), .B0(M2[12]), .B1(n8909), .C0(n8909), .C1(n8920), .Y(n8910) );
  OAI21XL U8963 ( .A0(n8912), .A1(n8911), .B0(n8910), .Y(n8913) );
endmodule


module Visible_Watermarking ( PADDR, PENABLE, PSEL, PWDATA, PWRITE, clk, rst, 
        Image_Done, Pixel_Data, new_pixel );
  input [9:0] PADDR;
  input [15:0] PWDATA;
  output [7:0] Pixel_Data;
  input PENABLE, PSEL, PWRITE, clk, rst;
  output Image_Done, new_pixel;
  wire   Block_Done, Ready, Image_Done1, ena_out, dout, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35;
  wire   [19:0] M2;
  wire   [31:0] block_out;
  wire   [31:0] Im_block;
  wire   [31:0] W_block;
  wire   [46:0] params;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16;

  Block_To_Pixel U_1 ( .clk(clk), .rst(n1), .M2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        M2[2:0]}), .block_in(block_out), .block_done(Block_Done), .Pixel_Data(
        Pixel_Data), .Ready(Ready), .new_pixel(new_pixel), .last_Block(
        Image_Done1), .Image_Done(Image_Done) );
  Equation_Implementation U_2 ( .Im_block(Im_block), .Ready(Ready), .W_block(
        W_block), .clk(clk), .ena_in(ena_out), .params(params), .rst(n1), 
        .block_done(Block_Done), .block_out(block_out), .M2({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, M2[2:0]}) );
  Control_And_Registers U_0 ( .clk(clk), .rst(n1), .ena_in(dout), .Address({
        n19, n18, n17, n16, n15, n14, n13, n12, n11, n10}), .data_in({n9, n8, 
        n7, n6, n5, n4, n3, n2, n34, n32, n30, n28, n26, n24, n22, n20}), 
        .ena_out(ena_out), .Image_Done(Image_Done1), .Block_Done(Block_Done), 
        .params(params), .Im_block(Im_block), .W_block(W_block) );
  INVX1 U2 ( .A(n21), .Y(n20) );
  INVX1 U3 ( .A(PWDATA[0]), .Y(n21) );
  INVX1 U4 ( .A(n23), .Y(n22) );
  INVX1 U5 ( .A(PWDATA[1]), .Y(n23) );
  INVX1 U6 ( .A(n25), .Y(n24) );
  INVX1 U7 ( .A(PWDATA[2]), .Y(n25) );
  INVX1 U8 ( .A(n27), .Y(n26) );
  INVX1 U9 ( .A(PWDATA[3]), .Y(n27) );
  INVX1 U10 ( .A(n29), .Y(n28) );
  INVX1 U11 ( .A(PWDATA[4]), .Y(n29) );
  INVX1 U12 ( .A(n31), .Y(n30) );
  INVX1 U13 ( .A(PWDATA[5]), .Y(n31) );
  INVX1 U14 ( .A(n33), .Y(n32) );
  INVX1 U15 ( .A(PWDATA[6]), .Y(n33) );
  INVX1 U16 ( .A(n35), .Y(n34) );
  INVX1 U17 ( .A(PWDATA[7]), .Y(n35) );
  BUFX3 U18 ( .A(PWDATA[8]), .Y(n2) );
  BUFX3 U19 ( .A(PWDATA[11]), .Y(n5) );
  BUFX3 U20 ( .A(PWDATA[10]), .Y(n4) );
  BUFX3 U21 ( .A(PWDATA[9]), .Y(n3) );
  BUFX3 U22 ( .A(PWDATA[12]), .Y(n6) );
  BUFX3 U23 ( .A(PWDATA[14]), .Y(n8) );
  BUFX3 U24 ( .A(PWDATA[13]), .Y(n7) );
  BUFX3 U25 ( .A(PWDATA[15]), .Y(n9) );
  BUFX3 U26 ( .A(PADDR[2]), .Y(n12) );
  BUFX3 U27 ( .A(PADDR[6]), .Y(n16) );
  BUFX3 U28 ( .A(PADDR[1]), .Y(n11) );
  BUFX3 U29 ( .A(PADDR[5]), .Y(n15) );
  BUFX3 U30 ( .A(PADDR[0]), .Y(n10) );
  BUFX3 U31 ( .A(PADDR[4]), .Y(n14) );
  BUFX3 U32 ( .A(PADDR[9]), .Y(n19) );
  BUFX3 U33 ( .A(PADDR[3]), .Y(n13) );
  BUFX3 U34 ( .A(PADDR[8]), .Y(n18) );
  BUFX3 U35 ( .A(PADDR[7]), .Y(n17) );
  AND3X2 U36 ( .A(PSEL), .B(PENABLE), .C(PWRITE), .Y(dout) );
  BUFX3 U37 ( .A(rst), .Y(n1) );
endmodule

